
module EXUNIT_N32 ( NPC1, RD1, A, B, IMM, S1_A_NPC, S2_IMM_B, ALU_OPCODE, CLK, 
        RST, JUMP_EN, EN_REGN_ALU_OUT, JUMP, ALUOUT, ALU_OUT_REGN, B_OUT_REGN, 
        NPC2, RD2_OUT_REGN );
  input [31:0] NPC1;
  input [4:0] RD1;
  input [31:0] A;
  input [31:0] B;
  input [31:0] IMM;
  input [5:0] ALU_OPCODE;
  input [1:0] JUMP_EN;
  output [31:0] ALUOUT;
  output [31:0] ALU_OUT_REGN;
  output [31:0] B_OUT_REGN;
  output [31:0] NPC2;
  output [4:0] RD2_OUT_REGN;
  input S1_A_NPC, S2_IMM_B, CLK, RST, EN_REGN_ALU_OUT;
  output JUMP;
  wire   \COMP_41_1MPX/n4 , \COMP_ALU/ADD_SUB/carries_s[0] ,
         \COMP_REGN_ALUOUT/ffi_31/n5 , \COMP_REGN_ALUOUT/ffi_31/n4 ,
         \COMP_REGN_ALUOUT/ffi_30/n5 , \COMP_REGN_ALUOUT/ffi_30/n4 ,
         \COMP_REGN_ALUOUT/ffi_29/n5 , \COMP_REGN_ALUOUT/ffi_29/n4 ,
         \COMP_REGN_ALUOUT/ffi_28/n5 , \COMP_REGN_ALUOUT/ffi_28/n4 ,
         \COMP_REGN_ALUOUT/ffi_27/n5 , \COMP_REGN_ALUOUT/ffi_27/n4 ,
         \COMP_REGN_ALUOUT/ffi_26/n5 , \COMP_REGN_ALUOUT/ffi_26/n4 ,
         \COMP_REGN_ALUOUT/ffi_25/n5 , \COMP_REGN_ALUOUT/ffi_25/n4 ,
         \COMP_REGN_ALUOUT/ffi_24/n5 , \COMP_REGN_ALUOUT/ffi_24/n4 ,
         \COMP_REGN_ALUOUT/ffi_23/n5 , \COMP_REGN_ALUOUT/ffi_23/n4 ,
         \COMP_REGN_ALUOUT/ffi_22/n5 , \COMP_REGN_ALUOUT/ffi_22/n4 ,
         \COMP_REGN_ALUOUT/ffi_21/n5 , \COMP_REGN_ALUOUT/ffi_21/n4 ,
         \COMP_REGN_ALUOUT/ffi_20/n5 , \COMP_REGN_ALUOUT/ffi_20/n4 ,
         \COMP_REGN_ALUOUT/ffi_19/n5 , \COMP_REGN_ALUOUT/ffi_19/n4 ,
         \COMP_REGN_ALUOUT/ffi_18/n5 , \COMP_REGN_ALUOUT/ffi_18/n4 ,
         \COMP_REGN_ALUOUT/ffi_17/n5 , \COMP_REGN_ALUOUT/ffi_17/n4 ,
         \COMP_REGN_ALUOUT/ffi_16/n5 , \COMP_REGN_ALUOUT/ffi_16/n4 ,
         \COMP_REGN_ALUOUT/ffi_15/n5 , \COMP_REGN_ALUOUT/ffi_15/n4 ,
         \COMP_REGN_ALUOUT/ffi_14/n5 , \COMP_REGN_ALUOUT/ffi_14/n4 ,
         \COMP_REGN_ALUOUT/ffi_13/n5 , \COMP_REGN_ALUOUT/ffi_13/n4 ,
         \COMP_REGN_ALUOUT/ffi_12/n5 , \COMP_REGN_ALUOUT/ffi_12/n4 ,
         \COMP_REGN_ALUOUT/ffi_11/n5 , \COMP_REGN_ALUOUT/ffi_11/n4 ,
         \COMP_REGN_ALUOUT/ffi_10/n5 , \COMP_REGN_ALUOUT/ffi_10/n4 ,
         \COMP_REGN_ALUOUT/ffi_9/n5 , \COMP_REGN_ALUOUT/ffi_9/n4 ,
         \COMP_REGN_ALUOUT/ffi_8/n5 , \COMP_REGN_ALUOUT/ffi_8/n4 ,
         \COMP_REGN_ALUOUT/ffi_7/n5 , \COMP_REGN_ALUOUT/ffi_7/n4 ,
         \COMP_REGN_ALUOUT/ffi_6/n5 , \COMP_REGN_ALUOUT/ffi_6/n4 ,
         \COMP_REGN_ALUOUT/ffi_5/n5 , \COMP_REGN_ALUOUT/ffi_5/n4 ,
         \COMP_REGN_ALUOUT/ffi_4/n5 , \COMP_REGN_ALUOUT/ffi_4/n4 ,
         \COMP_REGN_ALUOUT/ffi_3/n5 , \COMP_REGN_ALUOUT/ffi_3/n4 ,
         \COMP_REGN_ALUOUT/ffi_2/n5 , \COMP_REGN_ALUOUT/ffi_2/n4 ,
         \COMP_REGN_ALUOUT/ffi_1/n5 , \COMP_REGN_ALUOUT/ffi_1/n4 ,
         \COMP_REGN_BOUT/ffi_31/n5 , \COMP_REGN_BOUT/ffi_31/n4 ,
         \COMP_REGN_BOUT/ffi_30/n5 , \COMP_REGN_BOUT/ffi_30/n4 ,
         \COMP_REGN_BOUT/ffi_29/n5 , \COMP_REGN_BOUT/ffi_29/n4 ,
         \COMP_REGN_BOUT/ffi_28/n5 , \COMP_REGN_BOUT/ffi_28/n4 ,
         \COMP_REGN_BOUT/ffi_27/n5 , \COMP_REGN_BOUT/ffi_27/n4 ,
         \COMP_REGN_BOUT/ffi_26/n5 , \COMP_REGN_BOUT/ffi_26/n4 ,
         \COMP_REGN_BOUT/ffi_25/n5 , \COMP_REGN_BOUT/ffi_25/n4 ,
         \COMP_REGN_BOUT/ffi_24/n5 , \COMP_REGN_BOUT/ffi_24/n4 ,
         \COMP_REGN_BOUT/ffi_23/n5 , \COMP_REGN_BOUT/ffi_23/n4 ,
         \COMP_REGN_BOUT/ffi_22/n5 , \COMP_REGN_BOUT/ffi_22/n4 ,
         \COMP_REGN_BOUT/ffi_21/n5 , \COMP_REGN_BOUT/ffi_21/n4 ,
         \COMP_REGN_BOUT/ffi_20/n5 , \COMP_REGN_BOUT/ffi_20/n4 ,
         \COMP_REGN_BOUT/ffi_19/n5 , \COMP_REGN_BOUT/ffi_19/n4 ,
         \COMP_REGN_BOUT/ffi_18/n5 , \COMP_REGN_BOUT/ffi_18/n4 ,
         \COMP_REGN_BOUT/ffi_17/n5 , \COMP_REGN_BOUT/ffi_17/n4 ,
         \COMP_REGN_BOUT/ffi_16/n5 , \COMP_REGN_BOUT/ffi_16/n4 ,
         \COMP_REGN_BOUT/ffi_15/n5 , \COMP_REGN_BOUT/ffi_15/n4 ,
         \COMP_REGN_BOUT/ffi_14/n5 , \COMP_REGN_BOUT/ffi_14/n4 ,
         \COMP_REGN_BOUT/ffi_13/n5 , \COMP_REGN_BOUT/ffi_13/n4 ,
         \COMP_REGN_BOUT/ffi_12/n5 , \COMP_REGN_BOUT/ffi_12/n4 ,
         \COMP_REGN_BOUT/ffi_11/n5 , \COMP_REGN_BOUT/ffi_11/n4 ,
         \COMP_REGN_BOUT/ffi_10/n5 , \COMP_REGN_BOUT/ffi_10/n4 ,
         \COMP_REGN_BOUT/ffi_9/n5 , \COMP_REGN_BOUT/ffi_9/n4 ,
         \COMP_REGN_BOUT/ffi_8/n5 , \COMP_REGN_BOUT/ffi_8/n4 ,
         \COMP_REGN_BOUT/ffi_7/n5 , \COMP_REGN_BOUT/ffi_7/n4 ,
         \COMP_REGN_BOUT/ffi_6/n5 , \COMP_REGN_BOUT/ffi_6/n4 ,
         \COMP_REGN_BOUT/ffi_5/n5 , \COMP_REGN_BOUT/ffi_5/n4 ,
         \COMP_REGN_BOUT/ffi_4/n5 , \COMP_REGN_BOUT/ffi_4/n4 ,
         \COMP_REGN_BOUT/ffi_3/n5 , \COMP_REGN_BOUT/ffi_3/n4 ,
         \COMP_REGN_BOUT/ffi_2/n5 , \COMP_REGN_BOUT/ffi_2/n4 ,
         \COMP_REGN_BOUT/ffi_1/n5 , \COMP_REGN_BOUT/ffi_1/n4 ,
         \COMP_REGN_BOUT/ffi_0/n5 , \COMP_REGN_BOUT/ffi_0/n4 , n2, n2394,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
  assign \COMP_ALU/ADD_SUB/carries_s[0]  = ALU_OPCODE[0];

  DFF_X1 \COMP_REGN_ALUOUT/ffi_31/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_31/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[31]), .QN(\COMP_REGN_ALUOUT/ffi_31/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_30/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_30/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[30]), .QN(\COMP_REGN_ALUOUT/ffi_30/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_29/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_29/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[29]), .QN(\COMP_REGN_ALUOUT/ffi_29/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_28/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_28/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[28]), .QN(\COMP_REGN_ALUOUT/ffi_28/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_27/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_27/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[27]), .QN(\COMP_REGN_ALUOUT/ffi_27/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_26/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_26/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[26]), .QN(\COMP_REGN_ALUOUT/ffi_26/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_25/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_25/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[25]), .QN(\COMP_REGN_ALUOUT/ffi_25/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_24/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_24/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[24]), .QN(\COMP_REGN_ALUOUT/ffi_24/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_23/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_23/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[23]), .QN(\COMP_REGN_ALUOUT/ffi_23/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_22/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_22/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[22]), .QN(\COMP_REGN_ALUOUT/ffi_22/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_21/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_21/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[21]), .QN(\COMP_REGN_ALUOUT/ffi_21/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_20/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_20/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[20]), .QN(\COMP_REGN_ALUOUT/ffi_20/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_19/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_19/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[19]), .QN(\COMP_REGN_ALUOUT/ffi_19/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_18/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_18/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[18]), .QN(\COMP_REGN_ALUOUT/ffi_18/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_17/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_17/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[17]), .QN(\COMP_REGN_ALUOUT/ffi_17/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_16/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_16/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[16]), .QN(\COMP_REGN_ALUOUT/ffi_16/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_15/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_15/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[15]), .QN(\COMP_REGN_ALUOUT/ffi_15/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_14/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_14/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[14]), .QN(\COMP_REGN_ALUOUT/ffi_14/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_13/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_13/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[13]), .QN(\COMP_REGN_ALUOUT/ffi_13/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_12/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_12/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[12]), .QN(\COMP_REGN_ALUOUT/ffi_12/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_11/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_11/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[11]), .QN(\COMP_REGN_ALUOUT/ffi_11/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_10/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_10/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[10]), .QN(\COMP_REGN_ALUOUT/ffi_10/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_8/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_8/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[8]), .QN(\COMP_REGN_ALUOUT/ffi_8/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_7/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_7/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[7]), .QN(\COMP_REGN_ALUOUT/ffi_7/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_4/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_4/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[4]), .QN(\COMP_REGN_ALUOUT/ffi_4/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_3/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_3/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[3]), .QN(\COMP_REGN_ALUOUT/ffi_3/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_2/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_2/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[2]), .QN(\COMP_REGN_ALUOUT/ffi_2/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_0/Q_reg  ( .D(n2), .CK(CLK), .Q(n2394) );
  DFF_X1 \COMP_REGN_BOUT/ffi_31/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_31/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[31]), .QN(\COMP_REGN_BOUT/ffi_31/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_30/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_30/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[30]), .QN(\COMP_REGN_BOUT/ffi_30/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_29/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_29/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[29]), .QN(\COMP_REGN_BOUT/ffi_29/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_28/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_28/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[28]), .QN(\COMP_REGN_BOUT/ffi_28/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_27/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_27/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[27]), .QN(\COMP_REGN_BOUT/ffi_27/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_26/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_26/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[26]), .QN(\COMP_REGN_BOUT/ffi_26/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_25/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_25/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[25]), .QN(\COMP_REGN_BOUT/ffi_25/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_24/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_24/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[24]), .QN(\COMP_REGN_BOUT/ffi_24/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_23/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_23/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[23]), .QN(\COMP_REGN_BOUT/ffi_23/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_22/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_22/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[22]), .QN(\COMP_REGN_BOUT/ffi_22/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_21/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_21/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[21]), .QN(\COMP_REGN_BOUT/ffi_21/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_20/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_20/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[20]), .QN(\COMP_REGN_BOUT/ffi_20/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_19/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_19/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[19]), .QN(\COMP_REGN_BOUT/ffi_19/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_18/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_18/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[18]), .QN(\COMP_REGN_BOUT/ffi_18/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_17/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_17/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[17]), .QN(\COMP_REGN_BOUT/ffi_17/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_16/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_16/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[16]), .QN(\COMP_REGN_BOUT/ffi_16/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_15/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_15/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[15]), .QN(\COMP_REGN_BOUT/ffi_15/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_14/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_14/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[14]), .QN(\COMP_REGN_BOUT/ffi_14/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_13/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_13/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[13]), .QN(\COMP_REGN_BOUT/ffi_13/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_12/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_12/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[12]), .QN(\COMP_REGN_BOUT/ffi_12/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_11/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_11/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[11]), .QN(\COMP_REGN_BOUT/ffi_11/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_10/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_10/n5 ), .CK(
        CLK), .Q(B_OUT_REGN[10]), .QN(\COMP_REGN_BOUT/ffi_10/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_9/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_9/n5 ), .CK(CLK), .Q(B_OUT_REGN[9]), .QN(\COMP_REGN_BOUT/ffi_9/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_8/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_8/n5 ), .CK(CLK), .Q(B_OUT_REGN[8]), .QN(\COMP_REGN_BOUT/ffi_8/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_7/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_7/n5 ), .CK(CLK), .Q(B_OUT_REGN[7]), .QN(\COMP_REGN_BOUT/ffi_7/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_6/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_6/n5 ), .CK(CLK), .Q(B_OUT_REGN[6]), .QN(\COMP_REGN_BOUT/ffi_6/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_5/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_5/n5 ), .CK(CLK), .Q(B_OUT_REGN[5]), .QN(\COMP_REGN_BOUT/ffi_5/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_4/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_4/n5 ), .CK(CLK), .Q(B_OUT_REGN[4]), .QN(\COMP_REGN_BOUT/ffi_4/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_3/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_3/n5 ), .CK(CLK), .Q(B_OUT_REGN[3]), .QN(\COMP_REGN_BOUT/ffi_3/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_2/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_2/n5 ), .CK(CLK), .Q(B_OUT_REGN[2]), .QN(\COMP_REGN_BOUT/ffi_2/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_1/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_1/n5 ), .CK(CLK), .Q(B_OUT_REGN[1]), .QN(\COMP_REGN_BOUT/ffi_1/n4 ) );
  DFF_X1 \COMP_REGN_BOUT/ffi_0/Q_reg  ( .D(\COMP_REGN_BOUT/ffi_0/n5 ), .CK(CLK), .Q(B_OUT_REGN[0]), .QN(\COMP_REGN_BOUT/ffi_0/n4 ) );
  DFF_X1 \COMP_NPC2/ffi_31/Q_reg  ( .D(n2393), .CK(CLK), .QN(NPC2[31]) );
  DFF_X1 \COMP_REG5_RD2OUT/ffi_4/Q_reg  ( .D(n2361), .CK(CLK), .QN(
        RD2_OUT_REGN[4]) );
  DFF_X1 \COMP_REG5_RD2OUT/ffi_3/Q_reg  ( .D(n2360), .CK(CLK), .QN(
        RD2_OUT_REGN[3]) );
  DFF_X1 \COMP_REG5_RD2OUT/ffi_2/Q_reg  ( .D(n2359), .CK(CLK), .QN(
        RD2_OUT_REGN[2]) );
  DFF_X1 \COMP_REG5_RD2OUT/ffi_1/Q_reg  ( .D(n2358), .CK(CLK), .QN(
        RD2_OUT_REGN[1]) );
  DFF_X1 \COMP_REG5_RD2OUT/ffi_0/Q_reg  ( .D(n2357), .CK(CLK), .QN(
        RD2_OUT_REGN[0]) );
  DFF_X1 \COMP_NPC2/ffi_30/Q_reg  ( .D(n2392), .CK(CLK), .QN(NPC2[30]) );
  DFF_X1 \COMP_NPC2/ffi_29/Q_reg  ( .D(n2391), .CK(CLK), .QN(NPC2[29]) );
  DFF_X1 \COMP_NPC2/ffi_28/Q_reg  ( .D(n2390), .CK(CLK), .QN(NPC2[28]) );
  DFF_X1 \COMP_NPC2/ffi_27/Q_reg  ( .D(n2389), .CK(CLK), .QN(NPC2[27]) );
  DFF_X1 \COMP_NPC2/ffi_26/Q_reg  ( .D(n2388), .CK(CLK), .QN(NPC2[26]) );
  DFF_X1 \COMP_NPC2/ffi_25/Q_reg  ( .D(n2387), .CK(CLK), .QN(NPC2[25]) );
  DFF_X1 \COMP_NPC2/ffi_24/Q_reg  ( .D(n2386), .CK(CLK), .QN(NPC2[24]) );
  DFF_X1 \COMP_NPC2/ffi_23/Q_reg  ( .D(n2385), .CK(CLK), .QN(NPC2[23]) );
  DFF_X1 \COMP_NPC2/ffi_22/Q_reg  ( .D(n2384), .CK(CLK), .QN(NPC2[22]) );
  DFF_X1 \COMP_NPC2/ffi_21/Q_reg  ( .D(n2383), .CK(CLK), .QN(NPC2[21]) );
  DFF_X1 \COMP_NPC2/ffi_20/Q_reg  ( .D(n2382), .CK(CLK), .QN(NPC2[20]) );
  DFF_X1 \COMP_NPC2/ffi_19/Q_reg  ( .D(n2381), .CK(CLK), .QN(NPC2[19]) );
  DFF_X1 \COMP_NPC2/ffi_18/Q_reg  ( .D(n2380), .CK(CLK), .QN(NPC2[18]) );
  DFF_X1 \COMP_NPC2/ffi_17/Q_reg  ( .D(n2379), .CK(CLK), .QN(NPC2[17]) );
  DFF_X1 \COMP_NPC2/ffi_16/Q_reg  ( .D(n2378), .CK(CLK), .QN(NPC2[16]) );
  DFF_X1 \COMP_NPC2/ffi_15/Q_reg  ( .D(n2377), .CK(CLK), .QN(NPC2[15]) );
  DFF_X1 \COMP_NPC2/ffi_14/Q_reg  ( .D(n2376), .CK(CLK), .QN(NPC2[14]) );
  DFF_X1 \COMP_NPC2/ffi_13/Q_reg  ( .D(n2375), .CK(CLK), .QN(NPC2[13]) );
  DFF_X1 \COMP_NPC2/ffi_12/Q_reg  ( .D(n2374), .CK(CLK), .QN(NPC2[12]) );
  DFF_X1 \COMP_NPC2/ffi_11/Q_reg  ( .D(n2373), .CK(CLK), .QN(NPC2[11]) );
  DFF_X1 \COMP_NPC2/ffi_10/Q_reg  ( .D(n2372), .CK(CLK), .QN(NPC2[10]) );
  DFF_X1 \COMP_NPC2/ffi_9/Q_reg  ( .D(n2371), .CK(CLK), .QN(NPC2[9]) );
  DFF_X1 \COMP_NPC2/ffi_8/Q_reg  ( .D(n2370), .CK(CLK), .QN(NPC2[8]) );
  DFF_X1 \COMP_NPC2/ffi_7/Q_reg  ( .D(n2369), .CK(CLK), .QN(NPC2[7]) );
  DFF_X1 \COMP_NPC2/ffi_6/Q_reg  ( .D(n2368), .CK(CLK), .QN(NPC2[6]) );
  DFF_X1 \COMP_NPC2/ffi_5/Q_reg  ( .D(n2367), .CK(CLK), .QN(NPC2[5]) );
  DFF_X1 \COMP_NPC2/ffi_4/Q_reg  ( .D(n2366), .CK(CLK), .QN(NPC2[4]) );
  DFF_X1 \COMP_NPC2/ffi_3/Q_reg  ( .D(n2365), .CK(CLK), .QN(NPC2[3]) );
  DFF_X1 \COMP_NPC2/ffi_2/Q_reg  ( .D(n2364), .CK(CLK), .QN(NPC2[2]) );
  DFF_X1 \COMP_NPC2/ffi_1/Q_reg  ( .D(n2363), .CK(CLK), .QN(NPC2[1]) );
  DFF_X1 \COMP_NPC2/ffi_0/Q_reg  ( .D(n2362), .CK(CLK), .QN(NPC2[0]) );
  DFFS_X1 \COMP_REGN_ALUOUT/ffi_9/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_9/n5 ), 
        .CK(CLK), .SN(1'b1), .Q(ALU_OUT_REGN[9]), .QN(
        \COMP_REGN_ALUOUT/ffi_9/n4 ) );
  DFFS_X1 \COMP_REGN_ALUOUT/ffi_5/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_5/n5 ), 
        .CK(CLK), .SN(1'b1), .Q(ALU_OUT_REGN[5]), .QN(
        \COMP_REGN_ALUOUT/ffi_5/n4 ) );
  DFFS_X1 \COMP_REGN_ALUOUT/ffi_1/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_1/n5 ), 
        .CK(CLK), .SN(1'b1), .QN(\COMP_REGN_ALUOUT/ffi_1/n4 ) );
  DFF_X1 \COMP_REGN_ALUOUT/ffi_6/Q_reg  ( .D(\COMP_REGN_ALUOUT/ffi_6/n5 ), 
        .CK(CLK), .Q(ALU_OUT_REGN[6]), .QN(\COMP_REGN_ALUOUT/ffi_6/n4 ) );
  BUF_X2 U1127 ( .A(S2_IMM_B), .Z(n1382) );
  BUF_X2 U1128 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .Z(n1372) );
  INV_X1 U1129 ( .A(n1739), .ZN(n1578) );
  NAND2_X1 U1130 ( .A1(n1568), .A2(n2103), .ZN(n1739) );
  XNOR2_X1 U1131 ( .A(n1944), .B(n1377), .ZN(n1568) );
  OAI21_X1 U1132 ( .B1(n1381), .B2(n1031), .A(n1030), .ZN(n1944) );
  NAND2_X1 U1133 ( .A1(n1381), .A2(B[16]), .ZN(n1030) );
  INV_X1 U1134 ( .A(IMM[16]), .ZN(n1031) );
  AND2_X2 U1135 ( .A1(n1035), .A2(n1034), .ZN(n1708) );
  NAND3_X2 U1136 ( .A1(n1035), .A2(n1034), .A3(n1245), .ZN(n1039) );
  NAND2_X1 U1137 ( .A1(n1033), .A2(n1032), .ZN(n1245) );
  INV_X1 U1138 ( .A(n1633), .ZN(n1032) );
  INV_X1 U1139 ( .A(n1600), .ZN(n1033) );
  INV_X1 U1140 ( .A(n1604), .ZN(n1034) );
  NAND2_X1 U1141 ( .A1(n1637), .A2(n1634), .ZN(n1035) );
  NAND2_X2 U1142 ( .A1(n1039), .A2(n1342), .ZN(n1341) );
  AND2_X2 U1143 ( .A1(n1039), .A2(n1036), .ZN(n1339) );
  INV_X2 U1144 ( .A(n1037), .ZN(n1036) );
  NAND2_X2 U1145 ( .A1(n1038), .A2(n1342), .ZN(n1037) );
  INV_X2 U1146 ( .A(n1620), .ZN(n1038) );
  OR2_X2 U1147 ( .A1(n2008), .A2(n2007), .ZN(n2154) );
  INV_X2 U1148 ( .A(n2199), .ZN(n2251) );
  NAND2_X2 U1149 ( .A1(n2235), .A2(n1429), .ZN(n2211) );
  NAND2_X2 U1150 ( .A1(n1950), .A2(n1949), .ZN(n2083) );
  BUF_X1 U1151 ( .A(n2135), .Z(n1040) );
  INV_X4 U1152 ( .A(n1365), .ZN(n1363) );
  AND2_X2 U1153 ( .A1(n1529), .A2(n1525), .ZN(n1549) );
  BUF_X2 U1154 ( .A(n2098), .Z(n1352) );
  INV_X1 U1155 ( .A(n2305), .ZN(n1181) );
  AND3_X1 U1156 ( .A1(n2144), .A2(n2055), .A3(n2077), .ZN(n1274) );
  INV_X1 U1157 ( .A(n2208), .ZN(n1041) );
  OAI21_X1 U1158 ( .B1(n1610), .B2(n1041), .A(n1611), .ZN(n1748) );
  AOI21_X1 U1159 ( .B1(n1145), .B2(n1701), .A(n1327), .ZN(n1042) );
  AOI21_X1 U1160 ( .B1(n1701), .B2(n1242), .A(n1042), .ZN(n1043) );
  OAI21_X1 U1161 ( .B1(n1736), .B2(n1143), .A(n1043), .ZN(n2019) );
  OAI21_X1 U1162 ( .B1(n2245), .B2(n2124), .A(n2211), .ZN(n1044) );
  OAI22_X1 U1163 ( .A1(n2244), .A2(n2122), .B1(n2121), .B2(n2239), .ZN(n1045)
         );
  AOI211_X1 U1164 ( .C1(n2123), .C2(n2210), .A(n1044), .B(n1045), .ZN(n2254)
         );
  OAI22_X1 U1165 ( .A1(n2110), .A2(n2227), .B1(n2111), .B2(n1240), .ZN(n1046)
         );
  NOR3_X1 U1166 ( .A1(n2113), .A2(n2114), .A3(n1046), .ZN(n1047) );
  INV_X1 U1167 ( .A(n2117), .ZN(n1048) );
  AOI22_X1 U1168 ( .A1(n2117), .A2(n2170), .B1(n2168), .B2(n1048), .ZN(n1049)
         );
  AOI221_X1 U1169 ( .B1(n2169), .B2(n1048), .C1(n2171), .C2(n2117), .A(n2118), 
        .ZN(n1050) );
  AOI21_X1 U1170 ( .B1(n2118), .B2(n1049), .A(n1050), .ZN(n1051) );
  NAND2_X1 U1171 ( .A1(n2115), .A2(n1161), .ZN(n1052) );
  OAI211_X1 U1172 ( .C1(n1047), .C2(n2268), .A(n1051), .B(n1052), .ZN(
        ALUOUT[24]) );
  NAND2_X1 U1173 ( .A1(n1487), .A2(n1154), .ZN(n1053) );
  OAI21_X1 U1174 ( .B1(n1053), .B2(n1512), .A(n1511), .ZN(n1528) );
  NAND3_X1 U1175 ( .A1(n1351), .A2(n1258), .A3(n1237), .ZN(n1054) );
  NAND2_X1 U1176 ( .A1(n1237), .A2(n1308), .ZN(n1055) );
  NAND3_X1 U1177 ( .A1(n1055), .A2(n1339), .A3(n1054), .ZN(n1719) );
  AOI211_X1 U1178 ( .C1(ALU_OPCODE[1]), .C2(n1768), .A(n1751), .B(
        ALU_OPCODE[3]), .ZN(n1056) );
  INV_X1 U1179 ( .A(n1056), .ZN(n1057) );
  AOI21_X1 U1180 ( .B1(ALU_OPCODE[2]), .B2(n1176), .A(n1057), .ZN(n1338) );
  MUX2_X1 U1181 ( .A(n1702), .B(n1145), .S(n1701), .Z(n2001) );
  OAI21_X1 U1182 ( .B1(n2245), .B2(n2134), .A(n2211), .ZN(n1058) );
  OAI22_X1 U1183 ( .A1(n2244), .A2(n2132), .B1(n2131), .B2(n2239), .ZN(n1059)
         );
  AOI211_X1 U1184 ( .C1(n2133), .C2(n2210), .A(n1058), .B(n1059), .ZN(n2261)
         );
  INV_X1 U1185 ( .A(n2119), .ZN(n1060) );
  AOI22_X1 U1186 ( .A1(n2119), .A2(n2170), .B1(n2168), .B2(n1060), .ZN(n1061)
         );
  AOI221_X1 U1187 ( .B1(n2171), .B2(n2119), .C1(n2169), .C2(n1060), .A(n2120), 
        .ZN(n1062) );
  AOI21_X1 U1188 ( .B1(n2120), .B2(n1061), .A(n1062), .ZN(n1063) );
  AOI22_X1 U1189 ( .A1(n2154), .A2(n1361), .B1(n2176), .B2(n1184), .ZN(n1064)
         );
  AOI22_X1 U1190 ( .A1(n2221), .A2(n2173), .B1(n2177), .B2(n2260), .ZN(n1065)
         );
  AOI22_X1 U1191 ( .A1(n2224), .A2(n1358), .B1(n2225), .B2(n1355), .ZN(n1066)
         );
  AOI22_X1 U1192 ( .A1(n1040), .A2(n1359), .B1(n2125), .B2(n2222), .ZN(n1067)
         );
  OAI211_X1 U1193 ( .C1(n2251), .C2(n2265), .A(n1066), .B(n1067), .ZN(n1068)
         );
  NAND2_X1 U1194 ( .A1(n1064), .A2(n1065), .ZN(n1069) );
  OAI21_X1 U1195 ( .B1(n1068), .B2(n1069), .A(n2230), .ZN(n1070) );
  OAI211_X1 U1196 ( .C1(n2126), .C2(n2276), .A(n1063), .B(n1070), .ZN(
        ALUOUT[25]) );
  INV_X1 U1197 ( .A(n1353), .ZN(n1071) );
  INV_X1 U1198 ( .A(n2050), .ZN(n1072) );
  OAI221_X1 U1199 ( .B1(n2050), .B2(n1071), .C1(n1072), .C2(n1353), .A(n2194), 
        .ZN(n1630) );
  NOR2_X1 U1200 ( .A1(n1170), .A2(n1556), .ZN(n1073) );
  NAND2_X1 U1201 ( .A1(n1557), .A2(n1073), .ZN(n1640) );
  INV_X1 U1202 ( .A(n2196), .ZN(n1074) );
  OAI21_X1 U1203 ( .B1(n1607), .B2(n1074), .A(n1710), .ZN(n1712) );
  INV_X1 U1204 ( .A(n1773), .ZN(n1075) );
  INV_X1 U1205 ( .A(n2262), .ZN(n1076) );
  AOI222_X1 U1206 ( .A1(n1075), .A2(n1076), .B1(n1852), .B2(n2173), .C1(n1360), 
        .C2(n1804), .ZN(n1517) );
  OAI22_X1 U1207 ( .A1(n2244), .A2(n1885), .B1(n1185), .B2(n2181), .ZN(n1077)
         );
  AOI211_X1 U1208 ( .C1(n1251), .C2(n2210), .A(n1930), .B(n1077), .ZN(n1078)
         );
  INV_X2 U1209 ( .A(n1078), .ZN(n2026) );
  INV_X1 U1210 ( .A(n2178), .ZN(n1079) );
  AOI22_X1 U1211 ( .A1(n2178), .A2(n2170), .B1(n2171), .B2(n1079), .ZN(n1080)
         );
  AOI221_X1 U1212 ( .B1(n2168), .B2(n2178), .C1(n2169), .C2(n1079), .A(n2172), 
        .ZN(n1081) );
  AOI21_X1 U1213 ( .B1(n2172), .B2(n1080), .A(n1081), .ZN(n1082) );
  OAI211_X1 U1214 ( .C1(n2265), .C2(n2217), .A(n2175), .B(n2174), .ZN(n1083)
         );
  OAI21_X1 U1215 ( .B1(n2190), .B2(n1083), .A(n2230), .ZN(n1084) );
  OAI211_X1 U1216 ( .C1(n2191), .C2(n2276), .A(n1082), .B(n1084), .ZN(
        ALUOUT[28]) );
  INV_X1 U1217 ( .A(n1550), .ZN(n1085) );
  NAND3_X1 U1218 ( .A1(n1335), .A2(n1334), .A3(n1178), .ZN(n1086) );
  NAND2_X1 U1219 ( .A1(n1086), .A2(n1085), .ZN(n1669) );
  OAI22_X1 U1220 ( .A1(n2244), .A2(n2193), .B1(n1185), .B2(n2040), .ZN(n1087)
         );
  AOI211_X1 U1221 ( .C1(n1897), .C2(n2210), .A(n1930), .B(n1087), .ZN(n1088)
         );
  INV_X2 U1222 ( .A(n1088), .ZN(n2043) );
  NOR2_X1 U1223 ( .A1(n1767), .A2(n1238), .ZN(n1089) );
  OAI21_X1 U1224 ( .B1(n1269), .B2(n1268), .A(n1338), .ZN(n1090) );
  NAND3_X1 U1225 ( .A1(n1266), .A2(n1089), .A3(n1090), .ZN(ALUOUT[0]) );
  NOR2_X1 U1226 ( .A1(n1626), .A2(n1179), .ZN(n1091) );
  AOI211_X1 U1227 ( .C1(n1727), .C2(n1743), .A(n1587), .B(n1091), .ZN(n1314)
         );
  AND3_X1 U1228 ( .A1(n1176), .A2(ALU_OPCODE[3]), .A3(n1770), .ZN(n1238) );
  OAI22_X1 U1229 ( .A1(n2244), .A2(n2213), .B1(n1185), .B2(n1914), .ZN(n1092)
         );
  AOI211_X1 U1230 ( .C1(n2061), .C2(n2210), .A(n1930), .B(n1092), .ZN(n1093)
         );
  INV_X2 U1231 ( .A(n1093), .ZN(n2067) );
  INV_X1 U1232 ( .A(n1341), .ZN(n1094) );
  AOI21_X1 U1233 ( .B1(n1210), .B2(n1094), .A(n1209), .ZN(n1095) );
  OAI21_X1 U1234 ( .B1(n1341), .B2(n1293), .A(n1095), .ZN(n1096) );
  NAND2_X1 U1235 ( .A1(n1719), .A2(n1096), .ZN(n2191) );
  OAI22_X1 U1236 ( .A1(n2263), .A2(n2227), .B1(n2255), .B2(n2261), .ZN(n1097)
         );
  OAI22_X1 U1237 ( .A1(n2254), .A2(n2217), .B1(n2216), .B2(n1357), .ZN(n1098)
         );
  OAI22_X1 U1238 ( .A1(n2202), .A2(n2262), .B1(n2265), .B2(n1240), .ZN(n1099)
         );
  OR4_X1 U1239 ( .A1(n2203), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1100) );
  INV_X1 U1240 ( .A(n2204), .ZN(n1101) );
  AOI22_X1 U1241 ( .A1(n2204), .A2(n2233), .B1(n2232), .B2(n1101), .ZN(n1102)
         );
  OAI221_X1 U1242 ( .B1(n2204), .B2(n2236), .C1(n1101), .C2(n2234), .A(n2205), 
        .ZN(n1103) );
  OAI21_X1 U1243 ( .B1(n2205), .B2(n1102), .A(n1103), .ZN(n1104) );
  AOI21_X1 U1244 ( .B1(n2230), .B2(n1100), .A(n1104), .ZN(n1105) );
  OAI21_X1 U1245 ( .B1(n2206), .B2(n2276), .A(n1105), .ZN(ALUOUT[29]) );
  OR3_X1 U1246 ( .A1(n2243), .A2(n1618), .A3(n2274), .ZN(n1106) );
  AOI221_X1 U1247 ( .B1(n1617), .B2(n1106), .C1(n2235), .C2(n1106), .A(n1716), 
        .ZN(n1302) );
  NOR2_X1 U1248 ( .A1(n1732), .A2(n1329), .ZN(n1107) );
  NAND2_X1 U1249 ( .A1(n1107), .A2(n1626), .ZN(n1108) );
  OAI21_X1 U1250 ( .B1(n1730), .B2(n1731), .A(n1108), .ZN(n1326) );
  INV_X1 U1251 ( .A(n1652), .ZN(n1109) );
  AOI21_X1 U1252 ( .B1(n1659), .B2(n1177), .A(n1109), .ZN(n1110) );
  NAND2_X1 U1253 ( .A1(n1153), .A2(n1661), .ZN(n1111) );
  XNOR2_X1 U1254 ( .A(n1111), .B(n1110), .ZN(n1802) );
  NAND2_X1 U1255 ( .A1(n1335), .A2(n1246), .ZN(n1112) );
  INV_X1 U1256 ( .A(n1678), .ZN(n1113) );
  NAND3_X1 U1257 ( .A1(n1113), .A2(n1112), .A3(n1158), .ZN(n1114) );
  OAI211_X1 U1258 ( .C1(n1112), .C2(n1113), .A(n1114), .B(n1680), .ZN(n1862)
         );
  NOR2_X1 U1259 ( .A1(n2084), .A2(n2132), .ZN(n1115) );
  OAI22_X1 U1260 ( .A1(n1990), .A2(n1363), .B1(n2245), .B2(n2131), .ZN(n1116)
         );
  AOI211_X1 U1261 ( .C1(n2210), .C2(n1989), .A(n1115), .B(n1116), .ZN(n1117)
         );
  NAND2_X1 U1262 ( .A1(n2083), .A2(n1117), .ZN(n2135) );
  AOI22_X1 U1263 ( .A1(n2221), .A2(n2222), .B1(n2224), .B2(n1359), .ZN(n1118)
         );
  AOI211_X1 U1264 ( .C1(n2253), .C2(n1358), .A(n2218), .B(n2219), .ZN(n1119)
         );
  AOI22_X1 U1265 ( .A1(n2225), .A2(n1184), .B1(n2226), .B2(n1362), .ZN(n1120)
         );
  NAND3_X1 U1266 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1121) );
  INV_X1 U1267 ( .A(n2228), .ZN(n1122) );
  AOI22_X1 U1268 ( .A1(n2228), .A2(n2233), .B1(n2232), .B2(n1122), .ZN(n1123)
         );
  OAI221_X1 U1269 ( .B1(n2228), .B2(n2236), .C1(n1122), .C2(n2234), .A(n2229), 
        .ZN(n1124) );
  OAI21_X1 U1270 ( .B1(n1123), .B2(n2229), .A(n1124), .ZN(n1125) );
  AOI21_X1 U1271 ( .B1(n2230), .B2(n1121), .A(n1125), .ZN(n1126) );
  OAI21_X1 U1272 ( .B1(n1159), .B2(n2276), .A(n1126), .ZN(ALUOUT[30]) );
  NAND2_X2 U1273 ( .A1(n1954), .A2(n1352), .ZN(n2244) );
  BUF_X2 U1274 ( .A(S1_A_NPC), .Z(n1148) );
  AND2_X1 U1275 ( .A1(n1158), .A2(n1547), .ZN(n1127) );
  NAND2_X1 U1276 ( .A1(n1326), .A2(n1735), .ZN(n1128) );
  INV_X2 U1277 ( .A(\COMP_REGN_ALUOUT/ffi_1/n4 ), .ZN(ALU_OUT_REGN[1]) );
  OR2_X1 U1281 ( .A1(n2061), .A2(n1412), .ZN(n1527) );
  BUF_X1 U1282 ( .A(n1276), .Z(n1133) );
  BUF_X1 U1283 ( .A(n1525), .Z(n1134) );
  AND2_X1 U1284 ( .A1(n1454), .A2(n2131), .ZN(n1658) );
  INV_X1 U1285 ( .A(n1234), .ZN(n1135) );
  BUF_X1 U1286 ( .A(n1655), .Z(n1136) );
  BUF_X1 U1287 ( .A(n1654), .Z(n1137) );
  BUF_X1 U1288 ( .A(n1323), .Z(n1138) );
  AOI21_X1 U1289 ( .B1(n1637), .B2(n1634), .A(n1604), .ZN(n1139) );
  AND2_X1 U1290 ( .A1(n1394), .A2(n1661), .ZN(n1140) );
  NAND2_X1 U1291 ( .A1(n1440), .A2(n1788), .ZN(n1141) );
  AND2_X1 U1292 ( .A1(n1163), .A2(n1207), .ZN(n1142) );
  INV_X1 U1293 ( .A(n1737), .ZN(n1143) );
  AND2_X1 U1294 ( .A1(n1415), .A2(n2240), .ZN(n1144) );
  INV_X1 U1295 ( .A(n1702), .ZN(n1145) );
  XOR2_X1 U1296 ( .A(n2050), .B(n1353), .Z(n1146) );
  INV_X2 U1297 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1353) );
  INV_X1 U1298 ( .A(n1165), .ZN(n1147) );
  INV_X1 U1299 ( .A(n1813), .ZN(n2148) );
  AND2_X1 U1300 ( .A1(n1643), .A2(n1562), .ZN(n1149) );
  BUF_X1 U1301 ( .A(n1518), .Z(n1150) );
  BUF_X1 U1302 ( .A(n1944), .Z(n1151) );
  BUF_X1 U1303 ( .A(n1670), .Z(n1152) );
  BUF_X1 U1304 ( .A(n1662), .Z(n1153) );
  BUF_X1 U1305 ( .A(n1313), .Z(n1154) );
  BUF_X1 U1306 ( .A(n1553), .Z(n1155) );
  BUF_X1 U1307 ( .A(n1986), .Z(n1156) );
  AOI21_X1 U1308 ( .B1(n1293), .B2(n1250), .A(n1283), .ZN(n1282) );
  INV_X1 U1309 ( .A(n1332), .ZN(n1157) );
  OR2_X1 U1310 ( .A1(n1418), .A2(n1253), .ZN(n1158) );
  OR2_X1 U1311 ( .A1(n1418), .A2(n1253), .ZN(n1677) );
  CLKBUF_X1 U1312 ( .A(n1478), .Z(n1195) );
  CLKBUF_X1 U1313 ( .A(n1968), .Z(n1197) );
  BUF_X1 U1314 ( .A(n2231), .Z(n1159) );
  INV_X1 U1315 ( .A(n1172), .ZN(n1160) );
  BUF_X1 U1316 ( .A(n2116), .Z(n1161) );
  BUF_X1 U1317 ( .A(n1540), .Z(n1162) );
  OR2_X1 U1318 ( .A1(S2_IMM_B), .A2(n1208), .ZN(n1163) );
  NAND2_X1 U1319 ( .A1(n1163), .A2(n1207), .ZN(n2099) );
  XNOR2_X1 U1320 ( .A(n1478), .B(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1164)
         );
  INV_X1 U1321 ( .A(n2148), .ZN(n1165) );
  CLKBUF_X3 U1322 ( .A(S1_A_NPC), .Z(n1383) );
  NAND2_X1 U1323 ( .A1(n1229), .A2(n1623), .ZN(n1216) );
  BUF_X1 U1324 ( .A(n1741), .Z(n1166) );
  INV_X1 U1325 ( .A(S2_IMM_B), .ZN(n1167) );
  INV_X1 U1326 ( .A(n1167), .ZN(n1168) );
  BUF_X1 U1327 ( .A(n1409), .Z(n1169) );
  NAND3_X1 U1328 ( .A1(n1649), .A2(n1548), .A3(n1678), .ZN(n1170) );
  OR2_X1 U1329 ( .A1(n1554), .A2(n1555), .ZN(n1171) );
  INV_X1 U1330 ( .A(S2_IMM_B), .ZN(n1172) );
  INV_X1 U1331 ( .A(n1172), .ZN(n1173) );
  OR2_X1 U1332 ( .A1(n1738), .A2(n1728), .ZN(n1174) );
  XOR2_X1 U1333 ( .A(n2032), .B(n1354), .Z(n1175) );
  OAI21_X1 U1334 ( .B1(n1285), .B2(n1286), .A(n1282), .ZN(n1176) );
  NAND2_X1 U1335 ( .A1(n1408), .A2(n1137), .ZN(n1177) );
  CLKBUF_X3 U1336 ( .A(S2_IMM_B), .Z(n1380) );
  CLKBUF_X3 U1337 ( .A(S2_IMM_B), .Z(n1381) );
  AND2_X1 U1338 ( .A1(n1678), .A2(n1547), .ZN(n1178) );
  INV_X2 U1339 ( .A(n2262), .ZN(n2222) );
  INV_X2 U1340 ( .A(n2217), .ZN(n2260) );
  INV_X1 U1341 ( .A(n1727), .ZN(n1179) );
  AND2_X1 U1342 ( .A1(n2308), .A2(n1271), .ZN(n2210) );
  OR2_X1 U1343 ( .A1(n1446), .A2(n1465), .ZN(n2223) );
  OR2_X1 U1344 ( .A1(n1455), .A2(n1234), .ZN(n2227) );
  OR2_X1 U1345 ( .A1(n2249), .A2(n1376), .ZN(n2186) );
  BUF_X2 U1346 ( .A(n2220), .Z(n1358) );
  BUF_X1 U1347 ( .A(n1947), .Z(n1185) );
  INV_X1 U1348 ( .A(n2306), .ZN(n1180) );
  OAI211_X1 U1349 ( .C1(n1216), .C2(n1740), .A(n1217), .B(n1219), .ZN(n1985)
         );
  INV_X1 U1350 ( .A(n1237), .ZN(n1210) );
  INV_X1 U1351 ( .A(n1620), .ZN(n1209) );
  INV_X1 U1352 ( .A(n2223), .ZN(n1359) );
  INV_X1 U1353 ( .A(n2227), .ZN(n1362) );
  BUF_X1 U1354 ( .A(n1742), .Z(n1219) );
  INV_X1 U1355 ( .A(n2223), .ZN(n1360) );
  INV_X1 U1356 ( .A(n1623), .ZN(n1182) );
  INV_X1 U1357 ( .A(n2244), .ZN(n1365) );
  INV_X1 U1358 ( .A(n1705), .ZN(n1183) );
  INV_X1 U1359 ( .A(n2255), .ZN(n2173) );
  AND2_X1 U1360 ( .A1(n1313), .A2(n1487), .ZN(n1510) );
  NAND2_X1 U1361 ( .A1(n1718), .A2(n1709), .ZN(n1620) );
  AND2_X1 U1362 ( .A1(n1142), .A2(n2308), .ZN(n1954) );
  NAND2_X1 U1363 ( .A1(n1406), .A2(n1405), .ZN(n1656) );
  INV_X2 U1364 ( .A(n1240), .ZN(n1184) );
  BUF_X1 U1365 ( .A(n1236), .Z(n1642) );
  OR2_X1 U1366 ( .A1(n1674), .A2(n2118), .ZN(n1349) );
  INV_X1 U1367 ( .A(n2232), .ZN(n2169) );
  INV_X1 U1368 ( .A(n1759), .ZN(n1465) );
  INV_X1 U1369 ( .A(n2243), .ZN(n2235) );
  BUF_X4 U1370 ( .A(n2394), .Z(ALU_OUT_REGN[0]) );
  BUF_X2 U1371 ( .A(n2306), .Z(n1186) );
  OR2_X1 U1372 ( .A1(n1768), .A2(ALU_OPCODE[3]), .ZN(n1201) );
  BUF_X1 U1373 ( .A(n1781), .Z(n1200) );
  BUF_X2 U1374 ( .A(n2305), .Z(n1187) );
  INV_X1 U1375 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1378) );
  BUF_X1 U1376 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .Z(n1376) );
  XOR2_X1 U1377 ( .A(n2320), .B(JUMP_EN[0]), .Z(\COMP_41_1MPX/n4 ) );
  INV_X1 U1378 ( .A(\COMP_41_1MPX/n4 ), .ZN(JUMP) );
  BUF_X1 U1379 ( .A(n1847), .Z(n1189) );
  BUF_X1 U1380 ( .A(n2014), .Z(n1190) );
  AND2_X1 U1381 ( .A1(n1191), .A2(n1630), .ZN(n1589) );
  NAND2_X1 U1382 ( .A1(n1146), .A2(n2040), .ZN(n1191) );
  BUF_X1 U1383 ( .A(n1827), .Z(n1192) );
  BUF_X1 U1384 ( .A(n1834), .Z(n1193) );
  BUF_X1 U1385 ( .A(n1559), .Z(n1194) );
  NAND2_X1 U1386 ( .A1(n1276), .A2(n1644), .ZN(n1561) );
  XNOR2_X1 U1387 ( .A(n1553), .B(n2038), .ZN(n1276) );
  OAI21_X1 U1388 ( .B1(n1350), .B2(n1595), .A(n1734), .ZN(n1258) );
  AND2_X1 U1389 ( .A1(n1625), .A2(n1596), .ZN(n1350) );
  NAND2_X1 U1390 ( .A1(n1196), .A2(n1638), .ZN(n2126) );
  NAND2_X1 U1391 ( .A1(n1704), .A2(n1639), .ZN(n1638) );
  OR2_X1 U1392 ( .A1(n1221), .A2(n1639), .ZN(n1196) );
  NAND3_X1 U1393 ( .A1(n1275), .A2(n1274), .A3(n1224), .ZN(n1269) );
  NOR2_X1 U1394 ( .A1(n1738), .A2(n1728), .ZN(n1583) );
  NAND2_X1 U1395 ( .A1(n1628), .A2(n1588), .ZN(n1738) );
  OAI21_X1 U1396 ( .B1(n1381), .B2(n1199), .A(n1198), .ZN(n1986) );
  NAND2_X1 U1397 ( .A1(n1382), .A2(B[18]), .ZN(n1198) );
  INV_X1 U1398 ( .A(IMM[18]), .ZN(n1199) );
  NAND2_X1 U1399 ( .A1(n1578), .A2(n1694), .ZN(n1742) );
  XNOR2_X1 U1400 ( .A(n1579), .B(n2123), .ZN(n1694) );
  OR2_X1 U1401 ( .A1(n1769), .A2(n1201), .ZN(n1244) );
  NAND2_X1 U1402 ( .A1(n1314), .A2(n1202), .ZN(n1632) );
  NAND2_X1 U1403 ( .A1(n1229), .A2(n1203), .ZN(n1202) );
  NOR2_X1 U1404 ( .A1(n1315), .A2(n1179), .ZN(n1203) );
  NAND2_X1 U1405 ( .A1(n1214), .A2(n1249), .ZN(n1213) );
  OAI21_X1 U1406 ( .B1(n1380), .B2(n1205), .A(n1204), .ZN(n1968) );
  NAND2_X1 U1407 ( .A1(n1168), .A2(B[17]), .ZN(n1204) );
  INV_X1 U1408 ( .A(IMM[17]), .ZN(n1205) );
  XNOR2_X1 U1409 ( .A(n1540), .B(n1206), .ZN(n1232) );
  INV_X1 U1410 ( .A(n1374), .ZN(n1206) );
  XNOR2_X1 U1411 ( .A(n2099), .B(n1353), .ZN(n1392) );
  NAND2_X1 U1412 ( .A1(S2_IMM_B), .A2(B[3]), .ZN(n1207) );
  INV_X1 U1413 ( .A(IMM[3]), .ZN(n1208) );
  NAND2_X1 U1414 ( .A1(n1293), .A2(n1237), .ZN(n1340) );
  NAND2_X1 U1415 ( .A1(n1676), .A2(n1349), .ZN(n1293) );
  NAND3_X1 U1416 ( .A1(n1128), .A2(n1212), .A3(n1211), .ZN(n2096) );
  NAND3_X1 U1417 ( .A1(n1216), .A2(n1249), .A3(n1735), .ZN(n1211) );
  NAND3_X1 U1418 ( .A1(n1213), .A2(n1215), .A3(n1328), .ZN(n1212) );
  INV_X1 U1419 ( .A(n1229), .ZN(n1214) );
  AOI21_X1 U1420 ( .B1(n1249), .B2(n1182), .A(n1735), .ZN(n1215) );
  NAND4_X1 U1421 ( .A1(n2037), .A2(n2019), .A3(n1985), .A4(n2096), .ZN(n1749)
         );
  NAND2_X1 U1422 ( .A1(n1166), .A2(n1218), .ZN(n1217) );
  AND2_X1 U1423 ( .A1(n1739), .A2(n1740), .ZN(n1218) );
  INV_X1 U1424 ( .A(n1744), .ZN(n1220) );
  NAND2_X1 U1425 ( .A1(n1254), .A2(n1300), .ZN(n1221) );
  NAND2_X1 U1426 ( .A1(n1254), .A2(n1300), .ZN(n1704) );
  AND2_X1 U1427 ( .A1(n1394), .A2(n1661), .ZN(n1485) );
  BUF_X1 U1428 ( .A(n1967), .Z(n1222) );
  BUF_X1 U1429 ( .A(n1579), .Z(n1223) );
  XNOR2_X1 U1430 ( .A(n1305), .B(n1225), .ZN(n1224) );
  XNOR2_X1 U1431 ( .A(n1717), .B(n2235), .ZN(n1225) );
  AND2_X2 U1432 ( .A1(n1559), .A2(n1560), .ZN(n1643) );
  NAND2_X1 U1433 ( .A1(n1347), .A2(n1566), .ZN(n1226) );
  INV_X1 U1434 ( .A(n1230), .ZN(n1227) );
  XOR2_X1 U1435 ( .A(n2072), .B(n1378), .Z(n1228) );
  NAND2_X1 U1436 ( .A1(n1343), .A2(n1344), .ZN(n1229) );
  NAND2_X1 U1437 ( .A1(n1343), .A2(n1344), .ZN(n1697) );
  INV_X1 U1438 ( .A(n1631), .ZN(n1230) );
  OAI21_X1 U1439 ( .B1(n1221), .B2(n1247), .A(n1322), .ZN(n1231) );
  NOR2_X1 U1440 ( .A1(n1550), .A2(n1551), .ZN(n1233) );
  INV_X1 U1441 ( .A(n1440), .ZN(n1234) );
  BUF_X1 U1442 ( .A(n2099), .Z(n1235) );
  INV_X2 U1443 ( .A(n2268), .ZN(n2230) );
  INV_X1 U1444 ( .A(n2234), .ZN(n2170) );
  INV_X1 U1445 ( .A(n2236), .ZN(n2171) );
  INV_X1 U1446 ( .A(n2233), .ZN(n2168) );
  OR2_X1 U1447 ( .A1(n1472), .A2(n1471), .ZN(n1240) );
  INV_X1 U1448 ( .A(n2305), .ZN(n1367) );
  INV_X1 U1449 ( .A(n2306), .ZN(n1370) );
  OR2_X1 U1450 ( .A1(n1975), .A2(n1974), .ZN(n2125) );
  INV_X1 U1451 ( .A(n2186), .ZN(n1356) );
  OR2_X1 U1452 ( .A1(n2025), .A2(n2024), .ZN(n2176) );
  INV_X1 U1453 ( .A(n2115), .ZN(n2276) );
  AND2_X1 U1454 ( .A1(EN_REGN_ALU_OUT), .A2(n1379), .ZN(n2306) );
  AND2_X1 U1455 ( .A1(n1376), .A2(n1477), .ZN(n2232) );
  INV_X1 U1456 ( .A(n2309), .ZN(n1477) );
  INV_X1 U1457 ( .A(n2186), .ZN(n1355) );
  AND3_X1 U1458 ( .A1(n1509), .A2(n1508), .A3(n1507), .ZN(n2322) );
  INV_X1 U1459 ( .A(n2305), .ZN(n1366) );
  INV_X1 U1460 ( .A(n2306), .ZN(n1369) );
  NOR2_X1 U1461 ( .A1(EN_REGN_ALU_OUT), .A2(RST), .ZN(n2305) );
  AND2_X1 U1462 ( .A1(ALU_OPCODE[3]), .A2(n1477), .ZN(n2234) );
  AND2_X1 U1463 ( .A1(ALU_OPCODE[2]), .A2(n1477), .ZN(n2233) );
  AND2_X1 U1464 ( .A1(ALU_OPCODE[1]), .A2(n1477), .ZN(n2236) );
  INV_X1 U1465 ( .A(n2227), .ZN(n1361) );
  INV_X1 U1466 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1377) );
  BUF_X1 U1467 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .Z(n1375) );
  INV_X1 U1468 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1354) );
  AND2_X1 U1469 ( .A1(n1524), .A2(n1523), .ZN(n2323) );
  INV_X1 U1470 ( .A(n2306), .ZN(n1368) );
  AND2_X1 U1471 ( .A1(n1426), .A2(ALU_OPCODE[4]), .ZN(n2115) );
  OR2_X1 U1472 ( .A1(ALU_OPCODE[4]), .A2(ALU_OPCODE[5]), .ZN(n2268) );
  INV_X1 U1473 ( .A(RST), .ZN(n1379) );
  INV_X1 U1474 ( .A(ALU_OPCODE[5]), .ZN(n1426) );
  NOR2_X2 U1475 ( .A1(n1466), .A2(n1465), .ZN(n2199) );
  OAI22_X1 U1476 ( .A1(n2289), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_16/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_16/n5 ) );
  INV_X1 U1477 ( .A(ALUOUT[16]), .ZN(n2289) );
  OAI22_X1 U1478 ( .A1(n2280), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_3/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_3/n5 ) );
  INV_X1 U1479 ( .A(ALUOUT[3]), .ZN(n2280) );
  OAI211_X1 U1480 ( .C1(n2276), .C2(n1818), .A(n1817), .B(n1816), .ZN(
        ALUOUT[3]) );
  OAI21_X1 U1481 ( .B1(n1812), .B2(n1811), .A(n2230), .ZN(n1817) );
  OAI22_X1 U1482 ( .A1(n1855), .A2(n2251), .B1(n2223), .B2(n1810), .ZN(n1811)
         );
  OAI211_X1 U1483 ( .C1(n1868), .C2(n2186), .A(n1809), .B(n1808), .ZN(n1812)
         );
  AOI21_X1 U1484 ( .B1(n1184), .B2(n1823), .A(n1807), .ZN(n1808) );
  OAI211_X1 U1485 ( .C1(n1147), .C2(n2262), .A(n1806), .B(n1805), .ZN(n1807)
         );
  NAND2_X1 U1486 ( .A1(n2260), .A2(n1804), .ZN(n1805) );
  NAND2_X1 U1487 ( .A1(n1362), .A2(n1803), .ZN(n1806) );
  AOI22_X1 U1488 ( .A1(n1358), .A2(n1851), .B1(n1837), .B2(n2173), .ZN(n1809)
         );
  INV_X1 U1489 ( .A(n1802), .ZN(n1818) );
  OAI22_X1 U1490 ( .A1(n2284), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_10/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_10/n5 ) );
  INV_X1 U1491 ( .A(ALUOUT[10]), .ZN(n2284) );
  OAI22_X1 U1492 ( .A1(n2282), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_8/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_8/n5 ) );
  INV_X1 U1493 ( .A(ALUOUT[8]), .ZN(n2282) );
  OAI22_X1 U1494 ( .A1(n2283), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_9/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_9/n5 ) );
  INV_X1 U1495 ( .A(ALUOUT[9]), .ZN(n2283) );
  OAI211_X1 U1496 ( .C1(n1862), .C2(n2276), .A(n1861), .B(n1860), .ZN(
        ALUOUT[9]) );
  OAI21_X1 U1497 ( .B1(n1859), .B2(n1858), .A(n2230), .ZN(n1860) );
  NAND2_X1 U1498 ( .A1(n1857), .A2(n1856), .ZN(n1858) );
  AOI22_X1 U1499 ( .A1(n1184), .A2(n1878), .B1(n1910), .B2(n2173), .ZN(n1856)
         );
  AOI22_X1 U1500 ( .A1(n1358), .A2(n1925), .B1(n1877), .B2(n2260), .ZN(n1857)
         );
  OAI211_X1 U1501 ( .C1(n1855), .C2(n2223), .A(n1854), .B(n1853), .ZN(n1859)
         );
  AOI22_X1 U1502 ( .A1(n1356), .A2(n1976), .B1(n1852), .B2(n1361), .ZN(n1853)
         );
  AOI22_X1 U1503 ( .A1(n2199), .A2(n1958), .B1(n1851), .B2(n2222), .ZN(n1854)
         );
  OAI22_X1 U1504 ( .A1(n2285), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_12/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_12/n5 ) );
  INV_X1 U1505 ( .A(ALUOUT[12]), .ZN(n2285) );
  OAI22_X1 U1506 ( .A1(n2286), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_13/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_13/n5 ) );
  INV_X1 U1507 ( .A(ALUOUT[13]), .ZN(n2286) );
  OAI211_X1 U1508 ( .C1(n1909), .C2(n2268), .A(n1908), .B(n1907), .ZN(
        ALUOUT[13]) );
  NOR3_X1 U1509 ( .A1(n1901), .A2(n1900), .A3(n1899), .ZN(n1909) );
  OAI22_X1 U1510 ( .A1(n1913), .A2(n2186), .B1(n1898), .B2(n2262), .ZN(n1899)
         );
  OAI22_X1 U1511 ( .A1(n1896), .A2(n1357), .B1(n1895), .B2(n1240), .ZN(n1900)
         );
  INV_X1 U1512 ( .A(n1958), .ZN(n1895) );
  INV_X1 U1513 ( .A(n2009), .ZN(n1896) );
  OAI211_X1 U1514 ( .C1(n1894), .C2(n2251), .A(n1893), .B(n1892), .ZN(n1901)
         );
  AOI22_X1 U1515 ( .A1(n1360), .A2(n1910), .B1(n1925), .B2(n1361), .ZN(n1892)
         );
  AOI22_X1 U1516 ( .A1(n2173), .A2(n1991), .B1(n1976), .B2(n2260), .ZN(n1893)
         );
  INV_X1 U1517 ( .A(n2026), .ZN(n1894) );
  OAI22_X1 U1518 ( .A1(n2287), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_14/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_14/n5 ) );
  INV_X1 U1519 ( .A(ALUOUT[14]), .ZN(n2287) );
  OAI22_X1 U1520 ( .A1(n2290), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_17/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_17/n5 ) );
  INV_X1 U1521 ( .A(ALUOUT[17]), .ZN(n2290) );
  OAI211_X1 U1522 ( .C1(n1985), .C2(n2276), .A(n1984), .B(n1983), .ZN(
        ALUOUT[17]) );
  OAI21_X1 U1523 ( .B1(n1982), .B2(n1981), .A(n2230), .ZN(n1983) );
  NAND2_X1 U1524 ( .A1(n1980), .A2(n1979), .ZN(n1981) );
  AOI22_X1 U1525 ( .A1(n1358), .A2(n2087), .B1(n2043), .B2(n2260), .ZN(n1979)
         );
  AOI22_X1 U1526 ( .A1(n1184), .A2(n2026), .B1(n2067), .B2(n2173), .ZN(n1980)
         );
  OAI211_X1 U1527 ( .C1(n2058), .C2(n2251), .A(n1978), .B(n1977), .ZN(n1982)
         );
  AOI22_X1 U1528 ( .A1(n1361), .A2(n2009), .B1(n1976), .B2(n2222), .ZN(n1977)
         );
  AOI22_X1 U1529 ( .A1(n2125), .A2(n1355), .B1(n1991), .B2(n1359), .ZN(n1978)
         );
  OAI22_X1 U1530 ( .A1(n2288), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_15/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_15/n5 ) );
  INV_X1 U1531 ( .A(ALUOUT[15]), .ZN(n2288) );
  OAI211_X1 U1532 ( .C1(n1943), .C2(n2276), .A(n1942), .B(n1941), .ZN(
        ALUOUT[15]) );
  OAI21_X1 U1533 ( .B1(n1937), .B2(n1936), .A(n2230), .ZN(n1942) );
  NAND2_X1 U1534 ( .A1(n1935), .A2(n1934), .ZN(n1936) );
  AOI22_X1 U1535 ( .A1(n1356), .A2(n2087), .B1(n2043), .B2(n1358), .ZN(n1934)
         );
  AOI22_X1 U1536 ( .A1(n1184), .A2(n1991), .B1(n2026), .B2(n2173), .ZN(n1935)
         );
  OAI211_X1 U1537 ( .C1(n1928), .C2(n2251), .A(n1927), .B(n1926), .ZN(n1937)
         );
  AOI22_X1 U1538 ( .A1(n1360), .A2(n1958), .B1(n1925), .B2(n2222), .ZN(n1926)
         );
  AOI22_X1 U1539 ( .A1(n1362), .A2(n1976), .B1(n2009), .B2(n2260), .ZN(n1927)
         );
  INV_X1 U1540 ( .A(n2067), .ZN(n1928) );
  OAI22_X1 U1541 ( .A1(n2279), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_2/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_2/n5 ) );
  INV_X1 U1542 ( .A(ALUOUT[2]), .ZN(n2279) );
  OAI211_X1 U1543 ( .C1(n2276), .C2(n1801), .A(n1800), .B(n1799), .ZN(
        ALUOUT[2]) );
  OAI21_X1 U1544 ( .B1(n1795), .B2(n1794), .A(n2230), .ZN(n1800) );
  OAI21_X1 U1545 ( .B1(n1840), .B2(n2251), .A(n1793), .ZN(n1794) );
  OAI211_X1 U1546 ( .C1(n1820), .C2(n2255), .A(n1792), .B(n1791), .ZN(n1795)
         );
  AOI22_X1 U1547 ( .A1(n1356), .A2(n1869), .B1(n1837), .B2(n1358), .ZN(n1791)
         );
  AOI21_X1 U1548 ( .B1(n1184), .B2(n1803), .A(n1790), .ZN(n1792) );
  OAI21_X1 U1549 ( .B1(n2227), .B2(n1810), .A(n1789), .ZN(n1790) );
  AOI22_X1 U1550 ( .A1(n2222), .A2(n1788), .B1(n1823), .B2(n2260), .ZN(n1789)
         );
  OAI22_X1 U1551 ( .A1(n2293), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_20/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_20/n5 ) );
  INV_X1 U1552 ( .A(ALUOUT[20]), .ZN(n2293) );
  OAI22_X1 U1553 ( .A1(n2303), .A2(n1369), .B1(\COMP_REGN_ALUOUT/ffi_30/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_30/n5 ) );
  INV_X1 U1554 ( .A(ALUOUT[30]), .ZN(n2303) );
  OAI22_X1 U1555 ( .A1(n2292), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_19/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_19/n5 ) );
  INV_X1 U1556 ( .A(ALUOUT[19]), .ZN(n2292) );
  OAI211_X1 U1557 ( .C1(n2019), .C2(n2276), .A(n2018), .B(n2017), .ZN(
        ALUOUT[19]) );
  OAI21_X1 U1558 ( .B1(n2013), .B2(n2012), .A(n2230), .ZN(n2018) );
  OAI211_X1 U1559 ( .C1(n2110), .C2(n2251), .A(n2011), .B(n2010), .ZN(n2012)
         );
  AOI22_X1 U1560 ( .A1(n1184), .A2(n2067), .B1(n2009), .B2(n2222), .ZN(n2010)
         );
  AOI22_X1 U1561 ( .A1(n1355), .A2(n2154), .B1(n2125), .B2(n1358), .ZN(n2011)
         );
  NAND2_X1 U1562 ( .A1(n2003), .A2(n2002), .ZN(n2013) );
  AOI22_X1 U1563 ( .A1(n1361), .A2(n2043), .B1(n2087), .B2(n2260), .ZN(n2002)
         );
  AOI22_X1 U1564 ( .A1(n2097), .A2(n2173), .B1(n1360), .B2(n2026), .ZN(n2003)
         );
  OAI22_X1 U1565 ( .A1(n2295), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_22/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_22/n5 ) );
  INV_X1 U1566 ( .A(ALUOUT[22]), .ZN(n2295) );
  OAI21_X1 U1567 ( .B1(n1964), .B2(n1963), .A(n2230), .ZN(n1965) );
  NAND2_X1 U1568 ( .A1(n1962), .A2(n1961), .ZN(n1963) );
  AOI22_X1 U1569 ( .A1(n1358), .A2(n2067), .B1(n2026), .B2(n2260), .ZN(n1961)
         );
  AOI22_X1 U1570 ( .A1(n1184), .A2(n2009), .B1(n2043), .B2(n2173), .ZN(n1962)
         );
  OAI211_X1 U1571 ( .C1(n2058), .C2(n2186), .A(n1960), .B(n1959), .ZN(n1964)
         );
  AOI22_X1 U1572 ( .A1(n1362), .A2(n1991), .B1(n1958), .B2(n2222), .ZN(n1959)
         );
  AOI22_X1 U1573 ( .A1(n1360), .A2(n1976), .B1(n2087), .B2(n2199), .ZN(n1960)
         );
  INV_X1 U1574 ( .A(n2322), .ZN(ALUOUT[4]) );
  OAI21_X1 U1575 ( .B1(n1506), .B2(n1505), .A(n2230), .ZN(n1507) );
  NAND4_X1 U1576 ( .A1(n1504), .A2(n1503), .A3(n1502), .A4(n1501), .ZN(n1505)
         );
  NAND2_X1 U1577 ( .A1(n1184), .A2(n1804), .ZN(n1501) );
  NAND2_X1 U1578 ( .A1(n1360), .A2(n1803), .ZN(n1502) );
  AOI22_X1 U1579 ( .A1(n2222), .A2(n1777), .B1(n1362), .B2(n1823), .ZN(n1503)
         );
  NAND2_X1 U1580 ( .A1(n1878), .A2(n1355), .ZN(n1504) );
  NAND4_X1 U1581 ( .A1(n1500), .A2(n1499), .A3(n1498), .A4(n1497), .ZN(n1506)
         );
  NAND2_X1 U1582 ( .A1(n1851), .A2(n2173), .ZN(n1497) );
  NAND2_X1 U1583 ( .A1(n1852), .A2(n2199), .ZN(n1498) );
  NAND2_X1 U1584 ( .A1(n1869), .A2(n1358), .ZN(n1499) );
  NAND2_X1 U1585 ( .A1(n1837), .A2(n2260), .ZN(n1500) );
  INV_X1 U1586 ( .A(n1489), .ZN(n1490) );
  OAI211_X1 U1587 ( .C1(n1189), .C2(n2276), .A(n1846), .B(n1845), .ZN(
        ALUOUT[8]) );
  OAI21_X1 U1588 ( .B1(n1844), .B2(n1843), .A(n2230), .ZN(n1845) );
  NAND2_X1 U1589 ( .A1(n1842), .A2(n1841), .ZN(n1843) );
  AOI22_X1 U1590 ( .A1(n1362), .A2(n1869), .B1(n1878), .B2(n2260), .ZN(n1841)
         );
  AOI22_X1 U1591 ( .A1(n1184), .A2(n1852), .B1(n1910), .B2(n1358), .ZN(n1842)
         );
  OAI211_X1 U1592 ( .C1(n1840), .C2(n2223), .A(n1839), .B(n1838), .ZN(n1844)
         );
  AOI22_X1 U1593 ( .A1(n1356), .A2(n1958), .B1(n1877), .B2(n2173), .ZN(n1838)
         );
  AOI22_X1 U1594 ( .A1(n2199), .A2(n1925), .B1(n1837), .B2(n2222), .ZN(n1839)
         );
  OAI211_X1 U1595 ( .C1(n1876), .C2(n2276), .A(n1875), .B(n1874), .ZN(
        ALUOUT[10]) );
  OAI21_X1 U1596 ( .B1(n1873), .B2(n1872), .A(n2230), .ZN(n1874) );
  NAND2_X1 U1597 ( .A1(n1871), .A2(n1870), .ZN(n1872) );
  AOI22_X1 U1598 ( .A1(n2222), .A2(n1869), .B1(n1910), .B2(n2260), .ZN(n1870)
         );
  AOI22_X1 U1599 ( .A1(n1184), .A2(n1877), .B1(n1925), .B2(n2173), .ZN(n1871)
         );
  OAI211_X1 U1600 ( .C1(n1868), .C2(n2223), .A(n1867), .B(n1866), .ZN(n1873)
         );
  AOI22_X1 U1601 ( .A1(n2199), .A2(n1976), .B1(n1878), .B2(n1361), .ZN(n1866)
         );
  AOI22_X1 U1602 ( .A1(n1356), .A2(n1991), .B1(n1958), .B2(n1358), .ZN(n1867)
         );
  OAI211_X1 U1603 ( .C1(n1891), .C2(n2276), .A(n1890), .B(n1889), .ZN(
        ALUOUT[12]) );
  OAI21_X1 U1604 ( .B1(n1884), .B2(n1883), .A(n2230), .ZN(n1890) );
  NAND2_X1 U1605 ( .A1(n1882), .A2(n1881), .ZN(n1883) );
  AOI22_X1 U1606 ( .A1(n1362), .A2(n1910), .B1(n1925), .B2(n1184), .ZN(n1881)
         );
  AOI22_X1 U1607 ( .A1(n1356), .A2(n2026), .B1(n1958), .B2(n2260), .ZN(n1882)
         );
  OAI211_X1 U1608 ( .C1(n1898), .C2(n2223), .A(n1880), .B(n1879), .ZN(n1884)
         );
  AOI22_X1 U1609 ( .A1(n2199), .A2(n2009), .B1(n1878), .B2(n2222), .ZN(n1879)
         );
  AOI22_X1 U1610 ( .A1(n2173), .A2(n1976), .B1(n1991), .B2(n1358), .ZN(n1880)
         );
  INV_X1 U1611 ( .A(n1877), .ZN(n1898) );
  OAI22_X1 U1612 ( .A1(n2299), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_26/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_26/n5 ) );
  INV_X1 U1613 ( .A(ALUOUT[26]), .ZN(n2299) );
  OAI22_X1 U1614 ( .A1(n2291), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_18/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_18/n5 ) );
  INV_X1 U1615 ( .A(ALUOUT[18]), .ZN(n2291) );
  OAI211_X1 U1616 ( .C1(n1924), .C2(n2276), .A(n1923), .B(n1922), .ZN(
        ALUOUT[14]) );
  OAI21_X1 U1617 ( .B1(n1918), .B2(n1917), .A(n2230), .ZN(n1923) );
  NAND2_X1 U1618 ( .A1(n1916), .A2(n1915), .ZN(n1917) );
  AOI22_X1 U1619 ( .A1(n1356), .A2(n2067), .B1(n2026), .B2(n1358), .ZN(n1915)
         );
  AOI22_X1 U1620 ( .A1(n1184), .A2(n1976), .B1(n2009), .B2(n2173), .ZN(n1916)
         );
  OAI211_X1 U1621 ( .C1(n1913), .C2(n2251), .A(n1912), .B(n1911), .ZN(n1918)
         );
  AOI22_X1 U1622 ( .A1(n1360), .A2(n1925), .B1(n1910), .B2(n2222), .ZN(n1911)
         );
  AOI22_X1 U1623 ( .A1(n1362), .A2(n1958), .B1(n1991), .B2(n2260), .ZN(n1912)
         );
  INV_X1 U1624 ( .A(n2043), .ZN(n1913) );
  OAI22_X1 U1625 ( .A1(n2297), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_24/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_24/n5 ) );
  INV_X1 U1626 ( .A(ALUOUT[24]), .ZN(n2297) );
  OAI22_X1 U1627 ( .A1(n2294), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_21/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_21/n5 ) );
  INV_X1 U1628 ( .A(ALUOUT[21]), .ZN(n2294) );
  OAI211_X1 U1629 ( .C1(n2055), .C2(n2276), .A(n2054), .B(n2053), .ZN(
        ALUOUT[21]) );
  OAI21_X1 U1630 ( .B1(n2049), .B2(n2048), .A(n2230), .ZN(n2054) );
  NAND2_X1 U1631 ( .A1(n2047), .A2(n2046), .ZN(n2048) );
  AOI22_X1 U1632 ( .A1(n2173), .A2(n1040), .B1(n2125), .B2(n2260), .ZN(n2046)
         );
  AOI22_X1 U1633 ( .A1(n2097), .A2(n1184), .B1(n1360), .B2(n2067), .ZN(n2047)
         );
  OAI211_X1 U1634 ( .C1(n2112), .C2(n2251), .A(n2045), .B(n2044), .ZN(n2049)
         );
  AOI22_X1 U1635 ( .A1(n1361), .A2(n2087), .B1(n2043), .B2(n2222), .ZN(n2044)
         );
  AOI22_X1 U1636 ( .A1(n2177), .A2(n1355), .B1(n1358), .B2(n2154), .ZN(n2045)
         );
  OAI22_X1 U1637 ( .A1(n2298), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_25/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_25/n5 ) );
  INV_X1 U1638 ( .A(ALUOUT[25]), .ZN(n2298) );
  OAI22_X1 U1639 ( .A1(n2301), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_28/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_28/n5 ) );
  INV_X1 U1640 ( .A(ALUOUT[28]), .ZN(n2301) );
  INV_X1 U1641 ( .A(n2321), .ZN(ALUOUT[11]) );
  AOI21_X1 U1642 ( .B1(n1693), .B2(n2115), .A(n1483), .ZN(n2321) );
  NAND2_X1 U1643 ( .A1(n1482), .A2(n1481), .ZN(n1483) );
  NAND2_X1 U1644 ( .A1(n1476), .A2(n2230), .ZN(n1482) );
  NAND4_X1 U1645 ( .A1(n1243), .A2(n1475), .A3(n1474), .A4(n1473), .ZN(n1476)
         );
  AOI22_X1 U1646 ( .A1(n2199), .A2(n1991), .B1(n1910), .B2(n1184), .ZN(n1473)
         );
  AOI22_X1 U1647 ( .A1(n2222), .A2(n1852), .B1(n1925), .B2(n2260), .ZN(n1474)
         );
  AOI22_X1 U1648 ( .A1(n1356), .A2(n2009), .B1(n1877), .B2(n1361), .ZN(n1475)
         );
  NAND2_X1 U1649 ( .A1(n1878), .A2(n1359), .ZN(n1447) );
  NAND2_X1 U1650 ( .A1(n1976), .A2(n1358), .ZN(n1448) );
  OAI211_X1 U1651 ( .C1(n1363), .C2(n2124), .A(n1439), .B(n1438), .ZN(n1976)
         );
  NOR2_X1 U1652 ( .A1(n1930), .A2(n1437), .ZN(n1439) );
  NAND2_X1 U1653 ( .A1(n1958), .A2(n2173), .ZN(n1449) );
  OAI211_X1 U1654 ( .C1(n1363), .C2(n2105), .A(n1432), .B(n1431), .ZN(n1958)
         );
  NAND2_X1 U1655 ( .A1(n2210), .A2(n1760), .ZN(n1431) );
  NOR2_X1 U1656 ( .A1(n1930), .A2(n1430), .ZN(n1432) );
  OAI22_X1 U1657 ( .A1(n2302), .A2(n1369), .B1(\COMP_REGN_ALUOUT/ffi_29/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_29/n5 ) );
  INV_X1 U1658 ( .A(ALUOUT[29]), .ZN(n2302) );
  OAI22_X1 U1659 ( .A1(n2281), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_5/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_5/n5 ) );
  INV_X1 U1660 ( .A(ALUOUT[5]), .ZN(n2281) );
  OAI21_X1 U1661 ( .B1(n1833), .B2(n2276), .A(n1832), .ZN(ALUOUT[5]) );
  AOI21_X1 U1662 ( .B1(n1831), .B2(n2230), .A(n1830), .ZN(n1832) );
  AOI22_X1 U1663 ( .A1(n1878), .A2(n2199), .B1(n1360), .B2(n1823), .ZN(n1824)
         );
  AOI22_X1 U1664 ( .A1(n1184), .A2(n1837), .B1(n1851), .B2(n2260), .ZN(n1825)
         );
  AOI211_X1 U1665 ( .C1(n1355), .C2(n1877), .A(n1822), .B(n1821), .ZN(n1826)
         );
  OAI22_X1 U1666 ( .A1(n1855), .A2(n2255), .B1(n1868), .B2(n1357), .ZN(n1821)
         );
  INV_X1 U1667 ( .A(n1852), .ZN(n1868) );
  INV_X1 U1668 ( .A(n1869), .ZN(n1855) );
  OAI22_X1 U1669 ( .A1(n2227), .A2(n1820), .B1(n1819), .B2(n2262), .ZN(n1822)
         );
  OAI22_X1 U1670 ( .A1(n2278), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_1/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_1/n5 ) );
  INV_X1 U1671 ( .A(ALUOUT[1]), .ZN(n2278) );
  OAI211_X1 U1672 ( .C1(n2276), .C2(n1787), .A(n1786), .B(n1785), .ZN(
        ALUOUT[1]) );
  NAND2_X1 U1673 ( .A1(n1780), .A2(n2230), .ZN(n1786) );
  AOI211_X1 U1674 ( .C1(n1184), .C2(n1777), .A(n1776), .B(n1775), .ZN(n1778)
         );
  OAI22_X1 U1675 ( .A1(n1774), .A2(n2251), .B1(n1840), .B2(n2186), .ZN(n1775)
         );
  INV_X1 U1676 ( .A(n1851), .ZN(n1840) );
  INV_X1 U1677 ( .A(n1837), .ZN(n1774) );
  OAI21_X1 U1678 ( .B1(n2255), .B2(n1773), .A(n1772), .ZN(n1776) );
  AOI22_X1 U1679 ( .A1(n1358), .A2(n1804), .B1(n2260), .B2(n1803), .ZN(n1772)
         );
  INV_X1 U1680 ( .A(n1819), .ZN(n1803) );
  INV_X1 U1681 ( .A(n1810), .ZN(n1777) );
  OAI211_X1 U1682 ( .C1(n2264), .C2(n2186), .A(n2201), .B(n2200), .ZN(n2203)
         );
  NAND2_X1 U1683 ( .A1(n2253), .A2(n2199), .ZN(n2200) );
  NAND2_X1 U1684 ( .A1(n2221), .A2(n1359), .ZN(n2201) );
  OAI22_X1 U1685 ( .A1(n2296), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_23/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_23/n5 ) );
  INV_X1 U1686 ( .A(ALUOUT[23]), .ZN(n2296) );
  OAI211_X1 U1687 ( .C1(n2096), .C2(n2276), .A(n2095), .B(n2094), .ZN(
        ALUOUT[23]) );
  OAI21_X1 U1688 ( .B1(n2093), .B2(n2092), .A(n2230), .ZN(n2094) );
  NAND2_X1 U1689 ( .A1(n2091), .A2(n2090), .ZN(n2092) );
  AOI22_X1 U1690 ( .A1(n2173), .A2(n2176), .B1(n2154), .B2(n2260), .ZN(n2090)
         );
  AOI22_X1 U1691 ( .A1(n1361), .A2(n2125), .B1(n1040), .B2(n1184), .ZN(n2091)
         );
  OAI211_X1 U1692 ( .C1(n2157), .C2(n2251), .A(n2089), .B(n2088), .ZN(n2093)
         );
  AOI22_X1 U1693 ( .A1(n2097), .A2(n1359), .B1(n2222), .B2(n2087), .ZN(n2088)
         );
  AOI22_X1 U1694 ( .A1(n1356), .A2(n2224), .B1(n2177), .B2(n1358), .ZN(n2089)
         );
  OAI22_X1 U1695 ( .A1(n2304), .A2(n1369), .B1(\COMP_REGN_ALUOUT/ffi_31/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_31/n5 ) );
  INV_X1 U1696 ( .A(ALUOUT[31]), .ZN(n2304) );
  OAI211_X1 U1697 ( .C1(n2037), .C2(n2276), .A(n2036), .B(n2035), .ZN(
        ALUOUT[20]) );
  OAI21_X1 U1698 ( .B1(n2030), .B2(n2029), .A(n2230), .ZN(n2036) );
  OAI211_X1 U1699 ( .C1(n2111), .C2(n2251), .A(n2028), .B(n2027), .ZN(n2029)
         );
  AOI22_X1 U1700 ( .A1(n1184), .A2(n2087), .B1(n2026), .B2(n2222), .ZN(n2027)
         );
  AOI22_X1 U1701 ( .A1(n1355), .A2(n2176), .B1(n2135), .B2(n1358), .ZN(n2028)
         );
  NAND2_X1 U1702 ( .A1(n2021), .A2(n2020), .ZN(n2030) );
  AOI22_X1 U1703 ( .A1(n1359), .A2(n2043), .B1(n2067), .B2(n1361), .ZN(n2020)
         );
  AOI22_X1 U1704 ( .A1(n2097), .A2(n2260), .B1(n2173), .B2(n2125), .ZN(n2021)
         );
  INV_X1 U1705 ( .A(n2323), .ZN(ALUOUT[6]) );
  AOI21_X1 U1706 ( .B1(n1522), .B2(n2230), .A(n1521), .ZN(n1523) );
  NAND4_X1 U1707 ( .A1(n1517), .A2(n1516), .A3(n1515), .A4(n1514), .ZN(n1522)
         );
  AOI22_X1 U1708 ( .A1(n1184), .A2(n1851), .B1(n1877), .B2(n2199), .ZN(n1514)
         );
  AOI22_X1 U1709 ( .A1(n1362), .A2(n1837), .B1(n1869), .B2(n2260), .ZN(n1515)
         );
  AOI22_X1 U1710 ( .A1(n1356), .A2(n1910), .B1(n1878), .B2(n1358), .ZN(n1516)
         );
  INV_X1 U1711 ( .A(n1823), .ZN(n1773) );
  OR2_X1 U1712 ( .A1(n1667), .A2(n2276), .ZN(n1524) );
  OAI22_X1 U1713 ( .A1(n2261), .A2(n2217), .B1(n2216), .B2(n2255), .ZN(n2218)
         );
  OAI22_X1 U1714 ( .A1(n2264), .A2(n2251), .B1(n2252), .B2(n2186), .ZN(n2219)
         );
  OAI211_X1 U1715 ( .C1(n2077), .C2(n2276), .A(n2076), .B(n2075), .ZN(
        ALUOUT[22]) );
  OAI21_X1 U1716 ( .B1(n2071), .B2(n2070), .A(n2230), .ZN(n2076) );
  OAI211_X1 U1717 ( .C1(n2202), .C2(n2251), .A(n2069), .B(n2068), .ZN(n2070)
         );
  AOI22_X1 U1718 ( .A1(n1359), .A2(n2087), .B1(n2067), .B2(n2222), .ZN(n2068)
         );
  AOI22_X1 U1719 ( .A1(n1358), .A2(n2176), .B1(n2221), .B2(n1355), .ZN(n2069)
         );
  OAI211_X1 U1720 ( .C1(n2058), .C2(n2227), .A(n2057), .B(n2056), .ZN(n2071)
         );
  NAND2_X1 U1721 ( .A1(n2125), .A2(n1184), .ZN(n2056) );
  AOI22_X1 U1722 ( .A1(n2173), .A2(n2154), .B1(n2135), .B2(n2260), .ZN(n2057)
         );
  OAI211_X1 U1723 ( .C1(n2144), .C2(n2276), .A(n2143), .B(n2142), .ZN(
        ALUOUT[26]) );
  OAI21_X1 U1724 ( .B1(n2141), .B2(n2140), .A(n2230), .ZN(n2142) );
  NAND2_X1 U1725 ( .A1(n2139), .A2(n2138), .ZN(n2140) );
  AOI22_X1 U1726 ( .A1(n2224), .A2(n2173), .B1(n2260), .B2(n2221), .ZN(n2138)
         );
  AOI22_X1 U1727 ( .A1(n2177), .A2(n1184), .B1(n1362), .B2(n2176), .ZN(n2139)
         );
  OAI211_X1 U1728 ( .C1(n2254), .C2(n2251), .A(n2137), .B(n2136), .ZN(n2141)
         );
  AOI22_X1 U1729 ( .A1(n1360), .A2(n2154), .B1(n2135), .B2(n2222), .ZN(n2136)
         );
  AOI22_X1 U1730 ( .A1(n1355), .A2(n2187), .B1(n2226), .B2(n1358), .ZN(n2137)
         );
  INV_X1 U1731 ( .A(n2324), .ZN(ALUOUT[7]) );
  AOI21_X1 U1732 ( .B1(n1668), .B2(n2115), .A(n1545), .ZN(n2324) );
  NAND2_X1 U1733 ( .A1(n1544), .A2(n1543), .ZN(n1545) );
  NAND2_X1 U1734 ( .A1(n1539), .A2(n2230), .ZN(n1544) );
  NAND4_X1 U1735 ( .A1(n1538), .A2(n1537), .A3(n1536), .A4(n1535), .ZN(n1539)
         );
  AOI22_X1 U1736 ( .A1(n1362), .A2(n1851), .B1(n1910), .B2(n2199), .ZN(n1535)
         );
  OAI211_X1 U1737 ( .C1(n2207), .C2(n1363), .A(n1496), .B(n1470), .ZN(n1910)
         );
  NAND2_X1 U1738 ( .A1(n1494), .A2(n2059), .ZN(n1470) );
  OAI211_X1 U1739 ( .C1(n2121), .C2(n2244), .A(n1496), .B(n1495), .ZN(n1851)
         );
  NAND2_X1 U1740 ( .A1(n1494), .A2(n1971), .ZN(n1495) );
  AOI22_X1 U1741 ( .A1(n1184), .A2(n1869), .B1(n1878), .B2(n2173), .ZN(n1536)
         );
  OAI211_X1 U1742 ( .C1(n2182), .C2(n1363), .A(n1496), .B(n1444), .ZN(n1878)
         );
  NAND2_X1 U1743 ( .A1(n1494), .A2(n2179), .ZN(n1444) );
  OAI211_X1 U1744 ( .C1(n2131), .C2(n2244), .A(n1496), .B(n1493), .ZN(n1869)
         );
  NAND2_X1 U1745 ( .A1(n1494), .A2(n1989), .ZN(n1493) );
  AOI22_X1 U1746 ( .A1(n1356), .A2(n1925), .B1(n1877), .B2(n1358), .ZN(n1537)
         );
  OAI211_X1 U1747 ( .C1(n2192), .C2(n1363), .A(n1496), .B(n1453), .ZN(n1877)
         );
  NAND2_X1 U1748 ( .A1(n1494), .A2(n2038), .ZN(n1453) );
  OAI211_X1 U1749 ( .C1(n2240), .C2(n1363), .A(n1496), .B(n1461), .ZN(n1925)
         );
  NAND2_X1 U1750 ( .A1(n1494), .A2(n2081), .ZN(n1461) );
  INV_X1 U1751 ( .A(n1534), .ZN(n1538) );
  OAI211_X1 U1752 ( .C1(n2262), .C2(n1820), .A(n1533), .B(n1532), .ZN(n1534)
         );
  NAND2_X1 U1753 ( .A1(n1852), .A2(n2260), .ZN(n1532) );
  OAI211_X1 U1754 ( .C1(n1363), .C2(n1147), .A(n1458), .B(n1496), .ZN(n1852)
         );
  NAND2_X1 U1755 ( .A1(n1494), .A2(n2004), .ZN(n1458) );
  NAND2_X1 U1756 ( .A1(n1837), .A2(n1359), .ZN(n1533) );
  INV_X1 U1757 ( .A(n1804), .ZN(n1820) );
  OAI211_X1 U1758 ( .C1(n2001), .C2(n2276), .A(n2000), .B(n1999), .ZN(
        ALUOUT[18]) );
  OAI21_X1 U1759 ( .B1(n1998), .B2(n1997), .A(n2230), .ZN(n1999) );
  NAND2_X1 U1760 ( .A1(n1996), .A2(n1995), .ZN(n1997) );
  AOI22_X1 U1761 ( .A1(n1360), .A2(n2009), .B1(n2067), .B2(n2260), .ZN(n1995)
         );
  OAI211_X1 U1762 ( .C1(n1363), .C2(n1325), .A(n1452), .B(n1451), .ZN(n2009)
         );
  NAND2_X1 U1763 ( .A1(n2210), .A2(n1813), .ZN(n1451) );
  NOR2_X1 U1764 ( .A1(n1930), .A2(n1450), .ZN(n1452) );
  AOI22_X1 U1765 ( .A1(n1361), .A2(n2026), .B1(n2087), .B2(n2173), .ZN(n1996)
         );
  OAI211_X1 U1766 ( .C1(n2244), .C2(n2246), .A(n1933), .B(n1932), .ZN(n2087)
         );
  NAND2_X1 U1767 ( .A1(n2210), .A2(n1931), .ZN(n1932) );
  NOR2_X1 U1768 ( .A1(n1930), .A2(n1929), .ZN(n1933) );
  OAI211_X1 U1769 ( .C1(n1994), .C2(n2251), .A(n1993), .B(n1992), .ZN(n1998)
         );
  AOI22_X1 U1770 ( .A1(n1184), .A2(n2043), .B1(n1991), .B2(n2222), .ZN(n1992)
         );
  OAI211_X1 U1771 ( .C1(n1363), .C2(n2134), .A(n1469), .B(n1468), .ZN(n1991)
         );
  NAND2_X1 U1772 ( .A1(n2210), .A2(n1788), .ZN(n1468) );
  NOR2_X1 U1773 ( .A1(n1930), .A2(n1467), .ZN(n1469) );
  NOR2_X1 U1774 ( .A1(n2211), .A2(n1352), .ZN(n1930) );
  AOI22_X1 U1775 ( .A1(n2097), .A2(n1358), .B1(n1356), .B2(n2135), .ZN(n1993)
         );
  INV_X1 U1776 ( .A(n2125), .ZN(n1994) );
  OAI22_X1 U1777 ( .A1(n2112), .A2(n2217), .B1(n2202), .B2(n2255), .ZN(n2113)
         );
  INV_X1 U1778 ( .A(n2176), .ZN(n2112) );
  INV_X1 U1779 ( .A(n2135), .ZN(n2110) );
  INV_X1 U1780 ( .A(n2154), .ZN(n2111) );
  OAI211_X1 U1781 ( .C1(n2263), .C2(n2251), .A(n2109), .B(n2108), .ZN(n2114)
         );
  AOI22_X1 U1782 ( .A1(n2226), .A2(n1355), .B1(n1358), .B2(n2221), .ZN(n2108)
         );
  INV_X1 U1783 ( .A(n2265), .ZN(n2226) );
  AOI22_X1 U1784 ( .A1(n2097), .A2(n2222), .B1(n1360), .B2(n2125), .ZN(n2109)
         );
  OAI22_X1 U1785 ( .A1(n1973), .A2(n1363), .B1(n2245), .B2(n2121), .ZN(n1974)
         );
  INV_X1 U1786 ( .A(n2123), .ZN(n1973) );
  OAI211_X1 U1787 ( .C1(n2084), .C2(n2122), .A(n2083), .B(n1972), .ZN(n1975)
         );
  NAND2_X1 U1788 ( .A1(n2210), .A2(n1971), .ZN(n1972) );
  INV_X1 U1789 ( .A(n2058), .ZN(n2097) );
  NOR2_X1 U1790 ( .A1(n1957), .A2(n1956), .ZN(n2058) );
  OAI22_X1 U1791 ( .A1(n1955), .A2(n1363), .B1(n2245), .B2(n2101), .ZN(n1956)
         );
  OAI211_X1 U1792 ( .C1(n2084), .C2(n2102), .A(n2083), .B(n1952), .ZN(n1957)
         );
  NAND2_X1 U1793 ( .A1(n2210), .A2(n1951), .ZN(n1952) );
  OAI211_X1 U1794 ( .C1(n2216), .C2(n2251), .A(n2189), .B(n2188), .ZN(n2190)
         );
  AOI22_X1 U1795 ( .A1(n2187), .A2(n1358), .B1(n1356), .B2(n2253), .ZN(n2188)
         );
  INV_X1 U1796 ( .A(n2261), .ZN(n2187) );
  AOI22_X1 U1797 ( .A1(n2177), .A2(n1359), .B1(n2222), .B2(n2176), .ZN(n2189)
         );
  INV_X1 U1798 ( .A(n2202), .ZN(n2177) );
  NAND2_X1 U1799 ( .A1(n2225), .A2(n2173), .ZN(n2174) );
  AOI22_X1 U1800 ( .A1(n2224), .A2(n1184), .B1(n1362), .B2(n2221), .ZN(n2175)
         );
  INV_X1 U1801 ( .A(n2263), .ZN(n2224) );
  OAI21_X1 U1802 ( .B1(n1224), .B2(n2276), .A(n2275), .ZN(ALUOUT[31]) );
  AOI211_X1 U1803 ( .C1(n2274), .C2(n2273), .A(n2272), .B(n2271), .ZN(n2275)
         );
  AOI21_X1 U1804 ( .B1(n2270), .B2(n2269), .A(n2268), .ZN(n2271) );
  NOR2_X1 U1805 ( .A1(n2267), .A2(n2266), .ZN(n2269) );
  OAI22_X1 U1806 ( .A1(n2265), .A2(n2223), .B1(n2264), .B2(n1357), .ZN(n2266)
         );
  INV_X1 U1807 ( .A(n2220), .ZN(n1357) );
  NOR2_X1 U1808 ( .A1(n2198), .A2(n2197), .ZN(n2264) );
  OAI211_X1 U1809 ( .C1(n1363), .C2(n2196), .A(n2195), .B(n2211), .ZN(n2197)
         );
  NAND2_X1 U1810 ( .A1(n2210), .A2(n2194), .ZN(n2195) );
  OAI22_X1 U1811 ( .A1(n2245), .A2(n2193), .B1(n2239), .B2(n2192), .ZN(n2198)
         );
  OAI22_X1 U1812 ( .A1(n2263), .A2(n2262), .B1(n2261), .B2(n1240), .ZN(n2267)
         );
  AOI211_X1 U1813 ( .C1(n2260), .C2(n2259), .A(n2258), .B(n2257), .ZN(n2270)
         );
  OAI22_X1 U1814 ( .A1(n2256), .A2(n2255), .B1(n2254), .B2(n2227), .ZN(n2257)
         );
  INV_X1 U1815 ( .A(n2253), .ZN(n2256) );
  NAND4_X1 U1816 ( .A1(n2185), .A2(n2184), .A3(n1239), .A4(n2183), .ZN(n2253)
         );
  OR2_X1 U1817 ( .A1(n2239), .A2(n2182), .ZN(n2183) );
  NAND2_X1 U1818 ( .A1(n2180), .A2(n2179), .ZN(n2184) );
  NAND2_X1 U1819 ( .A1(n1364), .A2(n2178), .ZN(n2185) );
  OAI22_X1 U1820 ( .A1(n2252), .A2(n2251), .B1(n2250), .B2(n2249), .ZN(n2258)
         );
  NOR2_X1 U1821 ( .A1(n2248), .A2(n2247), .ZN(n2250) );
  OAI22_X1 U1822 ( .A1(n2246), .A2(n2245), .B1(n2244), .B2(n2243), .ZN(n2247)
         );
  OAI22_X1 U1823 ( .A1(n2242), .A2(n2241), .B1(n2240), .B2(n2239), .ZN(n2248)
         );
  INV_X1 U1824 ( .A(n2210), .ZN(n2242) );
  NOR2_X1 U1825 ( .A1(n2215), .A2(n2214), .ZN(n2252) );
  OAI211_X1 U1826 ( .C1(n2245), .C2(n2213), .A(n2212), .B(n2211), .ZN(n2214)
         );
  INV_X1 U1827 ( .A(n2059), .ZN(n2213) );
  OAI22_X1 U1828 ( .A1(n2244), .A2(n2208), .B1(n2239), .B2(n2207), .ZN(n2215)
         );
  AOI21_X1 U1829 ( .B1(n2238), .B2(n2237), .A(n2274), .ZN(n2272) );
  NAND2_X1 U1830 ( .A1(n2243), .A2(n2236), .ZN(n2237) );
  NAND2_X1 U1831 ( .A1(n2235), .A2(n2234), .ZN(n2238) );
  OAI22_X1 U1832 ( .A1(n2300), .A2(n1368), .B1(\COMP_REGN_ALUOUT/ffi_27/n4 ), 
        .B2(n1181), .ZN(\COMP_REGN_ALUOUT/ffi_27/n5 ) );
  INV_X1 U1833 ( .A(ALUOUT[27]), .ZN(n2300) );
  OAI21_X1 U1834 ( .B1(n2167), .B2(n2276), .A(n2166), .ZN(ALUOUT[27]) );
  AOI211_X1 U1835 ( .C1(n2165), .C2(n2164), .A(n2163), .B(n2162), .ZN(n2166)
         );
  NOR2_X1 U1836 ( .A1(n2161), .A2(n2268), .ZN(n2162) );
  NOR3_X1 U1837 ( .A1(n2160), .A2(n2159), .A3(n2158), .ZN(n2161) );
  OAI22_X1 U1838 ( .A1(n2263), .A2(n2217), .B1(n2265), .B2(n2255), .ZN(n2158)
         );
  NOR2_X1 U1839 ( .A1(n2107), .A2(n2106), .ZN(n2265) );
  OAI211_X1 U1840 ( .C1(n2245), .C2(n2105), .A(n2104), .B(n2211), .ZN(n2106)
         );
  NAND2_X1 U1841 ( .A1(n2210), .A2(n2103), .ZN(n2104) );
  OAI22_X1 U1842 ( .A1(n2244), .A2(n2102), .B1(n2239), .B2(n2101), .ZN(n2107)
         );
  INV_X1 U1843 ( .A(n2118), .ZN(n2102) );
  NOR2_X1 U1844 ( .A1(n2086), .A2(n2085), .ZN(n2263) );
  OAI22_X1 U1845 ( .A1(n2241), .A2(n1363), .B1(n2245), .B2(n2240), .ZN(n2085)
         );
  OAI211_X1 U1846 ( .C1(n2084), .C2(n2243), .A(n2083), .B(n2082), .ZN(n2086)
         );
  NAND2_X1 U1847 ( .A1(n2210), .A2(n2081), .ZN(n2082) );
  OAI22_X1 U1848 ( .A1(n2157), .A2(n1240), .B1(n2202), .B2(n2227), .ZN(n2159)
         );
  NOR2_X1 U1849 ( .A1(n2042), .A2(n2041), .ZN(n2202) );
  OAI22_X1 U1850 ( .A1(n2040), .A2(n1363), .B1(n2245), .B2(n2192), .ZN(n2041)
         );
  OAI211_X1 U1851 ( .C1(n2084), .C2(n2196), .A(n2083), .B(n2039), .ZN(n2042)
         );
  NAND2_X1 U1852 ( .A1(n2210), .A2(n2038), .ZN(n2039) );
  INV_X1 U1853 ( .A(n2221), .ZN(n2157) );
  NAND4_X1 U1854 ( .A1(n2066), .A2(n2065), .A3(n2064), .A4(n2063), .ZN(n2221)
         );
  NAND2_X1 U1855 ( .A1(n2062), .A2(n2228), .ZN(n2063) );
  INV_X1 U1856 ( .A(n2084), .ZN(n2062) );
  NAND2_X1 U1857 ( .A1(n2180), .A2(n2061), .ZN(n2064) );
  INV_X1 U1858 ( .A(n2245), .ZN(n2180) );
  AND2_X1 U1859 ( .A1(n2083), .A2(n2060), .ZN(n2066) );
  NAND2_X1 U1860 ( .A1(n2210), .A2(n2059), .ZN(n2060) );
  OAI211_X1 U1861 ( .C1(n2261), .C2(n2251), .A(n2156), .B(n2155), .ZN(n2160)
         );
  AOI22_X1 U1862 ( .A1(n1360), .A2(n2176), .B1(n2154), .B2(n2222), .ZN(n2155)
         );
  OAI22_X1 U1863 ( .A1(n2006), .A2(n1363), .B1(n2245), .B2(n1147), .ZN(n2007)
         );
  OAI211_X1 U1864 ( .C1(n2084), .C2(n2149), .A(n2083), .B(n2005), .ZN(n2008)
         );
  NAND2_X1 U1865 ( .A1(n2210), .A2(n2004), .ZN(n2005) );
  OAI22_X1 U1866 ( .A1(n2181), .A2(n1363), .B1(n2245), .B2(n2182), .ZN(n2024)
         );
  OAI211_X1 U1867 ( .C1(n2084), .C2(n2023), .A(n2083), .B(n2022), .ZN(n2025)
         );
  NAND2_X1 U1868 ( .A1(n2210), .A2(n2179), .ZN(n2022) );
  NAND2_X1 U1869 ( .A1(n1948), .A2(n1142), .ZN(n2084) );
  AOI22_X1 U1870 ( .A1(n1355), .A2(n2259), .B1(n2225), .B2(n1358), .ZN(n2156)
         );
  INV_X1 U1871 ( .A(n2254), .ZN(n2225) );
  INV_X1 U1872 ( .A(n1971), .ZN(n2124) );
  INV_X1 U1873 ( .A(n2120), .ZN(n2122) );
  INV_X1 U1874 ( .A(n2216), .ZN(n2259) );
  NOR2_X1 U1875 ( .A1(n2153), .A2(n2152), .ZN(n2216) );
  OAI211_X1 U1876 ( .C1(n2245), .C2(n1325), .A(n2151), .B(n2211), .ZN(n2152)
         );
  NAND2_X1 U1877 ( .A1(n2210), .A2(n2150), .ZN(n2151) );
  OAI22_X1 U1878 ( .A1(n2244), .A2(n2149), .B1(n2239), .B2(n2148), .ZN(n2153)
         );
  INV_X1 U1879 ( .A(n1989), .ZN(n2134) );
  NAND2_X1 U1880 ( .A1(n1954), .A2(n1953), .ZN(n2245) );
  AOI21_X1 U1881 ( .B1(n2147), .B2(n2146), .A(n2165), .ZN(n2163) );
  NAND2_X1 U1882 ( .A1(n2149), .A2(n2232), .ZN(n2146) );
  NAND2_X1 U1883 ( .A1(n2145), .A2(n2233), .ZN(n2147) );
  AND2_X1 U1884 ( .A1(n2305), .A2(ALU_OUT_REGN[0]), .ZN(n1272) );
  AOI21_X1 U1885 ( .B1(n1764), .B2(n2115), .A(n1763), .ZN(n1765) );
  INV_X1 U1886 ( .A(n1758), .ZN(n1764) );
  AOI211_X1 U1887 ( .C1(n2199), .C2(n1804), .A(n1757), .B(n1756), .ZN(n1766)
         );
  OAI211_X1 U1888 ( .C1(n2255), .C2(n1819), .A(n1754), .B(n1753), .ZN(n1757)
         );
  NAND2_X1 U1889 ( .A1(n1837), .A2(n1355), .ZN(n1753) );
  NAND2_X1 U1890 ( .A1(n1457), .A2(n1465), .ZN(n2249) );
  OAI211_X1 U1891 ( .C1(n2101), .C2(n2244), .A(n1496), .B(n1492), .ZN(n1837)
         );
  NAND2_X1 U1892 ( .A1(n1494), .A2(n1951), .ZN(n1492) );
  NAND2_X1 U1893 ( .A1(n1142), .A2(n1375), .ZN(n1441) );
  NAND2_X1 U1894 ( .A1(n1950), .A2(n1264), .ZN(n1496) );
  NOR2_X1 U1895 ( .A1(n1352), .A2(n1142), .ZN(n1264) );
  AND2_X1 U1896 ( .A1(n1376), .A2(ALU_OPCODE[1]), .ZN(n1429) );
  AOI21_X1 U1897 ( .B1(n1358), .B2(n1823), .A(n1752), .ZN(n1754) );
  OAI22_X1 U1898 ( .A1(n2262), .A2(n2101), .B1(n2217), .B2(n1810), .ZN(n1752)
         );
  NAND2_X1 U1899 ( .A1(n1251), .A2(n1375), .ZN(n1810) );
  INV_X1 U1900 ( .A(n1760), .ZN(n2101) );
  NAND2_X1 U1901 ( .A1(n1457), .A2(n1456), .ZN(n2262) );
  INV_X1 U1902 ( .A(n1464), .ZN(n1457) );
  AND2_X1 U1903 ( .A1(n2061), .A2(n1376), .ZN(n1823) );
  NAND2_X1 U1904 ( .A1(n1782), .A2(n1465), .ZN(n1455) );
  NAND2_X1 U1905 ( .A1(n1436), .A2(n1435), .ZN(n2255) );
  INV_X1 U1906 ( .A(n1472), .ZN(n1436) );
  NAND2_X1 U1907 ( .A1(n1464), .A2(n1759), .ZN(n1472) );
  AND2_X1 U1908 ( .A1(n1931), .A2(n1376), .ZN(n1804) );
  NAND2_X1 U1909 ( .A1(n1782), .A2(n1796), .ZN(n1463) );
  INV_X1 U1910 ( .A(n1445), .ZN(n1796) );
  INV_X1 U1911 ( .A(n1462), .ZN(n1782) );
  NAND2_X1 U1912 ( .A1(n1462), .A2(n1445), .ZN(n1464) );
  INV_X1 U1913 ( .A(n1771), .ZN(n1337) );
  OAI21_X1 U1914 ( .B1(ALU_OPCODE[2]), .B2(ALU_OPCODE[1]), .A(n1770), .ZN(
        n1771) );
  INV_X1 U1915 ( .A(n1751), .ZN(n1770) );
  AND2_X1 U1916 ( .A1(n1336), .A2(n2167), .ZN(n1273) );
  XNOR2_X1 U1917 ( .A(n1725), .B(n1724), .ZN(n2167) );
  XNOR2_X1 U1918 ( .A(n1723), .B(n2145), .ZN(n1724) );
  INV_X1 U1919 ( .A(n2149), .ZN(n2145) );
  NAND2_X1 U1920 ( .A1(n1722), .A2(n1721), .ZN(n1725) );
  XNOR2_X1 U1921 ( .A(n1304), .B(n1720), .ZN(n2206) );
  AND2_X1 U1922 ( .A1(n2231), .A2(n2191), .ZN(n1336) );
  XNOR2_X1 U1923 ( .A(n1231), .B(n1748), .ZN(n2231) );
  OAI21_X1 U1924 ( .B1(n1637), .B2(n1636), .A(n1722), .ZN(n2144) );
  OAI21_X1 U1925 ( .B1(n1704), .B2(n1296), .A(n1294), .ZN(n1722) );
  NOR2_X1 U1926 ( .A1(n1600), .A2(n1295), .ZN(n1294) );
  NOR2_X1 U1927 ( .A1(n1639), .A2(n1296), .ZN(n1295) );
  INV_X1 U1928 ( .A(n1635), .ZN(n1296) );
  INV_X1 U1929 ( .A(n1634), .ZN(n1635) );
  XNOR2_X1 U1930 ( .A(n1747), .B(n1746), .ZN(n2055) );
  AND2_X1 U1931 ( .A1(n1316), .A2(n1744), .ZN(n1292) );
  XNOR2_X1 U1932 ( .A(n1632), .B(n1227), .ZN(n2077) );
  INV_X1 U1933 ( .A(n1316), .ZN(n1315) );
  XNOR2_X1 U1934 ( .A(n1674), .B(n2118), .ZN(n1675) );
  INV_X1 U1935 ( .A(n1669), .ZN(n1671) );
  XNOR2_X1 U1936 ( .A(n1531), .B(n1530), .ZN(n1668) );
  AND2_X1 U1937 ( .A1(n1529), .A2(n1548), .ZN(n1530) );
  AOI21_X1 U1938 ( .B1(n1528), .B2(n1527), .A(n1526), .ZN(n1531) );
  XNOR2_X1 U1939 ( .A(n1528), .B(n1513), .ZN(n1667) );
  AOI211_X1 U1940 ( .C1(n1665), .C2(n1664), .A(n1663), .B(n1802), .ZN(n1666)
         );
  XNOR2_X1 U1941 ( .A(n1657), .B(n1656), .ZN(n1787) );
  XNOR2_X1 U1942 ( .A(n1759), .B(n1760), .ZN(n1758) );
  NAND2_X1 U1943 ( .A1(n1141), .A2(n1652), .ZN(n1653) );
  NAND2_X1 U1944 ( .A1(n1512), .A2(n1488), .ZN(n1664) );
  NAND2_X1 U1945 ( .A1(n1665), .A2(n1650), .ZN(n1651) );
  OR2_X1 U1946 ( .A1(n1512), .A2(n1488), .ZN(n1665) );
  OAI21_X1 U1947 ( .B1(n1144), .B2(n1416), .A(n1331), .ZN(n1333) );
  AOI21_X1 U1948 ( .B1(n1334), .B2(n1332), .A(n1127), .ZN(n1331) );
  INV_X1 U1949 ( .A(n1549), .ZN(n1332) );
  NAND2_X1 U1950 ( .A1(n1903), .A2(n1902), .ZN(n1673) );
  OR2_X1 U1951 ( .A1(n1646), .A2(n1133), .ZN(n1902) );
  NAND2_X1 U1952 ( .A1(n1646), .A2(n1133), .ZN(n1903) );
  OAI21_X1 U1953 ( .B1(n1321), .B2(n1643), .A(n1644), .ZN(n1320) );
  INV_X1 U1954 ( .A(n1321), .ZN(n1319) );
  NAND2_X1 U1955 ( .A1(n1642), .A2(n1645), .ZN(n1321) );
  INV_X1 U1956 ( .A(n1633), .ZN(n1639) );
  NOR2_X1 U1957 ( .A1(n1692), .A2(n1693), .ZN(n1703) );
  NAND4_X1 U1958 ( .A1(n1943), .A2(n1862), .A3(n1924), .A4(n1891), .ZN(n1692)
         );
  XNOR2_X1 U1959 ( .A(n1691), .B(n1690), .ZN(n1891) );
  XNOR2_X1 U1960 ( .A(n1689), .B(n2179), .ZN(n1690) );
  XNOR2_X1 U1961 ( .A(n1688), .B(n1687), .ZN(n1924) );
  AOI21_X1 U1962 ( .B1(n1686), .B2(n1149), .A(n1171), .ZN(n1688) );
  XNOR2_X1 U1963 ( .A(n1681), .B(n2081), .ZN(n1682) );
  NAND2_X1 U1964 ( .A1(n1335), .A2(n1246), .ZN(n1679) );
  XNOR2_X1 U1965 ( .A(n1425), .B(n1424), .ZN(n1693) );
  NAND2_X1 U1966 ( .A1(n1669), .A2(n1422), .ZN(n1672) );
  INV_X1 U1967 ( .A(n1152), .ZN(n1422) );
  INV_X1 U1968 ( .A(n1556), .ZN(n1513) );
  INV_X1 U1969 ( .A(n1326), .ZN(n1328) );
  INV_X1 U1970 ( .A(n1729), .ZN(n1730) );
  NOR2_X1 U1971 ( .A1(n1746), .A2(n1629), .ZN(n1727) );
  INV_X1 U1972 ( .A(n1628), .ZN(n1629) );
  INV_X1 U1973 ( .A(n1627), .ZN(n1329) );
  NAND2_X1 U1974 ( .A1(n1734), .A2(n1733), .ZN(n1735) );
  INV_X1 U1975 ( .A(n1732), .ZN(n1330) );
  INV_X1 U1976 ( .A(n1726), .ZN(n1732) );
  NAND2_X1 U1977 ( .A1(n1582), .A2(n1736), .ZN(n1327) );
  INV_X1 U1978 ( .A(n1280), .ZN(n1279) );
  OAI21_X1 U1979 ( .B1(n1344), .B2(n1241), .A(n1699), .ZN(n1280) );
  INV_X1 U1980 ( .A(n1698), .ZN(n1699) );
  OR2_X1 U1981 ( .A1(n1740), .A2(n1696), .ZN(n1241) );
  INV_X1 U1982 ( .A(n1695), .ZN(n1696) );
  NAND2_X1 U1983 ( .A1(n1291), .A2(n1626), .ZN(n1745) );
  NAND2_X1 U1984 ( .A1(n1229), .A2(n1316), .ZN(n1291) );
  NOR2_X1 U1985 ( .A1(n1627), .A2(n1182), .ZN(n1316) );
  NAND2_X1 U1986 ( .A1(n1624), .A2(n1700), .ZN(n1627) );
  INV_X1 U1987 ( .A(n1345), .ZN(n1344) );
  OAI21_X1 U1988 ( .B1(n1566), .B2(n1346), .A(n1622), .ZN(n1345) );
  OAI21_X1 U1989 ( .B1(n1714), .B2(n1183), .A(n1713), .ZN(n1715) );
  OAI21_X1 U1990 ( .B1(n1712), .B2(n1711), .A(n1710), .ZN(n1713) );
  INV_X1 U1991 ( .A(n1709), .ZN(n1711) );
  AOI21_X1 U1992 ( .B1(n1708), .B2(n1245), .A(n1707), .ZN(n1714) );
  INV_X1 U1993 ( .A(n1139), .ZN(n1706) );
  AND2_X1 U1994 ( .A1(n1577), .A2(n1349), .ZN(n1299) );
  AND2_X1 U1995 ( .A1(n1256), .A2(n1255), .ZN(n1254) );
  AND2_X1 U1996 ( .A1(n1734), .A2(n1349), .ZN(n1257) );
  INV_X1 U1997 ( .A(ALU_OPCODE[2]), .ZN(n1768) );
  NAND2_X1 U1998 ( .A1(n1750), .A2(ALU_OPCODE[5]), .ZN(n1751) );
  INV_X1 U1999 ( .A(ALU_OPCODE[4]), .ZN(n1750) );
  INV_X1 U2000 ( .A(n1284), .ZN(n1281) );
  AND2_X1 U2001 ( .A1(n1619), .A2(n1288), .ZN(n1287) );
  NAND2_X1 U2002 ( .A1(n1302), .A2(n1748), .ZN(n1288) );
  AOI21_X1 U2003 ( .B1(n1616), .B2(n1716), .A(n1615), .ZN(n1619) );
  OAI21_X1 U2004 ( .B1(n1617), .B2(n1614), .A(n1613), .ZN(n1615) );
  NAND2_X1 U2005 ( .A1(n1612), .A2(n1716), .ZN(n1613) );
  INV_X1 U2006 ( .A(n1618), .ZN(n1614) );
  NOR2_X1 U2007 ( .A1(n1303), .A2(n1748), .ZN(n1289) );
  INV_X1 U2008 ( .A(n2228), .ZN(n2208) );
  NAND2_X1 U2009 ( .A1(n1610), .A2(n2228), .ZN(n1611) );
  NOR2_X1 U2010 ( .A1(n1546), .A2(n1617), .ZN(n1612) );
  INV_X1 U2011 ( .A(n1717), .ZN(n1546) );
  NOR3_X1 U2012 ( .A1(n1618), .A2(n1717), .A3(n2274), .ZN(n1616) );
  INV_X1 U2013 ( .A(n1617), .ZN(n2274) );
  NOR2_X1 U2014 ( .A1(n1717), .A2(n2243), .ZN(n1618) );
  INV_X1 U2015 ( .A(NPC1[31]), .ZN(n1427) );
  INV_X1 U2016 ( .A(A[31]), .ZN(n1428) );
  XNOR2_X1 U2017 ( .A(n1617), .B(n1374), .ZN(n1717) );
  NOR2_X1 U2018 ( .A1(n1324), .A2(n1712), .ZN(n1323) );
  INV_X1 U2019 ( .A(n1339), .ZN(n1324) );
  NAND2_X1 U2020 ( .A1(n1606), .A2(n2023), .ZN(n1709) );
  INV_X1 U2021 ( .A(n2178), .ZN(n2023) );
  INV_X1 U2022 ( .A(n1605), .ZN(n1606) );
  INV_X1 U2023 ( .A(n1707), .ZN(n1342) );
  AND2_X1 U2024 ( .A1(n1723), .A2(n2149), .ZN(n1707) );
  XNOR2_X1 U2025 ( .A(n1601), .B(n2120), .ZN(n1633) );
  INV_X1 U2026 ( .A(n1710), .ZN(n1608) );
  INV_X1 U2027 ( .A(n1718), .ZN(n1609) );
  NAND2_X1 U2028 ( .A1(n1605), .A2(n2178), .ZN(n1718) );
  INV_X1 U2029 ( .A(n1712), .ZN(n1720) );
  INV_X1 U2030 ( .A(n2204), .ZN(n2196) );
  NAND2_X1 U2031 ( .A1(n1607), .A2(n2204), .ZN(n1710) );
  AND2_X1 U2032 ( .A1(n1139), .A2(n1348), .ZN(n1237) );
  OAI21_X1 U2033 ( .B1(n1723), .B2(n2149), .A(n1721), .ZN(n1604) );
  INV_X1 U2034 ( .A(NPC1[27]), .ZN(n1602) );
  INV_X1 U2035 ( .A(A[27]), .ZN(n1603) );
  XNOR2_X1 U2036 ( .A(n2165), .B(n1372), .ZN(n1723) );
  AND2_X1 U2037 ( .A1(n1601), .A2(n2120), .ZN(n1634) );
  NAND2_X1 U2038 ( .A1(n1721), .A2(n1599), .ZN(n1600) );
  NAND2_X1 U2039 ( .A1(n1598), .A2(n2132), .ZN(n1599) );
  INV_X1 U2040 ( .A(n2128), .ZN(n2132) );
  INV_X1 U2041 ( .A(n1597), .ZN(n1598) );
  NAND2_X1 U2042 ( .A1(n1597), .A2(n2128), .ZN(n1721) );
  NAND2_X1 U2043 ( .A1(n1351), .A2(n1258), .ZN(n1676) );
  NAND2_X1 U2044 ( .A1(n1593), .A2(n1592), .ZN(n1733) );
  INV_X1 U2045 ( .A(n2241), .ZN(n1592) );
  INV_X1 U2046 ( .A(n1591), .ZN(n1593) );
  AND2_X1 U2047 ( .A1(n1729), .A2(n1590), .ZN(n1726) );
  AOI21_X1 U2048 ( .B1(n1631), .B2(n1587), .A(n1586), .ZN(n1729) );
  NOR2_X1 U2049 ( .A1(n1228), .A2(n1914), .ZN(n1586) );
  NAND2_X1 U2050 ( .A1(n1584), .A2(n2081), .ZN(n1622) );
  INV_X1 U2051 ( .A(n2246), .ZN(n2081) );
  INV_X1 U2052 ( .A(n1681), .ZN(n1584) );
  NOR2_X1 U2053 ( .A1(n1174), .A2(n1746), .ZN(n1596) );
  INV_X1 U2054 ( .A(n1589), .ZN(n1746) );
  INV_X1 U2055 ( .A(n1702), .ZN(n1700) );
  NAND2_X1 U2056 ( .A1(n1580), .A2(n2123), .ZN(n1581) );
  INV_X1 U2057 ( .A(n2150), .ZN(n2006) );
  NAND2_X1 U2058 ( .A1(n1734), .A2(n1621), .ZN(n1576) );
  NAND2_X1 U2059 ( .A1(n1681), .A2(n2246), .ZN(n1621) );
  INV_X1 U2060 ( .A(NPC1[15]), .ZN(n1459) );
  INV_X1 U2061 ( .A(A[15]), .ZN(n1460) );
  XNOR2_X1 U2062 ( .A(n1938), .B(n1373), .ZN(n1681) );
  NAND2_X1 U2063 ( .A1(n1591), .A2(n2241), .ZN(n1734) );
  INV_X1 U2064 ( .A(NPC1[23]), .ZN(n1574) );
  INV_X1 U2065 ( .A(A[23]), .ZN(n1575) );
  XNOR2_X1 U2066 ( .A(n2078), .B(n1373), .ZN(n1591) );
  NAND2_X1 U2067 ( .A1(n1571), .A2(n1990), .ZN(n1572) );
  INV_X1 U2068 ( .A(n2133), .ZN(n1990) );
  NAND2_X1 U2069 ( .A1(n1569), .A2(n1955), .ZN(n1695) );
  INV_X1 U2070 ( .A(n2103), .ZN(n1955) );
  INV_X1 U2071 ( .A(n2194), .ZN(n2040) );
  NAND2_X1 U2072 ( .A1(n1175), .A2(n2181), .ZN(n1628) );
  BUF_X1 U2073 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .Z(n1373) );
  NAND2_X1 U2074 ( .A1(n1565), .A2(n2059), .ZN(n1566) );
  XNOR2_X1 U2075 ( .A(n1565), .B(n2059), .ZN(n1687) );
  INV_X1 U2076 ( .A(n1561), .ZN(n1562) );
  INV_X1 U2077 ( .A(n2061), .ZN(n2207) );
  AOI21_X1 U2078 ( .B1(n1313), .B2(n1486), .A(n1410), .ZN(n1511) );
  INV_X1 U2079 ( .A(n1897), .ZN(n2192) );
  AND2_X1 U2080 ( .A1(n1252), .A2(n1251), .ZN(n1486) );
  NAND2_X1 U2081 ( .A1(n1385), .A2(n1947), .ZN(n1252) );
  INV_X1 U2082 ( .A(n2131), .ZN(n1788) );
  INV_X1 U2083 ( .A(n1402), .ZN(n1403) );
  INV_X1 U2084 ( .A(n1401), .ZN(n1404) );
  OAI21_X1 U2085 ( .B1(n1402), .B2(n1401), .A(n1400), .ZN(n1406) );
  OAI21_X1 U2086 ( .B1(S1_A_NPC), .B2(A[0]), .A(n1399), .ZN(n1400) );
  NAND2_X1 U2087 ( .A1(S1_A_NPC), .A2(n1398), .ZN(n1399) );
  INV_X1 U2088 ( .A(NPC1[0]), .ZN(n1398) );
  INV_X1 U2089 ( .A(IMM[0]), .ZN(n1397) );
  INV_X1 U2090 ( .A(IMM[1]), .ZN(n1433) );
  INV_X1 U2091 ( .A(NPC1[2]), .ZN(n1390) );
  INV_X1 U2092 ( .A(A[2]), .ZN(n1391) );
  INV_X1 U2093 ( .A(IMM[2]), .ZN(n1434) );
  XNOR2_X1 U2094 ( .A(n1409), .B(n1897), .ZN(n1313) );
  XNOR2_X1 U2095 ( .A(n1827), .B(n1372), .ZN(n1409) );
  INV_X1 U2096 ( .A(NPC1[4]), .ZN(n1386) );
  INV_X1 U2097 ( .A(A[4]), .ZN(n1387) );
  INV_X1 U2098 ( .A(IMM[4]), .ZN(n1384) );
  NOR2_X1 U2099 ( .A1(n1555), .A2(n1554), .ZN(n1685) );
  NOR2_X1 U2100 ( .A1(n1561), .A2(n1236), .ZN(n1554) );
  INV_X1 U2101 ( .A(n2038), .ZN(n2193) );
  INV_X1 U2102 ( .A(n1885), .ZN(n2179) );
  INV_X1 U2103 ( .A(n1689), .ZN(n1552) );
  INV_X1 U2104 ( .A(NPC1[12]), .ZN(n1442) );
  INV_X1 U2105 ( .A(A[12]), .ZN(n1443) );
  XNOR2_X1 U2106 ( .A(n1886), .B(n1375), .ZN(n1689) );
  NAND2_X1 U2107 ( .A1(n1680), .A2(n1421), .ZN(n1550) );
  NAND2_X1 U2108 ( .A1(n1420), .A2(n1971), .ZN(n1421) );
  INV_X1 U2109 ( .A(n1158), .ZN(n1419) );
  NAND2_X1 U2110 ( .A1(n1277), .A2(n1989), .ZN(n1558) );
  INV_X1 U2111 ( .A(n2240), .ZN(n1931) );
  INV_X1 U2112 ( .A(NPC1[7]), .ZN(n1413) );
  INV_X1 U2113 ( .A(A[7]), .ZN(n1414) );
  BUF_X1 U2114 ( .A(\COMP_ALU/ADD_SUB/carries_s[0] ), .Z(n1374) );
  INV_X1 U2115 ( .A(n1951), .ZN(n2105) );
  OR2_X1 U2116 ( .A1(n1164), .A2(n1325), .ZN(n1236) );
  INV_X1 U2117 ( .A(n1588), .ZN(n1743) );
  INV_X1 U2118 ( .A(n2211), .ZN(n1950) );
  AND2_X1 U2119 ( .A1(n2211), .A2(n1270), .ZN(n1239) );
  NAND2_X1 U2120 ( .A1(n1689), .A2(n1885), .ZN(n1644) );
  AND2_X1 U2121 ( .A1(n1145), .A2(n1309), .ZN(n1242) );
  AND3_X1 U2122 ( .A1(n1449), .A2(n1448), .A3(n1447), .ZN(n1243) );
  INV_X1 U2123 ( .A(n2031), .ZN(n2181) );
  INV_X1 U2124 ( .A(n1611), .ZN(n1716) );
  MUX2_X1 U2125 ( .A(n1387), .B(n1386), .S(S1_A_NPC), .Z(n2182) );
  INV_X1 U2126 ( .A(n2182), .ZN(n1251) );
  AND2_X1 U2127 ( .A1(n1334), .A2(n1127), .ZN(n1246) );
  INV_X1 U2128 ( .A(n1144), .ZN(n1334) );
  OR2_X1 U2129 ( .A1(n1706), .A2(n1183), .ZN(n1247) );
  INV_X1 U2130 ( .A(n1600), .ZN(n1637) );
  AND2_X1 U2131 ( .A1(n2206), .A2(n1337), .ZN(n1248) );
  NAND2_X1 U2132 ( .A1(n1552), .A2(n2179), .ZN(n1645) );
  AND2_X1 U2133 ( .A1(n1626), .A2(n1330), .ZN(n1249) );
  INV_X1 U2134 ( .A(n1621), .ZN(n1346) );
  INV_X1 U2135 ( .A(n1738), .ZN(n1744) );
  INV_X1 U2136 ( .A(n1348), .ZN(n1301) );
  AND2_X1 U2137 ( .A1(n1281), .A2(n1237), .ZN(n1250) );
  NAND3_X1 U2138 ( .A1(n1385), .A2(n1947), .A3(n2182), .ZN(n1487) );
  INV_X1 U2139 ( .A(n1951), .ZN(n1253) );
  XNOR2_X1 U2140 ( .A(n1834), .B(n1372), .ZN(n1418) );
  AOI21_X1 U2141 ( .B1(n1595), .B2(n1257), .A(n1301), .ZN(n1256) );
  NAND2_X1 U2142 ( .A1(n1350), .A2(n1257), .ZN(n1255) );
  NOR2_X1 U2143 ( .A1(n1259), .A2(n2116), .ZN(n1307) );
  NAND4_X1 U2144 ( .A1(n1967), .A2(n1673), .A3(n1262), .A4(n1876), .ZN(n1259)
         );
  NAND2_X1 U2145 ( .A1(n1261), .A2(n1672), .ZN(n1876) );
  NAND2_X1 U2146 ( .A1(n1260), .A2(n1741), .ZN(n1967) );
  NAND2_X1 U2147 ( .A1(n1697), .A2(n1623), .ZN(n1741) );
  NAND2_X1 U2148 ( .A1(n1648), .A2(n1647), .ZN(n1260) );
  NAND2_X1 U2149 ( .A1(n1671), .A2(n1152), .ZN(n1261) );
  NOR2_X1 U2150 ( .A1(n1263), .A2(n1668), .ZN(n1262) );
  NAND4_X1 U2151 ( .A1(n1847), .A2(n1833), .A3(n1666), .A4(n1667), .ZN(n1263)
         );
  NAND3_X1 U2152 ( .A1(n1336), .A2(n2206), .A3(n2167), .ZN(n1268) );
  NAND4_X1 U2153 ( .A1(n1265), .A2(n1273), .A3(n1267), .A4(n1244), .ZN(n1266)
         );
  AND2_X1 U2154 ( .A1(n1275), .A2(n1224), .ZN(n1265) );
  AND2_X1 U2155 ( .A1(n1248), .A2(n1274), .ZN(n1267) );
  NAND2_X1 U2156 ( .A1(n2210), .A2(n2031), .ZN(n1270) );
  NOR2_X1 U2157 ( .A1(n1953), .A2(n1142), .ZN(n1271) );
  AOI21_X1 U2158 ( .B1(ALUOUT[0]), .B2(n2306), .A(n1272), .ZN(n2277) );
  NOR2_X1 U2159 ( .A1(n1749), .A2(n1306), .ZN(n1275) );
  NAND2_X1 U2160 ( .A1(n1558), .A2(n1670), .ZN(n1560) );
  XNOR2_X1 U2161 ( .A(n1277), .B(n1989), .ZN(n1670) );
  XNOR2_X1 U2162 ( .A(n1863), .B(n1353), .ZN(n1277) );
  OAI22_X1 U2163 ( .A1(n1582), .A2(n1736), .B1(n2006), .B2(n1278), .ZN(n1312)
         );
  INV_X1 U2164 ( .A(n1737), .ZN(n1582) );
  XNOR2_X1 U2165 ( .A(n1278), .B(n2150), .ZN(n1737) );
  XNOR2_X1 U2166 ( .A(n2014), .B(n1373), .ZN(n1278) );
  OAI21_X1 U2167 ( .B1(n1241), .B2(n1343), .A(n1279), .ZN(n1701) );
  OAI21_X1 U2168 ( .B1(n1323), .B2(n1284), .A(n1287), .ZN(n1283) );
  NAND2_X1 U2169 ( .A1(n1705), .A2(n1302), .ZN(n1284) );
  NOR2_X1 U2170 ( .A1(n1340), .A2(n1183), .ZN(n1285) );
  OAI21_X1 U2171 ( .B1(n1138), .B2(n1183), .A(n1289), .ZN(n1286) );
  AOI21_X1 U2172 ( .B1(n1229), .B2(n1292), .A(n1290), .ZN(n1747) );
  OAI21_X1 U2173 ( .B1(n1626), .B2(n1220), .A(n1588), .ZN(n1290) );
  NAND2_X1 U2174 ( .A1(n1638), .A2(n1635), .ZN(n1636) );
  XNOR2_X1 U2175 ( .A(n1518), .B(n1377), .ZN(n1412) );
  OAI21_X1 U2176 ( .B1(n1380), .B2(n1298), .A(n1297), .ZN(n1518) );
  NAND2_X1 U2177 ( .A1(n1160), .A2(B[6]), .ZN(n1297) );
  INV_X1 U2178 ( .A(IMM[6]), .ZN(n1298) );
  NAND2_X1 U2179 ( .A1(n1683), .A2(n1577), .ZN(n1351) );
  NAND2_X1 U2180 ( .A1(n1347), .A2(n1566), .ZN(n1683) );
  NAND2_X1 U2181 ( .A1(n1226), .A2(n1299), .ZN(n1300) );
  NOR2_X1 U2182 ( .A1(n1176), .A2(ALU_OPCODE[1]), .ZN(n1769) );
  NOR2_X1 U2183 ( .A1(n1616), .A2(n1612), .ZN(n1303) );
  NAND2_X1 U2184 ( .A1(n1719), .A2(n1718), .ZN(n1304) );
  OAI21_X1 U2185 ( .B1(n1231), .B2(n1748), .A(n1611), .ZN(n1305) );
  NAND4_X1 U2186 ( .A1(n1307), .A2(n2126), .A3(n1703), .A4(n2001), .ZN(n1306)
         );
  INV_X1 U2187 ( .A(n1349), .ZN(n1308) );
  INV_X1 U2188 ( .A(n1143), .ZN(n1309) );
  NAND3_X1 U2189 ( .A1(n1698), .A2(n1309), .A3(n1700), .ZN(n1310) );
  NAND2_X1 U2190 ( .A1(n1311), .A2(n1310), .ZN(n1625) );
  INV_X1 U2191 ( .A(n1312), .ZN(n1311) );
  XNOR2_X1 U2192 ( .A(n1651), .B(n1154), .ZN(n1833) );
  AOI21_X1 U2193 ( .B1(n1317), .B2(n1319), .A(n1320), .ZN(n1646) );
  INV_X1 U2194 ( .A(n1686), .ZN(n1317) );
  NAND2_X1 U2195 ( .A1(n1318), .A2(n1642), .ZN(n1691) );
  NAND2_X1 U2196 ( .A1(n1643), .A2(n1686), .ZN(n1318) );
  INV_X1 U2197 ( .A(n1715), .ZN(n1322) );
  INV_X1 U2198 ( .A(n2004), .ZN(n1325) );
  XNOR2_X1 U2199 ( .A(n1478), .B(\COMP_ALU/ADD_SUB/carries_s[0] ), .ZN(n1423)
         );
  NAND2_X1 U2200 ( .A1(n1416), .A2(n1157), .ZN(n1335) );
  NAND2_X1 U2201 ( .A1(n1679), .A2(n1333), .ZN(n1847) );
  NAND3_X1 U2202 ( .A1(n1564), .A2(n1621), .A3(n1563), .ZN(n1343) );
  NAND2_X1 U2203 ( .A1(n1564), .A2(n1563), .ZN(n1347) );
  NAND2_X1 U2204 ( .A1(n1674), .A2(n2118), .ZN(n1348) );
  INV_X1 U2205 ( .A(n2277), .ZN(n2) );
  NOR2_X1 U2206 ( .A1(n2192), .A2(n1169), .ZN(n1410) );
  INV_X1 U2207 ( .A(n1134), .ZN(n1526) );
  NAND2_X1 U2208 ( .A1(n1525), .A2(n1527), .ZN(n1556) );
  NAND2_X1 U2209 ( .A1(n1643), .A2(n1562), .ZN(n1684) );
  NAND2_X1 U2210 ( .A1(n1567), .A2(n2031), .ZN(n1588) );
  XNOR2_X1 U2211 ( .A(n1417), .B(n1971), .ZN(n1678) );
  XNOR2_X1 U2212 ( .A(n1848), .B(n1374), .ZN(n1417) );
  NAND2_X1 U2213 ( .A1(n1232), .A2(n1931), .ZN(n1529) );
  NOR2_X1 U2214 ( .A1(n1455), .A2(n1135), .ZN(n2220) );
  NAND2_X1 U2215 ( .A1(n1440), .A2(n1788), .ZN(n1659) );
  INV_X1 U2216 ( .A(n1647), .ZN(n1623) );
  NAND2_X1 U2217 ( .A1(n2210), .A2(n2209), .ZN(n2212) );
  NAND2_X1 U2218 ( .A1(n1364), .A2(n2209), .ZN(n2065) );
  INV_X1 U2219 ( .A(n2209), .ZN(n1914) );
  NAND2_X1 U2220 ( .A1(n1393), .A2(n2148), .ZN(n1661) );
  INV_X1 U2221 ( .A(n1658), .ZN(n1652) );
  NAND2_X1 U2222 ( .A1(n1742), .A2(n1581), .ZN(n1698) );
  INV_X1 U2223 ( .A(n1223), .ZN(n1580) );
  XNOR2_X1 U2224 ( .A(n1968), .B(n1376), .ZN(n1579) );
  AND2_X1 U2225 ( .A1(n1677), .A2(n1547), .ZN(n1649) );
  NAND2_X1 U2226 ( .A1(n1418), .A2(n2105), .ZN(n1547) );
  NAND2_X1 U2227 ( .A1(n1739), .A2(n1695), .ZN(n1647) );
  NAND2_X1 U2228 ( .A1(n1897), .A2(n1375), .ZN(n1819) );
  NAND2_X1 U2229 ( .A1(n1678), .A2(n1419), .ZN(n1680) );
  NOR2_X1 U2230 ( .A1(n1647), .A2(n1702), .ZN(n1573) );
  INV_X1 U2231 ( .A(n1454), .ZN(n1440) );
  XNOR2_X1 U2232 ( .A(n1389), .B(n1372), .ZN(n1454) );
  INV_X1 U2233 ( .A(n1194), .ZN(n1424) );
  XNOR2_X1 U2234 ( .A(n1423), .B(n2004), .ZN(n1559) );
  NAND2_X1 U2235 ( .A1(n1736), .A2(n1572), .ZN(n1702) );
  INV_X1 U2236 ( .A(n1694), .ZN(n1740) );
  AND2_X1 U2237 ( .A1(n1737), .A2(n1694), .ZN(n1624) );
  AOI21_X1 U2238 ( .B1(n1685), .B2(n1684), .A(n1687), .ZN(n1563) );
  NOR2_X1 U2239 ( .A1(n1551), .A2(n1550), .ZN(n1641) );
  OAI22_X1 U2240 ( .A1(n1561), .A2(n1645), .B1(n2193), .B2(n1155), .ZN(n1555)
         );
  NAND2_X1 U2241 ( .A1(n1136), .A2(n1137), .ZN(n1657) );
  INV_X1 U2242 ( .A(n1630), .ZN(n1587) );
  INV_X1 U2243 ( .A(n1625), .ZN(n1626) );
  NAND2_X1 U2244 ( .A1(n1662), .A2(n1658), .ZN(n1394) );
  NAND2_X1 U2245 ( .A1(n1412), .A2(n2061), .ZN(n1525) );
  XNOR2_X1 U2246 ( .A(n1904), .B(n1373), .ZN(n1553) );
  INV_X1 U2247 ( .A(n1570), .ZN(n1571) );
  NAND2_X1 U2248 ( .A1(n2133), .A2(n1570), .ZN(n1736) );
  XNOR2_X1 U2249 ( .A(n1745), .B(n1744), .ZN(n2037) );
  OAI211_X1 U2250 ( .C1(n1222), .C2(n2276), .A(n1966), .B(n1965), .ZN(
        ALUOUT[16]) );
  NAND2_X1 U2251 ( .A1(n1415), .A2(n2240), .ZN(n1548) );
  XNOR2_X1 U2252 ( .A(n1540), .B(n1374), .ZN(n1415) );
  INV_X1 U2253 ( .A(n1568), .ZN(n1569) );
  NAND2_X1 U2254 ( .A1(n2098), .A2(n1375), .ZN(n1947) );
  NAND2_X1 U2255 ( .A1(n1484), .A2(n1140), .ZN(n1512) );
  AND2_X1 U2256 ( .A1(S2_IMM_B), .A2(B[0]), .ZN(n1402) );
  OAI21_X1 U2257 ( .B1(n1170), .B2(n1549), .A(n1558), .ZN(n1551) );
  NAND2_X1 U2258 ( .A1(n1672), .A2(n1558), .ZN(n1425) );
  XNOR2_X1 U2259 ( .A(n1848), .B(n1378), .ZN(n1420) );
  NOR2_X1 U2260 ( .A1(n1759), .A2(n1354), .ZN(n1456) );
  NOR2_X1 U2261 ( .A1(n1755), .A2(n1353), .ZN(n1756) );
  OAI21_X1 U2262 ( .B1(n1779), .B2(n1354), .A(n1778), .ZN(n1780) );
  NAND2_X1 U2263 ( .A1(n1407), .A2(n1781), .ZN(n1655) );
  NAND2_X1 U2264 ( .A1(n2210), .A2(n1200), .ZN(n1438) );
  AOI222_X1 U2265 ( .A1(n1359), .A2(n1200), .B1(n1184), .B2(n1813), .C1(n1788), 
        .C2(n1361), .ZN(n1755) );
  AOI222_X1 U2266 ( .A1(n1359), .A2(n1788), .B1(n2222), .B2(n1200), .C1(n1362), 
        .C2(n1813), .ZN(n1779) );
  NOR2_X1 U2267 ( .A1(n1179), .A2(n1230), .ZN(n1731) );
  XNOR2_X1 U2268 ( .A(n2229), .B(n1377), .ZN(n1610) );
  XNOR2_X1 U2269 ( .A(n2117), .B(n1353), .ZN(n1674) );
  XNOR2_X1 U2270 ( .A(n2172), .B(n1377), .ZN(n1605) );
  XNOR2_X1 U2271 ( .A(n2119), .B(n1378), .ZN(n1601) );
  XNOR2_X1 U2272 ( .A(n2205), .B(n1354), .ZN(n1607) );
  XNOR2_X1 U2273 ( .A(n2127), .B(n1353), .ZN(n1597) );
  INV_X1 U2274 ( .A(n1728), .ZN(n1631) );
  XNOR2_X1 U2275 ( .A(n1919), .B(n1377), .ZN(n1565) );
  XNOR2_X1 U2276 ( .A(n1585), .B(n2209), .ZN(n1728) );
  XNOR2_X1 U2277 ( .A(n2032), .B(n1354), .ZN(n1567) );
  XNOR2_X1 U2278 ( .A(n1986), .B(n1354), .ZN(n1570) );
  XNOR2_X1 U2279 ( .A(n2072), .B(n1378), .ZN(n1585) );
  OR2_X1 U2280 ( .A1(n1781), .A2(n1407), .ZN(n1654) );
  XNOR2_X1 U2281 ( .A(n1396), .B(n1378), .ZN(n1407) );
  INV_X1 U2282 ( .A(n1200), .ZN(n2121) );
  AOI21_X1 U2283 ( .B1(n1720), .B2(n1609), .A(n1608), .ZN(n1705) );
  OAI21_X1 U2284 ( .B1(n1766), .B2(n2268), .A(n1765), .ZN(n1767) );
  NAND2_X1 U2285 ( .A1(n1655), .A2(n1656), .ZN(n1408) );
  NAND2_X1 U2286 ( .A1(n1487), .A2(n1650), .ZN(n1488) );
  INV_X1 U2287 ( .A(n1486), .ZN(n1650) );
  INV_X1 U2288 ( .A(n1697), .ZN(n1648) );
  NAND2_X1 U2289 ( .A1(n1953), .A2(n1354), .ZN(n1385) );
  NAND2_X1 U2290 ( .A1(n1408), .A2(n1654), .ZN(n1660) );
  XNOR2_X1 U2291 ( .A(n1676), .B(n1675), .ZN(n2116) );
  XNOR2_X1 U2292 ( .A(n1177), .B(n1653), .ZN(n1801) );
  OAI211_X1 U2293 ( .C1(n1594), .C2(n1622), .A(n1726), .B(n1733), .ZN(n1595)
         );
  NOR2_X1 U2294 ( .A1(n1594), .A2(n1576), .ZN(n1577) );
  NAND4_X1 U2295 ( .A1(n1583), .A2(n1624), .A3(n1589), .A4(n1573), .ZN(n1594)
         );
  NAND2_X1 U2296 ( .A1(n2100), .A2(n1235), .ZN(n2239) );
  NAND2_X1 U2297 ( .A1(n1640), .A2(n1233), .ZN(n1686) );
  INV_X1 U2298 ( .A(n1392), .ZN(n1393) );
  NAND2_X1 U2299 ( .A1(n1392), .A2(n1813), .ZN(n1662) );
  NAND2_X1 U2300 ( .A1(n1557), .A2(n1513), .ZN(n1416) );
  XNOR2_X1 U2301 ( .A(n1226), .B(n1682), .ZN(n1943) );
  NAND2_X1 U2302 ( .A1(n1411), .A2(n1511), .ZN(n1557) );
  OAI21_X1 U2303 ( .B1(n1434), .B2(S2_IMM_B), .A(n1388), .ZN(n1389) );
  NAND2_X1 U2304 ( .A1(S2_IMM_B), .A2(B[2]), .ZN(n1388) );
  OAI21_X1 U2305 ( .B1(n1433), .B2(S2_IMM_B), .A(n1395), .ZN(n1396) );
  NOR2_X1 U2306 ( .A1(n1397), .A2(S2_IMM_B), .ZN(n1401) );
  NAND2_X1 U2307 ( .A1(S2_IMM_B), .A2(B[1]), .ZN(n1395) );
  OAI22_X1 U2308 ( .A1(n1185), .A2(n2309), .B1(n1352), .B2(n2171), .ZN(n1489)
         );
  NOR2_X1 U2309 ( .A1(n1185), .A2(n1990), .ZN(n1467) );
  NOR2_X1 U2310 ( .A1(n1185), .A2(n2006), .ZN(n1450) );
  NOR2_X1 U2311 ( .A1(n1185), .A2(n2241), .ZN(n1929) );
  NOR2_X1 U2312 ( .A1(n1185), .A2(n1955), .ZN(n1430) );
  NOR2_X1 U2313 ( .A1(n1185), .A2(n1973), .ZN(n1437) );
  NAND2_X1 U2314 ( .A1(n1185), .A2(n1441), .ZN(n1494) );
  NAND2_X1 U2315 ( .A1(n1142), .A2(n1352), .ZN(n1949) );
  INV_X1 U2316 ( .A(n1185), .ZN(n1948) );
  NOR2_X1 U2317 ( .A1(n1352), .A2(n2307), .ZN(n2100) );
  INV_X1 U2318 ( .A(n2098), .ZN(n1953) );
  INV_X1 U2319 ( .A(n2244), .ZN(n1364) );
  MUX2_X1 U2320 ( .A(IMM[5]), .B(B[5]), .S(S2_IMM_B), .Z(n1827) );
  MUX2_X1 U2321 ( .A(A[5]), .B(NPC1[5]), .S(S1_A_NPC), .Z(n1897) );
  MUX2_X1 U2322 ( .A(n1384), .B(n2351), .S(S2_IMM_B), .Z(n2098) );
  MUX2_X1 U2323 ( .A(A[3]), .B(NPC1[3]), .S(S1_A_NPC), .Z(n1813) );
  MUX2_X1 U2324 ( .A(n1391), .B(n1390), .S(S1_A_NPC), .Z(n2131) );
  MUX2_X1 U2325 ( .A(A[1]), .B(NPC1[1]), .S(S1_A_NPC), .Z(n1781) );
  NAND3_X1 U2326 ( .A1(n1404), .A2(n1377), .A3(n1403), .ZN(n1405) );
  NAND3_X1 U2327 ( .A1(n1660), .A2(n1662), .A3(n1659), .ZN(n1484) );
  NAND3_X1 U2328 ( .A1(n1510), .A2(n1484), .A3(n1485), .ZN(n1411) );
  MUX2_X1 U2329 ( .A(A[6]), .B(NPC1[6]), .S(S1_A_NPC), .Z(n2061) );
  MUX2_X1 U2330 ( .A(IMM[7]), .B(B[7]), .S(n1382), .Z(n1540) );
  MUX2_X1 U2331 ( .A(n1414), .B(n1413), .S(S1_A_NPC), .Z(n2240) );
  MUX2_X1 U2332 ( .A(IMM[9]), .B(B[9]), .S(S2_IMM_B), .Z(n1848) );
  MUX2_X1 U2333 ( .A(A[9]), .B(NPC1[9]), .S(S1_A_NPC), .Z(n1971) );
  MUX2_X1 U2334 ( .A(IMM[8]), .B(B[8]), .S(S2_IMM_B), .Z(n1834) );
  MUX2_X1 U2335 ( .A(A[8]), .B(NPC1[8]), .S(S1_A_NPC), .Z(n1951) );
  MUX2_X1 U2336 ( .A(IMM[10]), .B(B[10]), .S(S2_IMM_B), .Z(n1863) );
  MUX2_X1 U2337 ( .A(A[10]), .B(NPC1[10]), .S(S1_A_NPC), .Z(n1989) );
  MUX2_X1 U2338 ( .A(IMM[11]), .B(B[11]), .S(n1382), .Z(n1478) );
  MUX2_X1 U2339 ( .A(A[11]), .B(NPC1[11]), .S(S1_A_NPC), .Z(n2004) );
  MUX2_X1 U2340 ( .A(n1428), .B(n1427), .S(n1148), .Z(n2243) );
  MUX2_X1 U2341 ( .A(A[16]), .B(NPC1[16]), .S(n1148), .Z(n2103) );
  MUX2_X1 U2342 ( .A(A[0]), .B(NPC1[0]), .S(n1383), .Z(n1760) );
  MUX2_X1 U2343 ( .A(n1433), .B(n2326), .S(n1173), .Z(n1462) );
  MUX2_X1 U2344 ( .A(n1434), .B(n2337), .S(n1173), .Z(n1445) );
  MUX2_X1 U2345 ( .A(IMM[0]), .B(B[0]), .S(n1380), .Z(n1759) );
  MUX2_X1 U2346 ( .A(n1445), .B(n1462), .S(n1376), .Z(n1435) );
  MUX2_X1 U2347 ( .A(A[17]), .B(NPC1[17]), .S(n1148), .Z(n2123) );
  MUX2_X1 U2348 ( .A(n1443), .B(n1442), .S(S1_A_NPC), .Z(n1885) );
  MUX2_X1 U2349 ( .A(n1464), .B(n1463), .S(n1378), .Z(n1446) );
  MUX2_X1 U2350 ( .A(A[19]), .B(NPC1[19]), .S(n1148), .Z(n2150) );
  MUX2_X1 U2351 ( .A(A[13]), .B(NPC1[13]), .S(S1_A_NPC), .Z(n2038) );
  MUX2_X1 U2352 ( .A(n1460), .B(n1459), .S(n1383), .Z(n2246) );
  NAND3_X1 U2353 ( .A1(n1796), .A2(n1465), .A3(n1462), .ZN(n2217) );
  MUX2_X1 U2354 ( .A(n1464), .B(n1463), .S(n1376), .Z(n1466) );
  MUX2_X1 U2355 ( .A(A[18]), .B(NPC1[18]), .S(n1148), .Z(n2133) );
  MUX2_X1 U2356 ( .A(A[14]), .B(NPC1[14]), .S(n1383), .Z(n2059) );
  MUX2_X1 U2357 ( .A(n1782), .B(n1796), .S(n1376), .Z(n1471) );
  MUX2_X1 U2358 ( .A(n2169), .B(n2168), .S(n2004), .Z(n1480) );
  MUX2_X1 U2359 ( .A(n2171), .B(n2170), .S(n2004), .Z(n1479) );
  MUX2_X1 U2360 ( .A(n1480), .B(n1479), .S(n1195), .Z(n1481) );
  NAND3_X1 U2361 ( .A1(n1665), .A2(n2115), .A3(n1664), .ZN(n1509) );
  MUX2_X1 U2362 ( .A(n2170), .B(n2168), .S(n1352), .Z(n1491) );
  MUX2_X1 U2363 ( .A(n1491), .B(n1490), .S(n2182), .Z(n1508) );
  MUX2_X1 U2364 ( .A(n2232), .B(n2233), .S(n2061), .Z(n1520) );
  MUX2_X1 U2365 ( .A(n2236), .B(n2234), .S(n2061), .Z(n1519) );
  MUX2_X1 U2366 ( .A(n1520), .B(n1519), .S(n1150), .Z(n1521) );
  MUX2_X1 U2367 ( .A(n2168), .B(n2169), .S(n2240), .Z(n1542) );
  MUX2_X1 U2368 ( .A(n2170), .B(n2171), .S(n2240), .Z(n1541) );
  MUX2_X1 U2369 ( .A(n1542), .B(n1541), .S(n1162), .Z(n1543) );
  MUX2_X1 U2370 ( .A(IMM[31]), .B(B[31]), .S(n1380), .Z(n1617) );
  MUX2_X1 U2371 ( .A(IMM[24]), .B(B[24]), .S(n1381), .Z(n2117) );
  MUX2_X1 U2372 ( .A(A[24]), .B(NPC1[24]), .S(n1383), .Z(n2118) );
  MUX2_X1 U2373 ( .A(IMM[13]), .B(B[13]), .S(S2_IMM_B), .Z(n1904) );
  MUX2_X1 U2374 ( .A(IMM[12]), .B(B[12]), .S(S2_IMM_B), .Z(n1886) );
  NAND3_X1 U2375 ( .A1(n1641), .A2(n1640), .A3(n1685), .ZN(n1564) );
  MUX2_X1 U2376 ( .A(IMM[14]), .B(B[14]), .S(n1380), .Z(n1919) );
  MUX2_X1 U2377 ( .A(IMM[19]), .B(B[19]), .S(n1382), .Z(n2014) );
  MUX2_X1 U2378 ( .A(IMM[22]), .B(B[22]), .S(S2_IMM_B), .Z(n2072) );
  MUX2_X1 U2379 ( .A(A[22]), .B(NPC1[22]), .S(S1_A_NPC), .Z(n2209) );
  MUX2_X1 U2380 ( .A(IMM[20]), .B(B[20]), .S(n1380), .Z(n2032) );
  MUX2_X1 U2381 ( .A(A[20]), .B(NPC1[20]), .S(n1383), .Z(n2031) );
  MUX2_X1 U2382 ( .A(IMM[21]), .B(B[21]), .S(n1160), .Z(n2050) );
  MUX2_X1 U2383 ( .A(A[21]), .B(NPC1[21]), .S(n1148), .Z(n2194) );
  MUX2_X1 U2384 ( .A(IMM[23]), .B(B[23]), .S(n1380), .Z(n2078) );
  MUX2_X1 U2385 ( .A(n1575), .B(n1574), .S(n1383), .Z(n2241) );
  MUX2_X1 U2386 ( .A(IMM[15]), .B(B[15]), .S(n1381), .Z(n1938) );
  NAND3_X1 U2387 ( .A1(n1631), .A2(n1589), .A3(n1743), .ZN(n1590) );
  MUX2_X1 U2388 ( .A(IMM[25]), .B(B[25]), .S(n1380), .Z(n2119) );
  MUX2_X1 U2389 ( .A(A[25]), .B(NPC1[25]), .S(n1383), .Z(n2120) );
  MUX2_X1 U2390 ( .A(IMM[26]), .B(B[26]), .S(n1168), .Z(n2127) );
  MUX2_X1 U2391 ( .A(A[26]), .B(NPC1[26]), .S(n1383), .Z(n2128) );
  MUX2_X1 U2392 ( .A(IMM[27]), .B(B[27]), .S(n1173), .Z(n2165) );
  MUX2_X1 U2393 ( .A(n1603), .B(n1602), .S(n1383), .Z(n2149) );
  MUX2_X1 U2394 ( .A(IMM[28]), .B(B[28]), .S(n1381), .Z(n2172) );
  MUX2_X1 U2395 ( .A(A[28]), .B(NPC1[28]), .S(n1383), .Z(n2178) );
  MUX2_X1 U2396 ( .A(IMM[29]), .B(B[29]), .S(n1173), .Z(n2205) );
  MUX2_X1 U2397 ( .A(A[29]), .B(NPC1[29]), .S(n1383), .Z(n2204) );
  MUX2_X1 U2398 ( .A(IMM[30]), .B(B[30]), .S(n1381), .Z(n2229) );
  MUX2_X1 U2399 ( .A(A[30]), .B(NPC1[30]), .S(n1383), .Z(n2228) );
  NAND3_X1 U2400 ( .A1(n1801), .A2(n1758), .A3(n1787), .ZN(n1663) );
  MUX2_X1 U2401 ( .A(n2232), .B(n2236), .S(n1759), .Z(n1762) );
  MUX2_X1 U2402 ( .A(n2233), .B(n2234), .S(n1759), .Z(n1761) );
  MUX2_X1 U2403 ( .A(n1762), .B(n1761), .S(n1760), .Z(n1763) );
  MUX2_X1 U2404 ( .A(n2169), .B(n2168), .S(n1200), .Z(n1784) );
  MUX2_X1 U2405 ( .A(n2171), .B(n2170), .S(n1200), .Z(n1783) );
  MUX2_X1 U2406 ( .A(n1784), .B(n1783), .S(n1782), .Z(n1785) );
  NAND3_X1 U2407 ( .A1(n1359), .A2(n1375), .A3(n1165), .ZN(n1793) );
  MUX2_X1 U2408 ( .A(n2168), .B(n2169), .S(n2131), .Z(n1798) );
  MUX2_X1 U2409 ( .A(n2170), .B(n2171), .S(n2131), .Z(n1797) );
  MUX2_X1 U2410 ( .A(n1798), .B(n1797), .S(n1796), .Z(n1799) );
  MUX2_X1 U2411 ( .A(n2169), .B(n2168), .S(n1165), .Z(n1815) );
  MUX2_X1 U2412 ( .A(n2171), .B(n2170), .S(n1813), .Z(n1814) );
  MUX2_X1 U2413 ( .A(n1815), .B(n1814), .S(n1235), .Z(n1816) );
  NAND3_X1 U2414 ( .A1(n1826), .A2(n1825), .A3(n1824), .ZN(n1831) );
  MUX2_X1 U2415 ( .A(n2232), .B(n2233), .S(n1897), .Z(n1829) );
  MUX2_X1 U2416 ( .A(n2236), .B(n2234), .S(n1897), .Z(n1828) );
  MUX2_X1 U2417 ( .A(n1829), .B(n1828), .S(n1192), .Z(n1830) );
  MUX2_X1 U2418 ( .A(n2169), .B(n2168), .S(n1951), .Z(n1836) );
  MUX2_X1 U2419 ( .A(n2171), .B(n2170), .S(n1951), .Z(n1835) );
  MUX2_X1 U2420 ( .A(n1836), .B(n1835), .S(n1193), .Z(n1846) );
  MUX2_X1 U2421 ( .A(n2169), .B(n2168), .S(n1971), .Z(n1850) );
  MUX2_X1 U2422 ( .A(n2171), .B(n2170), .S(n1971), .Z(n1849) );
  MUX2_X1 U2423 ( .A(n1850), .B(n1849), .S(n1848), .Z(n1861) );
  MUX2_X1 U2424 ( .A(n2169), .B(n2168), .S(n1989), .Z(n1865) );
  MUX2_X1 U2425 ( .A(n2171), .B(n2170), .S(n1989), .Z(n1864) );
  MUX2_X1 U2426 ( .A(n1865), .B(n1864), .S(n1863), .Z(n1875) );
  MUX2_X1 U2427 ( .A(n2168), .B(n2169), .S(n1885), .Z(n1888) );
  MUX2_X1 U2428 ( .A(n2170), .B(n2171), .S(n1885), .Z(n1887) );
  MUX2_X1 U2429 ( .A(n1888), .B(n1887), .S(n1886), .Z(n1889) );
  NAND3_X1 U2430 ( .A1(n1903), .A2(n1902), .A3(n2115), .ZN(n1908) );
  MUX2_X1 U2431 ( .A(n2169), .B(n2168), .S(n2038), .Z(n1906) );
  MUX2_X1 U2432 ( .A(n2171), .B(n2170), .S(n2038), .Z(n1905) );
  MUX2_X1 U2433 ( .A(n1906), .B(n1905), .S(n1904), .Z(n1907) );
  MUX2_X1 U2434 ( .A(n2169), .B(n2168), .S(n2059), .Z(n1921) );
  MUX2_X1 U2435 ( .A(n2171), .B(n2170), .S(n2059), .Z(n1920) );
  MUX2_X1 U2436 ( .A(n1921), .B(n1920), .S(n1919), .Z(n1922) );
  MUX2_X1 U2437 ( .A(n2168), .B(n2169), .S(n2246), .Z(n1940) );
  MUX2_X1 U2438 ( .A(n2170), .B(n2171), .S(n2246), .Z(n1939) );
  MUX2_X1 U2439 ( .A(n1940), .B(n1939), .S(n1938), .Z(n1941) );
  MUX2_X1 U2440 ( .A(n2169), .B(n2168), .S(n2103), .Z(n1946) );
  MUX2_X1 U2441 ( .A(n2171), .B(n2170), .S(n2103), .Z(n1945) );
  MUX2_X1 U2442 ( .A(n1946), .B(n1945), .S(n1151), .Z(n1966) );
  MUX2_X1 U2443 ( .A(n2169), .B(n2168), .S(n2123), .Z(n1970) );
  MUX2_X1 U2444 ( .A(n2171), .B(n2170), .S(n2123), .Z(n1969) );
  MUX2_X1 U2445 ( .A(n1970), .B(n1969), .S(n1197), .Z(n1984) );
  MUX2_X1 U2446 ( .A(n2169), .B(n2168), .S(n2133), .Z(n1988) );
  MUX2_X1 U2447 ( .A(n2171), .B(n2170), .S(n2133), .Z(n1987) );
  MUX2_X1 U2448 ( .A(n1988), .B(n1987), .S(n1156), .Z(n2000) );
  MUX2_X1 U2449 ( .A(n2169), .B(n2168), .S(n2150), .Z(n2016) );
  MUX2_X1 U2450 ( .A(n2171), .B(n2170), .S(n2150), .Z(n2015) );
  MUX2_X1 U2451 ( .A(n2016), .B(n2015), .S(n1190), .Z(n2017) );
  MUX2_X1 U2452 ( .A(n2169), .B(n2168), .S(n2031), .Z(n2034) );
  MUX2_X1 U2453 ( .A(n2171), .B(n2170), .S(n2031), .Z(n2033) );
  MUX2_X1 U2454 ( .A(n2034), .B(n2033), .S(n2032), .Z(n2035) );
  MUX2_X1 U2455 ( .A(n2169), .B(n2168), .S(n2194), .Z(n2052) );
  MUX2_X1 U2456 ( .A(n2171), .B(n2170), .S(n2194), .Z(n2051) );
  MUX2_X1 U2457 ( .A(n2052), .B(n2051), .S(n2050), .Z(n2053) );
  MUX2_X1 U2458 ( .A(n2169), .B(n2168), .S(n2209), .Z(n2074) );
  MUX2_X1 U2459 ( .A(n2171), .B(n2170), .S(n2209), .Z(n2073) );
  MUX2_X1 U2460 ( .A(n2074), .B(n2073), .S(n2072), .Z(n2075) );
  MUX2_X1 U2461 ( .A(n2168), .B(n2169), .S(n2241), .Z(n2080) );
  MUX2_X1 U2462 ( .A(n2170), .B(n2171), .S(n2241), .Z(n2079) );
  MUX2_X1 U2463 ( .A(n2080), .B(n2079), .S(n2078), .Z(n2095) );
  MUX2_X1 U2464 ( .A(n2169), .B(n2171), .S(n2127), .Z(n2130) );
  MUX2_X1 U2465 ( .A(n2168), .B(n2170), .S(n2127), .Z(n2129) );
  MUX2_X1 U2466 ( .A(n2130), .B(n2129), .S(n2128), .Z(n2143) );
  MUX2_X1 U2467 ( .A(n2234), .B(n2236), .S(n2149), .Z(n2164) );
  MUX2_X1 U2468 ( .A(n2233), .B(n2232), .S(n2243), .Z(n2273) );
  NOR2_X1 U2469 ( .A1(ALU_OPCODE[1]), .A2(n1376), .ZN(n2308) );
  NAND2_X1 U2470 ( .A1(ALU_OPCODE[4]), .A2(ALU_OPCODE[5]), .ZN(n2309) );
  INV_X1 U2471 ( .A(n2308), .ZN(n2307) );
  NOR4_X1 U2472 ( .A1(A[28]), .A2(A[30]), .A3(A[29]), .A4(A[15]), .ZN(n2313)
         );
  NOR4_X1 U2473 ( .A1(A[31]), .A2(A[27]), .A3(A[26]), .A4(A[25]), .ZN(n2312)
         );
  NOR4_X1 U2474 ( .A1(A[17]), .A2(A[19]), .A3(A[23]), .A4(A[20]), .ZN(n2311)
         );
  NOR4_X1 U2475 ( .A1(A[14]), .A2(A[13]), .A3(A[16]), .A4(A[18]), .ZN(n2310)
         );
  NAND4_X1 U2476 ( .A1(n2313), .A2(n2312), .A3(n2311), .A4(n2310), .ZN(n2319)
         );
  NOR4_X1 U2477 ( .A1(A[10]), .A2(A[5]), .A3(A[4]), .A4(A[0]), .ZN(n2317) );
  NOR4_X1 U2478 ( .A1(A[21]), .A2(A[22]), .A3(A[24]), .A4(A[6]), .ZN(n2316) );
  NOR4_X1 U2479 ( .A1(A[12]), .A2(A[2]), .A3(A[3]), .A4(A[1]), .ZN(n2315) );
  NOR4_X1 U2480 ( .A1(A[11]), .A2(A[9]), .A3(A[7]), .A4(A[8]), .ZN(n2314) );
  NAND4_X1 U2481 ( .A1(n2317), .A2(n2316), .A3(n2315), .A4(n2314), .ZN(n2318)
         );
  OAI21_X1 U2482 ( .B1(n2319), .B2(n2318), .A(JUMP_EN[1]), .ZN(n2320) );
  OAI22_X1 U2483 ( .A1(n2321), .A2(n1180), .B1(\COMP_REGN_ALUOUT/ffi_11/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_11/n5 ) );
  OAI22_X1 U2484 ( .A1(n2322), .A2(n1370), .B1(\COMP_REGN_ALUOUT/ffi_4/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_4/n5 ) );
  OAI22_X1 U2485 ( .A1(n2323), .A2(n1370), .B1(\COMP_REGN_ALUOUT/ffi_6/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_6/n5 ) );
  OAI22_X1 U2486 ( .A1(n2324), .A2(n1370), .B1(\COMP_REGN_ALUOUT/ffi_7/n4 ), 
        .B2(n1366), .ZN(\COMP_REGN_ALUOUT/ffi_7/n5 ) );
  INV_X1 U2487 ( .A(B[0]), .ZN(n2325) );
  OAI22_X1 U2488 ( .A1(\COMP_REGN_BOUT/ffi_0/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2325), .ZN(\COMP_REGN_BOUT/ffi_0/n5 ) );
  INV_X1 U2489 ( .A(B[1]), .ZN(n2326) );
  OAI22_X1 U2490 ( .A1(\COMP_REGN_BOUT/ffi_1/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2326), .ZN(\COMP_REGN_BOUT/ffi_1/n5 ) );
  INV_X1 U2491 ( .A(B[10]), .ZN(n2327) );
  OAI22_X1 U2492 ( .A1(\COMP_REGN_BOUT/ffi_10/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2327), .ZN(\COMP_REGN_BOUT/ffi_10/n5 ) );
  INV_X1 U2493 ( .A(B[11]), .ZN(n2328) );
  OAI22_X1 U2494 ( .A1(\COMP_REGN_BOUT/ffi_11/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2328), .ZN(\COMP_REGN_BOUT/ffi_11/n5 ) );
  INV_X1 U2495 ( .A(B[12]), .ZN(n2329) );
  OAI22_X1 U2496 ( .A1(\COMP_REGN_BOUT/ffi_12/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2329), .ZN(\COMP_REGN_BOUT/ffi_12/n5 ) );
  INV_X1 U2497 ( .A(B[13]), .ZN(n2330) );
  OAI22_X1 U2498 ( .A1(\COMP_REGN_BOUT/ffi_13/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2330), .ZN(\COMP_REGN_BOUT/ffi_13/n5 ) );
  INV_X1 U2499 ( .A(B[14]), .ZN(n2331) );
  OAI22_X1 U2500 ( .A1(\COMP_REGN_BOUT/ffi_14/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2331), .ZN(\COMP_REGN_BOUT/ffi_14/n5 ) );
  INV_X1 U2501 ( .A(B[15]), .ZN(n2332) );
  OAI22_X1 U2502 ( .A1(\COMP_REGN_BOUT/ffi_15/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2332), .ZN(\COMP_REGN_BOUT/ffi_15/n5 ) );
  INV_X1 U2503 ( .A(B[16]), .ZN(n2333) );
  OAI22_X1 U2504 ( .A1(\COMP_REGN_BOUT/ffi_16/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2333), .ZN(\COMP_REGN_BOUT/ffi_16/n5 ) );
  INV_X1 U2505 ( .A(B[17]), .ZN(n2334) );
  OAI22_X1 U2506 ( .A1(\COMP_REGN_BOUT/ffi_17/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2334), .ZN(\COMP_REGN_BOUT/ffi_17/n5 ) );
  INV_X1 U2507 ( .A(B[18]), .ZN(n2335) );
  OAI22_X1 U2508 ( .A1(\COMP_REGN_BOUT/ffi_18/n4 ), .A2(n1366), .B1(n1370), 
        .B2(n2335), .ZN(\COMP_REGN_BOUT/ffi_18/n5 ) );
  INV_X1 U2509 ( .A(B[19]), .ZN(n2336) );
  OAI22_X1 U2510 ( .A1(\COMP_REGN_BOUT/ffi_19/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2336), .ZN(\COMP_REGN_BOUT/ffi_19/n5 ) );
  INV_X1 U2511 ( .A(B[2]), .ZN(n2337) );
  OAI22_X1 U2512 ( .A1(\COMP_REGN_BOUT/ffi_2/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2337), .ZN(\COMP_REGN_BOUT/ffi_2/n5 ) );
  INV_X1 U2513 ( .A(B[20]), .ZN(n2338) );
  OAI22_X1 U2514 ( .A1(\COMP_REGN_BOUT/ffi_20/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2338), .ZN(\COMP_REGN_BOUT/ffi_20/n5 ) );
  INV_X1 U2515 ( .A(B[21]), .ZN(n2339) );
  OAI22_X1 U2516 ( .A1(\COMP_REGN_BOUT/ffi_21/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2339), .ZN(\COMP_REGN_BOUT/ffi_21/n5 ) );
  INV_X1 U2517 ( .A(B[22]), .ZN(n2340) );
  OAI22_X1 U2518 ( .A1(\COMP_REGN_BOUT/ffi_22/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2340), .ZN(\COMP_REGN_BOUT/ffi_22/n5 ) );
  INV_X1 U2519 ( .A(B[23]), .ZN(n2341) );
  OAI22_X1 U2520 ( .A1(\COMP_REGN_BOUT/ffi_23/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2341), .ZN(\COMP_REGN_BOUT/ffi_23/n5 ) );
  INV_X1 U2521 ( .A(B[24]), .ZN(n2342) );
  OAI22_X1 U2522 ( .A1(\COMP_REGN_BOUT/ffi_24/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2342), .ZN(\COMP_REGN_BOUT/ffi_24/n5 ) );
  INV_X1 U2523 ( .A(B[25]), .ZN(n2343) );
  OAI22_X1 U2524 ( .A1(\COMP_REGN_BOUT/ffi_25/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2343), .ZN(\COMP_REGN_BOUT/ffi_25/n5 ) );
  INV_X1 U2525 ( .A(B[26]), .ZN(n2344) );
  OAI22_X1 U2526 ( .A1(\COMP_REGN_BOUT/ffi_26/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2344), .ZN(\COMP_REGN_BOUT/ffi_26/n5 ) );
  INV_X1 U2527 ( .A(B[27]), .ZN(n2345) );
  OAI22_X1 U2528 ( .A1(\COMP_REGN_BOUT/ffi_27/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2345), .ZN(\COMP_REGN_BOUT/ffi_27/n5 ) );
  INV_X1 U2529 ( .A(B[28]), .ZN(n2346) );
  OAI22_X1 U2530 ( .A1(\COMP_REGN_BOUT/ffi_28/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2346), .ZN(\COMP_REGN_BOUT/ffi_28/n5 ) );
  INV_X1 U2531 ( .A(B[29]), .ZN(n2347) );
  OAI22_X1 U2532 ( .A1(\COMP_REGN_BOUT/ffi_29/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2347), .ZN(\COMP_REGN_BOUT/ffi_29/n5 ) );
  INV_X1 U2533 ( .A(B[3]), .ZN(n2348) );
  OAI22_X1 U2534 ( .A1(\COMP_REGN_BOUT/ffi_3/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2348), .ZN(\COMP_REGN_BOUT/ffi_3/n5 ) );
  INV_X1 U2535 ( .A(B[30]), .ZN(n2349) );
  OAI22_X1 U2536 ( .A1(\COMP_REGN_BOUT/ffi_30/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2349), .ZN(\COMP_REGN_BOUT/ffi_30/n5 ) );
  INV_X1 U2537 ( .A(B[31]), .ZN(n2350) );
  OAI22_X1 U2538 ( .A1(\COMP_REGN_BOUT/ffi_31/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2350), .ZN(\COMP_REGN_BOUT/ffi_31/n5 ) );
  INV_X1 U2539 ( .A(B[4]), .ZN(n2351) );
  OAI22_X1 U2540 ( .A1(\COMP_REGN_BOUT/ffi_4/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2351), .ZN(\COMP_REGN_BOUT/ffi_4/n5 ) );
  INV_X1 U2541 ( .A(B[5]), .ZN(n2352) );
  OAI22_X1 U2542 ( .A1(\COMP_REGN_BOUT/ffi_5/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2352), .ZN(\COMP_REGN_BOUT/ffi_5/n5 ) );
  INV_X1 U2543 ( .A(B[6]), .ZN(n2353) );
  OAI22_X1 U2544 ( .A1(\COMP_REGN_BOUT/ffi_6/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2353), .ZN(\COMP_REGN_BOUT/ffi_6/n5 ) );
  INV_X1 U2545 ( .A(B[7]), .ZN(n2354) );
  OAI22_X1 U2546 ( .A1(\COMP_REGN_BOUT/ffi_7/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2354), .ZN(\COMP_REGN_BOUT/ffi_7/n5 ) );
  INV_X1 U2547 ( .A(B[8]), .ZN(n2355) );
  OAI22_X1 U2548 ( .A1(\COMP_REGN_BOUT/ffi_8/n4 ), .A2(n1367), .B1(n1369), 
        .B2(n2355), .ZN(\COMP_REGN_BOUT/ffi_8/n5 ) );
  INV_X1 U2549 ( .A(B[9]), .ZN(n2356) );
  OAI22_X1 U2550 ( .A1(\COMP_REGN_BOUT/ffi_9/n4 ), .A2(n1367), .B1(n1370), 
        .B2(n2356), .ZN(\COMP_REGN_BOUT/ffi_9/n5 ) );
  AOI22_X1 U2551 ( .A1(n1186), .A2(RD1[0]), .B1(n1187), .B2(RD2_OUT_REGN[0]), 
        .ZN(n2357) );
  AOI22_X1 U2552 ( .A1(n1186), .A2(RD1[1]), .B1(n1187), .B2(RD2_OUT_REGN[1]), 
        .ZN(n2358) );
  AOI22_X1 U2553 ( .A1(n1186), .A2(RD1[2]), .B1(n1187), .B2(RD2_OUT_REGN[2]), 
        .ZN(n2359) );
  AOI22_X1 U2554 ( .A1(n1186), .A2(RD1[3]), .B1(n1187), .B2(RD2_OUT_REGN[3]), 
        .ZN(n2360) );
  AOI22_X1 U2555 ( .A1(n1186), .A2(RD1[4]), .B1(n1187), .B2(RD2_OUT_REGN[4]), 
        .ZN(n2361) );
  AOI22_X1 U2556 ( .A1(n1186), .A2(NPC1[0]), .B1(n1187), .B2(NPC2[0]), .ZN(
        n2362) );
  AOI22_X1 U2557 ( .A1(n1186), .A2(NPC1[1]), .B1(n1187), .B2(NPC2[1]), .ZN(
        n2363) );
  AOI22_X1 U2558 ( .A1(n1186), .A2(NPC1[2]), .B1(n1187), .B2(NPC2[2]), .ZN(
        n2364) );
  AOI22_X1 U2559 ( .A1(n1186), .A2(NPC1[3]), .B1(n1187), .B2(NPC2[3]), .ZN(
        n2365) );
  AOI22_X1 U2560 ( .A1(n1186), .A2(NPC1[4]), .B1(n1187), .B2(NPC2[4]), .ZN(
        n2366) );
  AOI22_X1 U2561 ( .A1(n1186), .A2(NPC1[5]), .B1(n1187), .B2(NPC2[5]), .ZN(
        n2367) );
  AOI22_X1 U2562 ( .A1(n1186), .A2(NPC1[6]), .B1(n1187), .B2(NPC2[6]), .ZN(
        n2368) );
  AOI22_X1 U2563 ( .A1(n1186), .A2(NPC1[7]), .B1(n1187), .B2(NPC2[7]), .ZN(
        n2369) );
  AOI22_X1 U2564 ( .A1(n1186), .A2(NPC1[8]), .B1(n1187), .B2(NPC2[8]), .ZN(
        n2370) );
  AOI22_X1 U2565 ( .A1(n1186), .A2(NPC1[9]), .B1(n1187), .B2(NPC2[9]), .ZN(
        n2371) );
  AOI22_X1 U2566 ( .A1(n1186), .A2(NPC1[10]), .B1(n1187), .B2(NPC2[10]), .ZN(
        n2372) );
  AOI22_X1 U2567 ( .A1(n1186), .A2(NPC1[11]), .B1(n1187), .B2(NPC2[11]), .ZN(
        n2373) );
  AOI22_X1 U2568 ( .A1(n1186), .A2(NPC1[12]), .B1(n1187), .B2(NPC2[12]), .ZN(
        n2374) );
  AOI22_X1 U2569 ( .A1(n1186), .A2(NPC1[13]), .B1(n1187), .B2(NPC2[13]), .ZN(
        n2375) );
  AOI22_X1 U2570 ( .A1(n1186), .A2(NPC1[14]), .B1(n1187), .B2(NPC2[14]), .ZN(
        n2376) );
  AOI22_X1 U2571 ( .A1(n1186), .A2(NPC1[15]), .B1(n1187), .B2(NPC2[15]), .ZN(
        n2377) );
  AOI22_X1 U2572 ( .A1(n1186), .A2(NPC1[16]), .B1(n1187), .B2(NPC2[16]), .ZN(
        n2378) );
  AOI22_X1 U2573 ( .A1(n1186), .A2(NPC1[17]), .B1(n1187), .B2(NPC2[17]), .ZN(
        n2379) );
  AOI22_X1 U2574 ( .A1(n1186), .A2(NPC1[18]), .B1(n1187), .B2(NPC2[18]), .ZN(
        n2380) );
  AOI22_X1 U2575 ( .A1(n1186), .A2(NPC1[19]), .B1(n1187), .B2(NPC2[19]), .ZN(
        n2381) );
  AOI22_X1 U2576 ( .A1(n1186), .A2(NPC1[20]), .B1(n1187), .B2(NPC2[20]), .ZN(
        n2382) );
  AOI22_X1 U2577 ( .A1(n1186), .A2(NPC1[21]), .B1(n1187), .B2(NPC2[21]), .ZN(
        n2383) );
  AOI22_X1 U2578 ( .A1(n1186), .A2(NPC1[22]), .B1(n1187), .B2(NPC2[22]), .ZN(
        n2384) );
  AOI22_X1 U2579 ( .A1(n1186), .A2(NPC1[23]), .B1(n1187), .B2(NPC2[23]), .ZN(
        n2385) );
  AOI22_X1 U2580 ( .A1(n1186), .A2(NPC1[24]), .B1(n1187), .B2(NPC2[24]), .ZN(
        n2386) );
  AOI22_X1 U2581 ( .A1(n1186), .A2(NPC1[25]), .B1(n1187), .B2(NPC2[25]), .ZN(
        n2387) );
  AOI22_X1 U2582 ( .A1(n1186), .A2(NPC1[26]), .B1(n1187), .B2(NPC2[26]), .ZN(
        n2388) );
  AOI22_X1 U2583 ( .A1(n1186), .A2(NPC1[27]), .B1(n1187), .B2(NPC2[27]), .ZN(
        n2389) );
  AOI22_X1 U2584 ( .A1(n1186), .A2(NPC1[28]), .B1(n1187), .B2(NPC2[28]), .ZN(
        n2390) );
  AOI22_X1 U2585 ( .A1(n1186), .A2(NPC1[29]), .B1(n1187), .B2(NPC2[29]), .ZN(
        n2391) );
  AOI22_X1 U2586 ( .A1(n1186), .A2(NPC1[30]), .B1(n1187), .B2(NPC2[30]), .ZN(
        n2392) );
  AOI22_X1 U2587 ( .A1(n1186), .A2(NPC1[31]), .B1(n2305), .B2(NPC2[31]), .ZN(
        n2393) );
endmodule


module dlx ( RST, CLK );
  input RST, CLK;
  wire   jump, \unit_control/n418 , \unit_control/n400 , \unit_control/n399 ,
         \unit_control/n398 , \unit_control/n393 , \unit_control/n392 ,
         \unit_control/n391 , \unit_control/n390 , \unit_control/n389 ,
         \unit_control/n387 , \unit_control/n386 , \unit_control/n385 ,
         \unit_control/n383 , \unit_control/n382 , \unit_control/n381 ,
         \unit_control/n379 , \unit_control/n378 , \unit_control/n373 ,
         \unit_control/n266 , \unit_control/uut_third_stage/ffi_11/n5 ,
         \unit_control/uut_third_stage/ffi_10/n5 ,
         \unit_control/uut_third_stage/ffi_9/n6 ,
         \unit_control/uut_fourth_stage/ffi_6/n6 ,
         \unit_control/uut_fourth_stage/ffi_3/n6 ,
         \unit_control/uut_second_stage/ffi_17/n5 ,
         \unit_control/uut_second_stage/ffi_15/n5 ,
         \unit_control/uut_second_stage/ffi_14/n5 ,
         \unit_control/uut_second_stage/ffi_13/n5 ,
         \unit_control/uut_second_stage/ffi_12/n5 ,
         \unit_control/uut_second_stage/ffi_11/n5 ,
         \unit_control/uut_second_stage/ffi_10/n5 ,
         \unit_control/uut_second_stage/ffi_9/n5 ,
         \unit_control/uut_second_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_15/n5 ,
         \unit_control/uut_third_stage/ffi_14/n5 ,
         \unit_control/uut_third_stage/ffi_13/n5 ,
         \unit_control/uut_third_stage/ffi_7/n5 ,
         \unit_control/uut_third_stage/ffi_6/n5 ,
         \unit_control/uut_third_stage/ffi_5/n5 ,
         \unit_control/uut_third_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_3/n5 ,
         \unit_control/uut_fourth_stage/ffi_7/n5 ,
         \unit_control/uut_fourth_stage/ffi_5/n5 ,
         \unit_control/uut_fourth_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_12/n5 ,
         \unit_control/uut_third_stage/ffi_12/n2 ,
         \unit_control/uut_third_stage/ffi_17/n6 ,
         \unit_control/uut_third_stage/ffi_17/n2 ,
         \unit_control/uut_third_stage/ffi_19/n6 ,
         \unit_control/uut_third_stage/ffi_19/n2 ,
         \unit_control/uut_second_stage/ffi_24/n5 ,
         \unit_control/next_state[1] , \unit_control/next_state[0] ,
         \unit_fetch/n682 , \unit_fetch/n674 , \unit_fetch/n462 ,
         \unit_fetch/n447 , \unit_fetch/n329 ,
         \unit_fetch/unit_programCounter/ffi_30/n5 ,
         \unit_fetch/unit_programCounter/ffi_29/n5 ,
         \unit_fetch/unit_programCounter/ffi_28/n5 ,
         \unit_fetch/unit_programCounter/ffi_27/n5 ,
         \unit_fetch/unit_programCounter/ffi_26/n5 ,
         \unit_fetch/unit_programCounter/ffi_25/n5 ,
         \unit_fetch/unit_programCounter/ffi_24/n5 ,
         \unit_fetch/unit_programCounter/ffi_23/n5 ,
         \unit_fetch/unit_programCounter/ffi_22/n5 ,
         \unit_fetch/unit_programCounter/ffi_21/n5 ,
         \unit_fetch/unit_programCounter/ffi_20/n5 ,
         \unit_fetch/unit_programCounter/ffi_19/n5 ,
         \unit_fetch/unit_programCounter/ffi_18/n5 ,
         \unit_fetch/unit_programCounter/ffi_17/n5 ,
         \unit_fetch/unit_programCounter/ffi_16/n5 ,
         \unit_fetch/unit_programCounter/ffi_15/n5 ,
         \unit_fetch/unit_programCounter/ffi_14/n5 ,
         \unit_fetch/unit_programCounter/ffi_13/n5 ,
         \unit_fetch/unit_programCounter/ffi_12/n5 ,
         \unit_fetch/unit_programCounter/ffi_11/n5 ,
         \unit_fetch/unit_programCounter/ffi_10/n5 ,
         \unit_fetch/unit_programCounter/ffi_9/n5 ,
         \unit_fetch/unit_programCounter/ffi_8/n5 ,
         \unit_fetch/unit_programCounter/ffi_7/n5 ,
         \unit_fetch/unit_programCounter/ffi_6/n5 ,
         \unit_fetch/unit_programCounter/ffi_5/n5 ,
         \unit_fetch/unit_programCounter/ffi_4/n5 ,
         \unit_fetch/unit_programCounter/ffi_3/n5 ,
         \unit_fetch/unit_programCounter/ffi_2/n5 ,
         \unit_fetch/unit_programCounter/ffi_1/n5 ,
         \unit_fetch/unit_programCounter/ffi_0/n5 ,
         \unit_fetch/unit_npcregister/ffi_31/n5 ,
         \unit_fetch/unit_npcregister/ffi_30/n5 ,
         \unit_fetch/unit_npcregister/ffi_29/n5 ,
         \unit_fetch/unit_npcregister/ffi_28/n5 ,
         \unit_fetch/unit_npcregister/ffi_27/n5 ,
         \unit_fetch/unit_npcregister/ffi_26/n5 ,
         \unit_fetch/unit_npcregister/ffi_25/n5 ,
         \unit_fetch/unit_npcregister/ffi_24/n5 ,
         \unit_fetch/unit_npcregister/ffi_23/n5 ,
         \unit_fetch/unit_npcregister/ffi_22/n5 ,
         \unit_fetch/unit_npcregister/ffi_21/n5 ,
         \unit_fetch/unit_npcregister/ffi_20/n5 ,
         \unit_fetch/unit_npcregister/ffi_19/n5 ,
         \unit_fetch/unit_npcregister/ffi_18/n5 ,
         \unit_fetch/unit_npcregister/ffi_17/n5 ,
         \unit_fetch/unit_npcregister/ffi_16/n5 ,
         \unit_fetch/unit_npcregister/ffi_15/n5 ,
         \unit_fetch/unit_npcregister/ffi_14/n5 ,
         \unit_fetch/unit_npcregister/ffi_13/n5 ,
         \unit_fetch/unit_npcregister/ffi_12/n5 ,
         \unit_fetch/unit_npcregister/ffi_11/n5 ,
         \unit_fetch/unit_npcregister/ffi_10/n5 ,
         \unit_fetch/unit_npcregister/ffi_9/n5 ,
         \unit_fetch/unit_npcregister/ffi_8/n5 ,
         \unit_fetch/unit_npcregister/ffi_7/n5 ,
         \unit_fetch/unit_npcregister/ffi_6/n5 ,
         \unit_fetch/unit_npcregister/ffi_5/n5 ,
         \unit_fetch/unit_npcregister/ffi_4/n5 ,
         \unit_fetch/unit_npcregister/ffi_3/n5 ,
         \unit_fetch/unit_npcregister/ffi_2/n5 ,
         \unit_fetch/unit_npcregister/ffi_1/n5 ,
         \unit_fetch/unit_npcregister/ffi_0/n5 ,
         \unit_fetch/unit_programCounter/ffi_31/n5 ,
         \unit_fetch/unit_instructionRegister/n67 ,
         \unit_fetch/unit_instructionRegister/n68 ,
         \unit_fetch/unit_instructionRegister/n69 ,
         \unit_fetch/unit_instructionRegister/n71 ,
         \unit_fetch/unit_instructionRegister/n72 ,
         \unit_fetch/unit_instructionRegister/n73 ,
         \unit_fetch/unit_instructionRegister/n74 ,
         \unit_fetch/unit_instructionRegister/n75 ,
         \unit_fetch/unit_instructionRegister/n79 ,
         \unit_fetch/unit_instructionRegister/n80 ,
         \unit_fetch/unit_instructionRegister/n81 ,
         \unit_fetch/unit_instructionRegister/n83 ,
         \unit_fetch/unit_instructionRegister/n84 ,
         \unit_fetch/unit_instructionRegister/n85 ,
         \unit_fetch/unit_instructionRegister/n87 ,
         \unit_fetch/unit_instructionRegister/n88 ,
         \unit_fetch/unit_instructionRegister/n89 ,
         \unit_fetch/unit_instructionRegister/n90 ,
         \unit_fetch/unit_instructionRegister/n91 ,
         \unit_fetch/unit_instructionRegister/n92 ,
         \unit_fetch/unit_instructionRegister/n93 ,
         \unit_fetch/unit_instructionRegister/n95 ,
         \unit_fetch/unit_instructionRegister/n96 ,
         \unit_fetch/unit_instructionRegister/n97 ,
         \unit_fetch/unit_instructionRegister/n98 , \unit_fetch/pc_regout[2] ,
         \unit_fetch/pc_regout[3] , \unit_fetch/pc_regout[4] ,
         \unit_fetch/pc_regout[5] , \unit_fetch/pc_regout[6] ,
         \unit_fetch/pc_regout[7] , \unit_fetch/pc_regout[8] ,
         \unit_fetch/pc_regout[10] , \unit_fetch/pc_regout[11] ,
         \unit_fetch/pc_regout[12] , \unit_fetch/pc_regout[14] ,
         \unit_fetch/pc_regout[15] , \unit_fetch/pc_regout[16] ,
         \unit_fetch/pc_regout[18] , \unit_fetch/pc_regout[19] ,
         \unit_fetch/pc_regout[20] , \unit_fetch/pc_regout[21] ,
         \unit_fetch/pc_regout[22] , \unit_fetch/pc_regout[23] ,
         \unit_fetch/pc_regout[24] , \unit_fetch/pc_regout[26] ,
         \unit_fetch/pc_regout[27] , \unit_fetch/pc_regout[28] ,
         \unit_fetch/pc_regout[29] , \unit_fetch/pc_regout[30] ,
         \unit_fetch/pc_regout[31] , \unit_decode/n4138 , \unit_decode/n4137 ,
         \unit_decode/n4136 , \unit_decode/n4135 , \unit_decode/n4134 ,
         \unit_decode/n4133 , \unit_decode/n4132 , \unit_decode/n4131 ,
         \unit_decode/n4130 , \unit_decode/n4129 , \unit_decode/n4128 ,
         \unit_decode/n4127 , \unit_decode/n4126 , \unit_decode/n4125 ,
         \unit_decode/n4124 , \unit_decode/n4123 , \unit_decode/n4122 ,
         \unit_decode/n4121 , \unit_decode/n4120 , \unit_decode/n4119 ,
         \unit_decode/n4118 , \unit_decode/n4117 , \unit_decode/n4116 ,
         \unit_decode/n4115 , \unit_decode/n4114 , \unit_decode/n4113 ,
         \unit_decode/n4112 , \unit_decode/n4111 , \unit_decode/n4110 ,
         \unit_decode/n4109 , \unit_decode/n4108 , \unit_decode/n4107 ,
         \unit_decode/n4106 , \unit_decode/n4105 , \unit_decode/n4104 ,
         \unit_decode/n4103 , \unit_decode/n4102 , \unit_decode/n4101 ,
         \unit_decode/n4100 , \unit_decode/n4099 , \unit_decode/n4098 ,
         \unit_decode/n4097 , \unit_decode/n4096 , \unit_decode/n4095 ,
         \unit_decode/n4094 , \unit_decode/n4093 , \unit_decode/n4092 ,
         \unit_decode/n4091 , \unit_decode/n4090 , \unit_decode/n4089 ,
         \unit_decode/n4088 , \unit_decode/n4087 , \unit_decode/n4086 ,
         \unit_decode/n4085 , \unit_decode/n4084 , \unit_decode/n4083 ,
         \unit_decode/n4082 , \unit_decode/n4081 , \unit_decode/n4080 ,
         \unit_decode/n4079 , \unit_decode/n4078 , \unit_decode/n4077 ,
         \unit_decode/n4076 , \unit_decode/n4075 , \unit_decode/n4074 ,
         \unit_decode/n4073 , \unit_decode/n4072 , \unit_decode/n4071 ,
         \unit_decode/n4070 , \unit_decode/n4069 , \unit_decode/n4068 ,
         \unit_decode/n4067 , \unit_decode/n4066 , \unit_decode/n4065 ,
         \unit_decode/n4064 , \unit_decode/n4063 , \unit_decode/n4062 ,
         \unit_decode/n4061 , \unit_decode/n4060 , \unit_decode/n4059 ,
         \unit_decode/n4058 , \unit_decode/n4057 , \unit_decode/n4056 ,
         \unit_decode/n4055 , \unit_decode/n4054 , \unit_decode/n4053 ,
         \unit_decode/n4052 , \unit_decode/n4051 , \unit_decode/n4050 ,
         \unit_decode/n4049 , \unit_decode/n4048 , \unit_decode/n4047 ,
         \unit_decode/n4046 , \unit_decode/n4045 , \unit_decode/n4044 ,
         \unit_decode/n4043 , \unit_decode/n4042 , \unit_decode/n4041 ,
         \unit_decode/n4040 , \unit_decode/n4039 , \unit_decode/n4038 ,
         \unit_decode/n4037 , \unit_decode/n4036 , \unit_decode/n4035 ,
         \unit_decode/n4034 , \unit_decode/n4033 , \unit_decode/n4032 ,
         \unit_decode/n4031 , \unit_decode/n4030 , \unit_decode/n4029 ,
         \unit_decode/n4028 , \unit_decode/n4027 , \unit_decode/n4026 ,
         \unit_decode/n4025 , \unit_decode/n4024 , \unit_decode/n4023 ,
         \unit_decode/n4022 , \unit_decode/n4021 , \unit_decode/n4020 ,
         \unit_decode/n4019 , \unit_decode/n4018 , \unit_decode/n4017 ,
         \unit_decode/n4016 , \unit_decode/n4015 , \unit_decode/n4014 ,
         \unit_decode/n4013 , \unit_decode/n4012 , \unit_decode/n4011 ,
         \unit_decode/n4006 , \unit_decode/n4005 , \unit_decode/n4000 ,
         \unit_decode/n3999 , \unit_decode/n3994 , \unit_decode/n3993 ,
         \unit_decode/n3988 , \unit_decode/n3987 , \unit_decode/n3982 ,
         \unit_decode/n3981 , \unit_decode/n3976 , \unit_decode/n3975 ,
         \unit_decode/n3970 , \unit_decode/n3969 , \unit_decode/n3964 ,
         \unit_decode/n3963 , \unit_decode/n3958 , \unit_decode/n3957 ,
         \unit_decode/n3952 , \unit_decode/n3951 , \unit_decode/n3946 ,
         \unit_decode/n3945 , \unit_decode/n3940 , \unit_decode/n3939 ,
         \unit_decode/n3934 , \unit_decode/n3933 , \unit_decode/n3928 ,
         \unit_decode/n3927 , \unit_decode/n3922 , \unit_decode/n3921 ,
         \unit_decode/n3916 , \unit_decode/n3915 , \unit_decode/n3910 ,
         \unit_decode/n3909 , \unit_decode/n3904 , \unit_decode/n3903 ,
         \unit_decode/n3898 , \unit_decode/n3897 , \unit_decode/n3892 ,
         \unit_decode/n3891 , \unit_decode/n3886 , \unit_decode/n3885 ,
         \unit_decode/n3880 , \unit_decode/n3879 , \unit_decode/n3874 ,
         \unit_decode/n3873 , \unit_decode/n3868 , \unit_decode/n3867 ,
         \unit_decode/n3862 , \unit_decode/n3861 , \unit_decode/n3856 ,
         \unit_decode/n3855 , \unit_decode/n3850 , \unit_decode/n3849 ,
         \unit_decode/n3844 , \unit_decode/n3843 , \unit_decode/n3838 ,
         \unit_decode/n3837 , \unit_decode/n3832 , \unit_decode/n3831 ,
         \unit_decode/n3826 , \unit_decode/n3825 , \unit_decode/n3820 ,
         \unit_decode/n3819 , \unit_decode/n3814 , \unit_decode/n3813 ,
         \unit_decode/n3808 , \unit_decode/n3807 , \unit_decode/n3802 ,
         \unit_decode/n3801 , \unit_decode/n3796 , \unit_decode/n3795 ,
         \unit_decode/n3790 , \unit_decode/n3789 , \unit_decode/n3784 ,
         \unit_decode/n3783 , \unit_decode/n3778 , \unit_decode/n3777 ,
         \unit_decode/n3772 , \unit_decode/n3771 , \unit_decode/n3766 ,
         \unit_decode/n3765 , \unit_decode/n3760 , \unit_decode/n3759 ,
         \unit_decode/n3754 , \unit_decode/n3753 , \unit_decode/n3748 ,
         \unit_decode/n3747 , \unit_decode/n3742 , \unit_decode/n3741 ,
         \unit_decode/n3736 , \unit_decode/n3735 , \unit_decode/n3730 ,
         \unit_decode/n3729 , \unit_decode/n3724 , \unit_decode/n3723 ,
         \unit_decode/n3718 , \unit_decode/n3717 , \unit_decode/n3712 ,
         \unit_decode/n3711 , \unit_decode/n3706 , \unit_decode/n3705 ,
         \unit_decode/n3700 , \unit_decode/n3699 , \unit_decode/n3694 ,
         \unit_decode/n3693 , \unit_decode/n3688 , \unit_decode/n3687 ,
         \unit_decode/n3682 , \unit_decode/n3681 , \unit_decode/n3676 ,
         \unit_decode/n3675 , \unit_decode/n3670 , \unit_decode/n3669 ,
         \unit_decode/n3664 , \unit_decode/n3663 , \unit_decode/n3658 ,
         \unit_decode/n3657 , \unit_decode/n3652 , \unit_decode/n3651 ,
         \unit_decode/n3646 , \unit_decode/n3645 , \unit_decode/n3640 ,
         \unit_decode/n3639 , \unit_decode/n3634 , \unit_decode/n3633 ,
         \unit_decode/n3628 , \unit_decode/n3627 , \unit_decode/n3626 ,
         \unit_decode/n3625 , \unit_decode/n3624 , \unit_decode/n3623 ,
         \unit_decode/n3622 , \unit_decode/n3621 , \unit_decode/n3620 ,
         \unit_decode/n3619 , \unit_decode/n3618 , \unit_decode/n3617 ,
         \unit_decode/n3616 , \unit_decode/n3615 , \unit_decode/n3614 ,
         \unit_decode/n3613 , \unit_decode/n3612 , \unit_decode/n3611 ,
         \unit_decode/n3610 , \unit_decode/n3609 , \unit_decode/n3608 ,
         \unit_decode/n3607 , \unit_decode/n3606 , \unit_decode/n3605 ,
         \unit_decode/n3604 , \unit_decode/n3603 , \unit_decode/n3602 ,
         \unit_decode/n3601 , \unit_decode/n3600 , \unit_decode/n3599 ,
         \unit_decode/n3598 , \unit_decode/n3597 , \unit_decode/n3596 ,
         \unit_decode/n3595 , \unit_decode/n3594 , \unit_decode/n3593 ,
         \unit_decode/n3592 , \unit_decode/n3591 , \unit_decode/n3590 ,
         \unit_decode/n3589 , \unit_decode/n3588 , \unit_decode/n3587 ,
         \unit_decode/n3586 , \unit_decode/n3585 , \unit_decode/n3584 ,
         \unit_decode/n3583 , \unit_decode/n3582 , \unit_decode/n3581 ,
         \unit_decode/n3580 , \unit_decode/n3579 , \unit_decode/n3578 ,
         \unit_decode/n3577 , \unit_decode/n3576 , \unit_decode/n3575 ,
         \unit_decode/n3574 , \unit_decode/n3573 , \unit_decode/n3572 ,
         \unit_decode/n3571 , \unit_decode/n3570 , \unit_decode/n3569 ,
         \unit_decode/n3568 , \unit_decode/n3567 , \unit_decode/n3566 ,
         \unit_decode/n3565 , \unit_decode/n3564 , \unit_decode/n3563 ,
         \unit_decode/n3562 , \unit_decode/n3561 , \unit_decode/n3560 ,
         \unit_decode/n3559 , \unit_decode/n3558 , \unit_decode/n3557 ,
         \unit_decode/n3556 , \unit_decode/n3555 , \unit_decode/n3554 ,
         \unit_decode/n3553 , \unit_decode/n3552 , \unit_decode/n3551 ,
         \unit_decode/n3550 , \unit_decode/n3549 , \unit_decode/n3548 ,
         \unit_decode/n3547 , \unit_decode/n3546 , \unit_decode/n3545 ,
         \unit_decode/n3544 , \unit_decode/n3543 , \unit_decode/n3542 ,
         \unit_decode/n3541 , \unit_decode/n3540 , \unit_decode/n3539 ,
         \unit_decode/n3538 , \unit_decode/n3537 , \unit_decode/n3536 ,
         \unit_decode/n3535 , \unit_decode/n3534 , \unit_decode/n3533 ,
         \unit_decode/n3532 , \unit_decode/n3531 , \unit_decode/n3530 ,
         \unit_decode/n3529 , \unit_decode/n3528 , \unit_decode/n3527 ,
         \unit_decode/n3526 , \unit_decode/n3525 , \unit_decode/n3524 ,
         \unit_decode/n3523 , \unit_decode/n3522 , \unit_decode/n3521 ,
         \unit_decode/n3520 , \unit_decode/n3519 , \unit_decode/n3517 ,
         \unit_decode/n3516 , \unit_decode/n3515 , \unit_decode/n3514 ,
         \unit_decode/n3513 , \unit_decode/n3512 , \unit_decode/n3511 ,
         \unit_decode/n3510 , \unit_decode/n3509 , \unit_decode/n3508 ,
         \unit_decode/n3507 , \unit_decode/n3506 , \unit_decode/n3505 ,
         \unit_decode/n3504 , \unit_decode/n3503 , \unit_decode/n3502 ,
         \unit_decode/n3501 , \unit_decode/n3500 , \unit_decode/n3499 ,
         \unit_decode/n3498 , \unit_decode/n3497 , \unit_decode/n3496 ,
         \unit_decode/n3495 , \unit_decode/n3494 , \unit_decode/n3493 ,
         \unit_decode/n3492 , \unit_decode/n3491 , \unit_decode/n3490 ,
         \unit_decode/n3489 , \unit_decode/n3488 , \unit_decode/n3487 ,
         \unit_decode/n3486 , \unit_decode/n3485 , \unit_decode/n3484 ,
         \unit_decode/n3483 , \unit_decode/n3482 , \unit_decode/n3481 ,
         \unit_decode/n3480 , \unit_decode/n3479 , \unit_decode/n3478 ,
         \unit_decode/n3477 , \unit_decode/n3476 , \unit_decode/n3475 ,
         \unit_decode/n3474 , \unit_decode/n3473 , \unit_decode/n3472 ,
         \unit_decode/n3471 , \unit_decode/n3470 , \unit_decode/n3469 ,
         \unit_decode/n3468 , \unit_decode/n3467 , \unit_decode/n3466 ,
         \unit_decode/n3465 , \unit_decode/n3464 , \unit_decode/n3463 ,
         \unit_decode/n3462 , \unit_decode/n3461 , \unit_decode/n3460 ,
         \unit_decode/n3459 , \unit_decode/n3458 , \unit_decode/n3457 ,
         \unit_decode/n3456 , \unit_decode/n3455 , \unit_decode/n3454 ,
         \unit_decode/n3453 , \unit_decode/n3452 , \unit_decode/n3451 ,
         \unit_decode/n3450 , \unit_decode/n3449 , \unit_decode/n3448 ,
         \unit_decode/n3447 , \unit_decode/n3446 , \unit_decode/n3445 ,
         \unit_decode/n3444 , \unit_decode/n3443 , \unit_decode/n3442 ,
         \unit_decode/n3441 , \unit_decode/n3440 , \unit_decode/n3439 ,
         \unit_decode/n3438 , \unit_decode/n3437 , \unit_decode/n3436 ,
         \unit_decode/n3435 , \unit_decode/n3434 , \unit_decode/n3433 ,
         \unit_decode/n3432 , \unit_decode/n3431 , \unit_decode/n3430 ,
         \unit_decode/n3429 , \unit_decode/n3428 , \unit_decode/n3427 ,
         \unit_decode/n3426 , \unit_decode/n3425 , \unit_decode/n3424 ,
         \unit_decode/n3423 , \unit_decode/n3422 , \unit_decode/n3421 ,
         \unit_decode/n3420 , \unit_decode/n3419 , \unit_decode/n3418 ,
         \unit_decode/n3417 , \unit_decode/n3416 , \unit_decode/n3415 ,
         \unit_decode/n3414 , \unit_decode/n3413 , \unit_decode/n3412 ,
         \unit_decode/n3411 , \unit_decode/n3410 , \unit_decode/n3409 ,
         \unit_decode/n3408 , \unit_decode/n3407 , \unit_decode/n3406 ,
         \unit_decode/n3405 , \unit_decode/n3404 , \unit_decode/n3403 ,
         \unit_decode/n3402 , \unit_decode/n3401 , \unit_decode/n3400 ,
         \unit_decode/n3399 , \unit_decode/n3398 , \unit_decode/n3397 ,
         \unit_decode/n3396 , \unit_decode/n3395 , \unit_decode/n3394 ,
         \unit_decode/n3393 , \unit_decode/n3392 , \unit_decode/n3391 ,
         \unit_decode/n3390 , \unit_decode/n3389 , \unit_decode/n3388 ,
         \unit_decode/n3387 , \unit_decode/n3386 , \unit_decode/n3385 ,
         \unit_decode/n3384 , \unit_decode/n3383 , \unit_decode/n3382 ,
         \unit_decode/n3381 , \unit_decode/n3380 , \unit_decode/n3379 ,
         \unit_decode/n3378 , \unit_decode/n3377 , \unit_decode/n3376 ,
         \unit_decode/n3375 , \unit_decode/n3374 , \unit_decode/n3373 ,
         \unit_decode/n3372 , \unit_decode/n3371 , \unit_decode/n3370 ,
         \unit_decode/n3369 , \unit_decode/n3368 , \unit_decode/n3367 ,
         \unit_decode/n3366 , \unit_decode/n3365 , \unit_decode/n3364 ,
         \unit_decode/n3363 , \unit_decode/n3362 , \unit_decode/n3361 ,
         \unit_decode/n3360 , \unit_decode/n3359 , \unit_decode/n3358 ,
         \unit_decode/n3357 , \unit_decode/n3356 , \unit_decode/n3355 ,
         \unit_decode/n3354 , \unit_decode/n3353 , \unit_decode/n3352 ,
         \unit_decode/n3351 , \unit_decode/n3350 , \unit_decode/n3349 ,
         \unit_decode/n3348 , \unit_decode/n3347 , \unit_decode/n3346 ,
         \unit_decode/n3345 , \unit_decode/n3344 , \unit_decode/n3343 ,
         \unit_decode/n3342 , \unit_decode/n3341 , \unit_decode/n3340 ,
         \unit_decode/n3339 , \unit_decode/n3338 , \unit_decode/n3337 ,
         \unit_decode/n3336 , \unit_decode/n3335 , \unit_decode/n3334 ,
         \unit_decode/n3333 , \unit_decode/n3332 , \unit_decode/n3331 ,
         \unit_decode/n3330 , \unit_decode/n3329 , \unit_decode/n3328 ,
         \unit_decode/n3327 , \unit_decode/n3326 , \unit_decode/n3325 ,
         \unit_decode/n3324 , \unit_decode/n3323 , \unit_decode/n3322 ,
         \unit_decode/n3321 , \unit_decode/n3320 , \unit_decode/n3319 ,
         \unit_decode/n3318 , \unit_decode/n3317 , \unit_decode/n3316 ,
         \unit_decode/n3315 , \unit_decode/n3314 , \unit_decode/n3313 ,
         \unit_decode/n3312 , \unit_decode/n3311 , \unit_decode/n3310 ,
         \unit_decode/n3309 , \unit_decode/n3308 , \unit_decode/n3307 ,
         \unit_decode/n3306 , \unit_decode/n3305 , \unit_decode/n3304 ,
         \unit_decode/n3303 , \unit_decode/n3302 , \unit_decode/n3301 ,
         \unit_decode/n3300 , \unit_decode/n3299 , \unit_decode/n3298 ,
         \unit_decode/n3297 , \unit_decode/n3296 , \unit_decode/n3295 ,
         \unit_decode/n3294 , \unit_decode/n3293 , \unit_decode/n3292 ,
         \unit_decode/n3291 , \unit_decode/n3290 , \unit_decode/n3289 ,
         \unit_decode/n3288 , \unit_decode/n3287 , \unit_decode/n3286 ,
         \unit_decode/n3285 , \unit_decode/n3284 , \unit_decode/n3283 ,
         \unit_decode/n3282 , \unit_decode/n3281 , \unit_decode/n3280 ,
         \unit_decode/n3279 , \unit_decode/n3278 , \unit_decode/n3277 ,
         \unit_decode/n3276 , \unit_decode/n3275 , \unit_decode/n3274 ,
         \unit_decode/n3273 , \unit_decode/n3272 , \unit_decode/n3271 ,
         \unit_decode/n3270 , \unit_decode/n3269 , \unit_decode/n3268 ,
         \unit_decode/n3267 , \unit_decode/n3266 , \unit_decode/n3265 ,
         \unit_decode/n3264 , \unit_decode/n3263 , \unit_decode/n3262 ,
         \unit_decode/n3261 , \unit_decode/n3260 , \unit_decode/n3259 ,
         \unit_decode/n3258 , \unit_decode/n3257 , \unit_decode/n3256 ,
         \unit_decode/n3255 , \unit_decode/n3254 , \unit_decode/n3253 ,
         \unit_decode/n3252 , \unit_decode/n3251 , \unit_decode/n3250 ,
         \unit_decode/n3249 , \unit_decode/n3248 , \unit_decode/n3247 ,
         \unit_decode/n3246 , \unit_decode/n3245 , \unit_decode/n3244 ,
         \unit_decode/n3243 , \unit_decode/n3242 , \unit_decode/n3241 ,
         \unit_decode/n3240 , \unit_decode/n3239 , \unit_decode/n3238 ,
         \unit_decode/n3237 , \unit_decode/n3236 , \unit_decode/n3235 ,
         \unit_decode/n3234 , \unit_decode/n3233 , \unit_decode/n3232 ,
         \unit_decode/n3231 , \unit_decode/n3230 , \unit_decode/n3229 ,
         \unit_decode/n3228 , \unit_decode/n3227 , \unit_decode/n3226 ,
         \unit_decode/n3225 , \unit_decode/n3224 , \unit_decode/n3223 ,
         \unit_decode/n3222 , \unit_decode/n3221 , \unit_decode/n3220 ,
         \unit_decode/n3219 , \unit_decode/n3218 , \unit_decode/n3217 ,
         \unit_decode/n3216 , \unit_decode/n3215 , \unit_decode/n3214 ,
         \unit_decode/n3213 , \unit_decode/n3212 , \unit_decode/n3211 ,
         \unit_decode/n3210 , \unit_decode/n3209 , \unit_decode/n3208 ,
         \unit_decode/n3207 , \unit_decode/n3206 , \unit_decode/n3205 ,
         \unit_decode/n3204 , \unit_decode/n3203 , \unit_decode/n3202 ,
         \unit_decode/n3201 , \unit_decode/n3200 , \unit_decode/n3199 ,
         \unit_decode/n3198 , \unit_decode/n3197 , \unit_decode/n3196 ,
         \unit_decode/n3195 , \unit_decode/n3194 , \unit_decode/n3193 ,
         \unit_decode/n3192 , \unit_decode/n3191 , \unit_decode/n3190 ,
         \unit_decode/n3189 , \unit_decode/n3188 , \unit_decode/n3187 ,
         \unit_decode/n3186 , \unit_decode/n3185 , \unit_decode/n3184 ,
         \unit_decode/n3183 , \unit_decode/n3182 , \unit_decode/n3181 ,
         \unit_decode/n3180 , \unit_decode/n3179 , \unit_decode/n3178 ,
         \unit_decode/n3177 , \unit_decode/n3176 , \unit_decode/n3175 ,
         \unit_decode/n3174 , \unit_decode/n3173 , \unit_decode/n3172 ,
         \unit_decode/n3171 , \unit_decode/n3170 , \unit_decode/n3169 ,
         \unit_decode/n3168 , \unit_decode/n3167 , \unit_decode/n3166 ,
         \unit_decode/n3165 , \unit_decode/n3164 , \unit_decode/n3163 ,
         \unit_decode/n3162 , \unit_decode/n3161 , \unit_decode/n3160 ,
         \unit_decode/n3159 , \unit_decode/n3158 , \unit_decode/n3157 ,
         \unit_decode/n3156 , \unit_decode/n3155 , \unit_decode/n3154 ,
         \unit_decode/n3153 , \unit_decode/n3152 , \unit_decode/n3151 ,
         \unit_decode/n3150 , \unit_decode/n3149 , \unit_decode/n3148 ,
         \unit_decode/n3147 , \unit_decode/n3146 , \unit_decode/n3145 ,
         \unit_decode/n3144 , \unit_decode/n3143 , \unit_decode/n3142 ,
         \unit_decode/n3141 , \unit_decode/n3140 , \unit_decode/n3139 ,
         \unit_decode/n3138 , \unit_decode/n3137 , \unit_decode/n3136 ,
         \unit_decode/n3135 , \unit_decode/n3134 , \unit_decode/n3133 ,
         \unit_decode/n3132 , \unit_decode/n3131 , \unit_decode/n3130 ,
         \unit_decode/n3129 , \unit_decode/n3128 , \unit_decode/n3127 ,
         \unit_decode/n3126 , \unit_decode/n3125 , \unit_decode/n3124 ,
         \unit_decode/n3123 , \unit_decode/n3122 , \unit_decode/n3121 ,
         \unit_decode/n3120 , \unit_decode/n3119 , \unit_decode/n3118 ,
         \unit_decode/n3117 , \unit_decode/n3116 , \unit_decode/n3115 ,
         \unit_decode/n3114 , \unit_decode/n3113 , \unit_decode/n3112 ,
         \unit_decode/n3111 , \unit_decode/n3110 , \unit_decode/n3109 ,
         \unit_decode/n3108 , \unit_decode/n3107 , \unit_decode/n3106 ,
         \unit_decode/n3105 , \unit_decode/n3104 , \unit_decode/n3103 ,
         \unit_decode/n3102 , \unit_decode/n3101 , \unit_decode/n3100 ,
         \unit_decode/n3099 , \unit_decode/n3098 , \unit_decode/n3097 ,
         \unit_decode/n3096 , \unit_decode/n3095 , \unit_decode/n3094 ,
         \unit_decode/n3093 , \unit_decode/n3092 , \unit_decode/n3091 ,
         \unit_decode/n3090 , \unit_decode/n3089 , \unit_decode/n3088 ,
         \unit_decode/n3087 , \unit_decode/n3086 , \unit_decode/n3085 ,
         \unit_decode/n3084 , \unit_decode/n3083 , \unit_decode/n3082 ,
         \unit_decode/n3081 , \unit_decode/n3080 , \unit_decode/n3079 ,
         \unit_decode/n3078 , \unit_decode/n3077 , \unit_decode/n3076 ,
         \unit_decode/n3075 , \unit_decode/n3074 , \unit_decode/n3073 ,
         \unit_decode/n3072 , \unit_decode/n3071 , \unit_decode/n3070 ,
         \unit_decode/n3069 , \unit_decode/n3068 , \unit_decode/n3067 ,
         \unit_decode/n3066 , \unit_decode/n3065 , \unit_decode/n3064 ,
         \unit_decode/n3063 , \unit_decode/n3062 , \unit_decode/n3061 ,
         \unit_decode/n3060 , \unit_decode/n3059 , \unit_decode/n3058 ,
         \unit_decode/n3057 , \unit_decode/n3056 , \unit_decode/n3055 ,
         \unit_decode/n3054 , \unit_decode/n3053 , \unit_decode/n3052 ,
         \unit_decode/n3051 , \unit_decode/n3050 , \unit_decode/n3049 ,
         \unit_decode/n3048 , \unit_decode/n3047 , \unit_decode/n3046 ,
         \unit_decode/n3045 , \unit_decode/n3044 , \unit_decode/n3043 ,
         \unit_decode/n3042 , \unit_decode/n3041 , \unit_decode/n3040 ,
         \unit_decode/n3039 , \unit_decode/n3038 , \unit_decode/n3037 ,
         \unit_decode/n3036 , \unit_decode/n3035 , \unit_decode/n3034 ,
         \unit_decode/n3033 , \unit_decode/n3032 , \unit_decode/n3031 ,
         \unit_decode/n3030 , \unit_decode/n3029 , \unit_decode/n3028 ,
         \unit_decode/n3027 , \unit_decode/n3026 , \unit_decode/n3025 ,
         \unit_decode/n3024 , \unit_decode/n3023 , \unit_decode/n3022 ,
         \unit_decode/n3021 , \unit_decode/n3020 , \unit_decode/n3019 ,
         \unit_decode/n3018 , \unit_decode/n3017 , \unit_decode/n3016 ,
         \unit_decode/n3015 , \unit_decode/n3014 , \unit_decode/n3013 ,
         \unit_decode/n3012 , \unit_decode/n3011 , \unit_decode/n3010 ,
         \unit_decode/n3009 , \unit_decode/n3008 , \unit_decode/n3007 ,
         \unit_decode/n3006 , \unit_decode/n3005 , \unit_decode/n3004 ,
         \unit_decode/n3003 , \unit_decode/n3002 , \unit_decode/n3001 ,
         \unit_decode/n3000 , \unit_decode/n2999 , \unit_decode/n2998 ,
         \unit_decode/n2997 , \unit_decode/n2996 , \unit_decode/n2995 ,
         \unit_decode/n2994 , \unit_decode/n2993 , \unit_decode/n2992 ,
         \unit_decode/n2991 , \unit_decode/n2990 , \unit_decode/n2989 ,
         \unit_decode/n2988 , \unit_decode/n2987 , \unit_decode/n2986 ,
         \unit_decode/n2985 , \unit_decode/n2984 , \unit_decode/n2983 ,
         \unit_decode/n2982 , \unit_decode/n2981 , \unit_decode/n2980 ,
         \unit_decode/n2979 , \unit_decode/n2978 , \unit_decode/n2977 ,
         \unit_decode/n2976 , \unit_decode/n2975 , \unit_decode/n2974 ,
         \unit_decode/n2973 , \unit_decode/n2972 , \unit_decode/n2971 ,
         \unit_decode/n2970 , \unit_decode/n2969 , \unit_decode/n2968 ,
         \unit_decode/n2967 , \unit_decode/n2966 , \unit_decode/n2965 ,
         \unit_decode/n2964 , \unit_decode/n2963 , \unit_decode/n2962 ,
         \unit_decode/n2961 , \unit_decode/n2960 , \unit_decode/n2959 ,
         \unit_decode/n2958 , \unit_decode/n2957 , \unit_decode/n2956 ,
         \unit_decode/n2955 , \unit_decode/n2954 , \unit_decode/n2953 ,
         \unit_decode/n2952 , \unit_decode/n2951 , \unit_decode/n2950 ,
         \unit_decode/n2949 , \unit_decode/n2948 , \unit_decode/n2947 ,
         \unit_decode/n2946 , \unit_decode/n2945 , \unit_decode/n2944 ,
         \unit_decode/n2943 , \unit_decode/n2942 , \unit_decode/n2941 ,
         \unit_decode/n2940 , \unit_decode/n2939 , \unit_decode/n2938 ,
         \unit_decode/n2937 , \unit_decode/n2936 , \unit_decode/n2935 ,
         \unit_decode/n2934 , \unit_decode/n2933 , \unit_decode/n2932 ,
         \unit_decode/n2931 , \unit_decode/n2930 , \unit_decode/n2929 ,
         \unit_decode/n2928 , \unit_decode/n2927 , \unit_decode/n2926 ,
         \unit_decode/n2925 , \unit_decode/n2924 , \unit_decode/n2923 ,
         \unit_decode/n2922 , \unit_decode/n2921 , \unit_decode/n2920 ,
         \unit_decode/n2919 , \unit_decode/n2918 , \unit_decode/n2917 ,
         \unit_decode/n2916 , \unit_decode/n2915 , \unit_decode/n2914 ,
         \unit_decode/n2913 , \unit_decode/n2912 , \unit_decode/n2911 ,
         \unit_decode/n2910 , \unit_decode/n2909 , \unit_decode/n2908 ,
         \unit_decode/n2907 , \unit_decode/n2906 , \unit_decode/n2905 ,
         \unit_decode/n2904 , \unit_decode/n2903 , \unit_decode/n2902 ,
         \unit_decode/n2901 , \unit_decode/n2900 , \unit_decode/n2899 ,
         \unit_decode/n2898 , \unit_decode/n2897 , \unit_decode/n2896 ,
         \unit_decode/n2895 , \unit_decode/n2894 , \unit_decode/n2893 ,
         \unit_decode/n2892 , \unit_decode/n2891 , \unit_decode/n2890 ,
         \unit_decode/n2889 , \unit_decode/n2888 , \unit_decode/n2887 ,
         \unit_decode/n2886 , \unit_decode/n2885 , \unit_decode/n2884 ,
         \unit_decode/n2883 , \unit_decode/n2882 , \unit_decode/n2881 ,
         \unit_decode/n2880 , \unit_decode/n2879 , \unit_decode/n2878 ,
         \unit_decode/n2877 , \unit_decode/n2876 , \unit_decode/n2875 ,
         \unit_decode/n2874 , \unit_decode/n2873 , \unit_decode/n2872 ,
         \unit_decode/n2871 , \unit_decode/n2870 , \unit_decode/n2869 ,
         \unit_decode/n2868 , \unit_decode/n2867 , \unit_decode/n2866 ,
         \unit_decode/n2865 , \unit_decode/n2864 , \unit_decode/n2863 ,
         \unit_decode/n2862 , \unit_decode/n2861 , \unit_decode/n2860 ,
         \unit_decode/n2859 , \unit_decode/n2858 , \unit_decode/n2857 ,
         \unit_decode/n2856 , \unit_decode/n2855 , \unit_decode/n2854 ,
         \unit_decode/n2853 , \unit_decode/n2852 , \unit_decode/n2851 ,
         \unit_decode/n2850 , \unit_decode/n2849 , \unit_decode/n2848 ,
         \unit_decode/n2847 , \unit_decode/n2846 , \unit_decode/n2845 ,
         \unit_decode/n2844 , \unit_decode/n2843 , \unit_decode/n2842 ,
         \unit_decode/n2841 , \unit_decode/n2840 , \unit_decode/n2839 ,
         \unit_decode/n2838 , \unit_decode/n2837 , \unit_decode/n2836 ,
         \unit_decode/n2835 , \unit_decode/n2834 , \unit_decode/n2833 ,
         \unit_decode/n2832 , \unit_decode/n2831 , \unit_decode/n2830 ,
         \unit_decode/n2829 , \unit_decode/n2828 , \unit_decode/n2827 ,
         \unit_decode/n2826 , \unit_decode/n2825 , \unit_decode/n2824 ,
         \unit_decode/n2823 , \unit_decode/n2822 , \unit_decode/n2821 ,
         \unit_decode/n2820 , \unit_decode/n2819 , \unit_decode/n2818 ,
         \unit_decode/n2817 , \unit_decode/n2816 , \unit_decode/n2815 ,
         \unit_decode/n2814 , \unit_decode/n2813 , \unit_decode/n2812 ,
         \unit_decode/n2811 , \unit_decode/n2810 , \unit_decode/n2809 ,
         \unit_decode/n2808 , \unit_decode/n2807 , \unit_decode/n2806 ,
         \unit_decode/n2805 , \unit_decode/n2804 , \unit_decode/n2803 ,
         \unit_decode/n2802 , \unit_decode/n2801 , \unit_decode/n2800 ,
         \unit_decode/n2799 , \unit_decode/n2798 , \unit_decode/n2797 ,
         \unit_decode/n2796 , \unit_decode/n2795 , \unit_decode/n2794 ,
         \unit_decode/n2793 , \unit_decode/n2792 , \unit_decode/n2791 ,
         \unit_decode/n2790 , \unit_decode/n2789 , \unit_decode/n2788 ,
         \unit_decode/n2787 , \unit_decode/n2786 , \unit_decode/n2785 ,
         \unit_decode/n2784 , \unit_decode/n2783 , \unit_decode/n2782 ,
         \unit_decode/n2781 , \unit_decode/n2780 , \unit_decode/n2779 ,
         \unit_decode/n2778 , \unit_decode/n2777 , \unit_decode/n2776 ,
         \unit_decode/n2775 , \unit_decode/n2774 , \unit_decode/n2773 ,
         \unit_decode/n2772 , \unit_decode/n2771 , \unit_decode/n2770 ,
         \unit_decode/n2769 , \unit_decode/n2768 , \unit_decode/n2767 ,
         \unit_decode/n2766 , \unit_decode/n2765 , \unit_decode/n2764 ,
         \unit_decode/n2763 , \unit_decode/n2762 , \unit_decode/n2761 ,
         \unit_decode/n2760 , \unit_decode/n2759 , \unit_decode/n2758 ,
         \unit_decode/n2757 , \unit_decode/n2756 , \unit_decode/n2755 ,
         \unit_decode/n2754 , \unit_decode/n2753 , \unit_decode/n2752 ,
         \unit_decode/n2751 , \unit_decode/n2750 , \unit_decode/n2749 ,
         \unit_decode/n2748 , \unit_decode/n2747 , \unit_decode/n2746 ,
         \unit_decode/n2745 , \unit_decode/n2744 , \unit_decode/n2743 ,
         \unit_decode/n2742 , \unit_decode/n2741 , \unit_decode/n2740 ,
         \unit_decode/n2739 , \unit_decode/n2738 , \unit_decode/n2737 ,
         \unit_decode/n2736 , \unit_decode/n2735 , \unit_decode/n2734 ,
         \unit_decode/n2733 , \unit_decode/n2732 , \unit_decode/n2731 ,
         \unit_decode/n2730 , \unit_decode/n2729 , \unit_decode/n2728 ,
         \unit_decode/n2727 , \unit_decode/n2726 , \unit_decode/n2725 ,
         \unit_decode/n2724 , \unit_decode/n2723 , \unit_decode/n2722 ,
         \unit_decode/n2721 , \unit_decode/n2720 , \unit_decode/n2719 ,
         \unit_decode/n2718 , \unit_decode/n2717 , \unit_decode/n2716 ,
         \unit_decode/n2715 , \unit_decode/n2714 , \unit_decode/n2713 ,
         \unit_decode/n2712 , \unit_decode/n2711 , \unit_decode/n2710 ,
         \unit_decode/n2709 , \unit_decode/n2708 , \unit_decode/n2707 ,
         \unit_decode/n2706 , \unit_decode/n2705 , \unit_decode/n2704 ,
         \unit_decode/n2703 , \unit_decode/n2702 , \unit_decode/n2701 ,
         \unit_decode/n2700 , \unit_decode/n2699 , \unit_decode/n2698 ,
         \unit_decode/n2697 , \unit_decode/n2696 , \unit_decode/n2695 ,
         \unit_decode/n2694 , \unit_decode/n2693 , \unit_decode/n2692 ,
         \unit_decode/n2691 , \unit_decode/n2690 , \unit_decode/n2689 ,
         \unit_decode/n2688 , \unit_decode/n2687 , \unit_decode/n2686 ,
         \unit_decode/n2685 , \unit_decode/n2684 , \unit_decode/n2683 ,
         \unit_decode/n2682 , \unit_decode/n2681 , \unit_decode/n2680 ,
         \unit_decode/n2679 , \unit_decode/n2678 , \unit_decode/n2677 ,
         \unit_decode/n2676 , \unit_decode/n2675 , \unit_decode/n2674 ,
         \unit_decode/n2673 , \unit_decode/n2672 , \unit_decode/n2671 ,
         \unit_decode/n2670 , \unit_decode/n2669 , \unit_decode/n2668 ,
         \unit_decode/n2667 , \unit_decode/n2666 , \unit_decode/n2665 ,
         \unit_decode/n2664 , \unit_decode/n2663 , \unit_decode/n2662 ,
         \unit_decode/n2661 , \unit_decode/n2660 , \unit_decode/n2659 ,
         \unit_decode/n2658 , \unit_decode/n2657 , \unit_decode/n2656 ,
         \unit_decode/n2655 , \unit_decode/n2654 , \unit_decode/n2653 ,
         \unit_decode/n2652 , \unit_decode/n2651 , \unit_decode/n2650 ,
         \unit_decode/n2649 , \unit_decode/n2648 , \unit_decode/n2647 ,
         \unit_decode/n2646 , \unit_decode/n2645 , \unit_decode/n2644 ,
         \unit_decode/n2643 , \unit_decode/n2642 , \unit_decode/n2641 ,
         \unit_decode/n2640 , \unit_decode/n2639 , \unit_decode/n2638 ,
         \unit_decode/n2637 , \unit_decode/n2636 , \unit_decode/n2635 ,
         \unit_decode/n2634 , \unit_decode/n2633 , \unit_decode/n2632 ,
         \unit_decode/n2631 , \unit_decode/n2630 , \unit_decode/n2629 ,
         \unit_decode/n2628 , \unit_decode/n2627 , \unit_decode/n2626 ,
         \unit_decode/n2625 , \unit_decode/n2624 , \unit_decode/n2623 ,
         \unit_decode/n2622 , \unit_decode/n2621 , \unit_decode/n2620 ,
         \unit_decode/n2619 , \unit_decode/n2618 , \unit_decode/n2617 ,
         \unit_decode/n2616 , \unit_decode/n2615 , \unit_decode/n2614 ,
         \unit_decode/n2613 , \unit_decode/n2612 , \unit_decode/n2611 ,
         \unit_decode/n2610 , \unit_decode/n2609 , \unit_decode/n2608 ,
         \unit_decode/n2607 , \unit_decode/n2606 , \unit_decode/n2605 ,
         \unit_decode/n2604 , \unit_decode/n2603 , \unit_decode/n2602 ,
         \unit_decode/n2601 , \unit_decode/n2600 , \unit_decode/n2599 ,
         \unit_decode/n2598 , \unit_decode/n2597 , \unit_decode/n2596 ,
         \unit_decode/n2595 , \unit_decode/n2594 , \unit_decode/n2593 ,
         \unit_decode/n2592 , \unit_decode/n2591 , \unit_decode/n2590 ,
         \unit_decode/n2589 , \unit_decode/n2588 , \unit_decode/n2587 ,
         \unit_decode/n2586 , \unit_decode/n2585 , \unit_decode/n2584 ,
         \unit_decode/n2583 , \unit_decode/n2582 , \unit_decode/n2581 ,
         \unit_decode/n2580 , \unit_decode/n2579 , \unit_decode/n2578 ,
         \unit_decode/n2577 , \unit_decode/n2576 , \unit_decode/n2575 ,
         \unit_decode/n2574 , \unit_decode/n2573 , \unit_decode/n2572 ,
         \unit_decode/n2571 , \unit_decode/n2570 , \unit_decode/n2569 ,
         \unit_decode/n2568 , \unit_decode/n2567 , \unit_decode/n2566 ,
         \unit_decode/n2565 , \unit_decode/n2564 , \unit_decode/n2563 ,
         \unit_decode/n2562 , \unit_decode/n2561 , \unit_decode/n2560 ,
         \unit_decode/n2559 , \unit_decode/n2558 , \unit_decode/n2557 ,
         \unit_decode/n2556 , \unit_decode/n2555 , \unit_decode/n2554 ,
         \unit_decode/n2553 , \unit_decode/n2552 , \unit_decode/n2551 ,
         \unit_decode/n2550 , \unit_decode/n2549 , \unit_decode/n2548 ,
         \unit_decode/n2547 , \unit_decode/n2546 , \unit_decode/n2545 ,
         \unit_decode/n2544 , \unit_decode/n2543 , \unit_decode/n2542 ,
         \unit_decode/n2541 , \unit_decode/n2540 , \unit_decode/n2539 ,
         \unit_decode/n2538 , \unit_decode/n2537 , \unit_decode/n2536 ,
         \unit_decode/n2535 , \unit_decode/n2534 , \unit_decode/n2533 ,
         \unit_decode/n2532 , \unit_decode/n2531 , \unit_decode/n2530 ,
         \unit_decode/n2529 , \unit_decode/n2528 , \unit_decode/n2527 ,
         \unit_decode/n2526 , \unit_decode/n2525 , \unit_decode/n2524 ,
         \unit_decode/n2523 , \unit_decode/n2522 , \unit_decode/n2521 ,
         \unit_decode/n2520 , \unit_decode/n2519 , \unit_decode/n2518 ,
         \unit_decode/n2517 , \unit_decode/n2516 , \unit_decode/n2515 ,
         \unit_decode/n2514 , \unit_decode/n2513 , \unit_decode/n2512 ,
         \unit_decode/n2511 , \unit_decode/n2510 , \unit_decode/n2509 ,
         \unit_decode/n2508 , \unit_decode/n2507 , \unit_decode/n2506 ,
         \unit_decode/n2505 , \unit_decode/n2504 , \unit_decode/n2503 ,
         \unit_decode/n2502 , \unit_decode/n2501 , \unit_decode/n2500 ,
         \unit_decode/n2499 , \unit_decode/n2498 , \unit_decode/n2497 ,
         \unit_decode/n2496 , \unit_decode/n2495 , \unit_decode/n2494 ,
         \unit_decode/n2493 , \unit_decode/n2492 , \unit_decode/n2491 ,
         \unit_decode/n2490 , \unit_decode/n2489 , \unit_decode/n2488 ,
         \unit_decode/n2487 , \unit_decode/n2486 , \unit_decode/n2485 ,
         \unit_decode/n2484 , \unit_decode/n2483 , \unit_decode/n2482 ,
         \unit_decode/n2481 , \unit_decode/n2480 , \unit_decode/n2479 ,
         \unit_decode/n2478 , \unit_decode/n2477 , \unit_decode/n2476 ,
         \unit_decode/n2475 , \unit_decode/n2474 , \unit_decode/n2473 ,
         \unit_decode/n2472 , \unit_decode/n2471 , \unit_decode/n2470 ,
         \unit_decode/n2469 , \unit_decode/n2468 , \unit_decode/n2467 ,
         \unit_decode/n2466 , \unit_decode/n2465 , \unit_decode/n2464 ,
         \unit_decode/n2463 , \unit_decode/n2462 , \unit_decode/n2461 ,
         \unit_decode/n2460 , \unit_decode/n2459 , \unit_decode/n2458 ,
         \unit_decode/n2457 , \unit_decode/n2456 , \unit_decode/n2455 ,
         \unit_decode/n2454 , \unit_decode/n2453 , \unit_decode/n2452 ,
         \unit_decode/n2451 , \unit_decode/n2450 , \unit_decode/n2449 ,
         \unit_decode/n2448 , \unit_decode/n2447 , \unit_decode/n2446 ,
         \unit_decode/n2445 , \unit_decode/n2444 , \unit_decode/n2443 ,
         \unit_decode/n2442 , \unit_decode/n2441 , \unit_decode/n2440 ,
         \unit_decode/n2439 , \unit_decode/n2438 , \unit_decode/n2437 ,
         \unit_decode/n2436 , \unit_decode/n2435 , \unit_decode/n2434 ,
         \unit_decode/n2433 , \unit_decode/n2432 , \unit_decode/n2431 ,
         \unit_decode/n2430 , \unit_decode/n2429 , \unit_decode/n2428 ,
         \unit_decode/n2427 , \unit_decode/n2426 , \unit_decode/n2425 ,
         \unit_decode/n2424 , \unit_decode/n2423 , \unit_decode/n2422 ,
         \unit_decode/n2421 , \unit_decode/n2420 , \unit_decode/n2419 ,
         \unit_decode/n2418 , \unit_decode/n2417 , \unit_decode/n2416 ,
         \unit_decode/n2415 , \unit_decode/n2414 , \unit_decode/n2413 ,
         \unit_decode/n2412 , \unit_decode/n2411 , \unit_decode/n2410 ,
         \unit_decode/n2409 , \unit_decode/n2408 , \unit_decode/n2407 ,
         \unit_decode/n2406 , \unit_decode/n2405 , \unit_decode/n2404 ,
         \unit_decode/n2403 , \unit_decode/n2402 , \unit_decode/n2401 ,
         \unit_decode/n2400 , \unit_decode/n2399 , \unit_decode/n2398 ,
         \unit_decode/n2397 , \unit_decode/n2396 , \unit_decode/n2395 ,
         \unit_decode/n2394 , \unit_decode/n2393 , \unit_decode/n2392 ,
         \unit_decode/n2391 , \unit_decode/n2390 , \unit_decode/n2389 ,
         \unit_decode/n2388 , \unit_decode/n2387 , \unit_decode/n2386 ,
         \unit_decode/n2385 , \unit_decode/n2384 , \unit_decode/n2383 ,
         \unit_decode/n2382 , \unit_decode/n2381 , \unit_decode/n2380 ,
         \unit_decode/n2379 , \unit_decode/n2378 , \unit_decode/n2377 ,
         \unit_decode/n2376 , \unit_decode/n2375 , \unit_decode/n2374 ,
         \unit_decode/n2373 , \unit_decode/n2372 , \unit_decode/n2371 ,
         \unit_decode/n2370 , \unit_decode/n2369 , \unit_decode/n2368 ,
         \unit_decode/n2367 , \unit_decode/n2366 , \unit_decode/n2365 ,
         \unit_decode/n2364 , \unit_decode/n2363 , \unit_decode/n2362 ,
         \unit_decode/n2361 , \unit_decode/n2360 , \unit_decode/n2359 ,
         \unit_decode/n2358 , \unit_decode/n2357 , \unit_decode/n2356 ,
         \unit_decode/n2355 , \unit_decode/n2354 , \unit_decode/n2353 ,
         \unit_decode/n2352 , \unit_decode/n2351 , \unit_decode/n2350 ,
         \unit_decode/n2349 , \unit_decode/n2348 , \unit_decode/n2347 ,
         \unit_decode/n2346 , \unit_decode/n2345 , \unit_decode/n2344 ,
         \unit_decode/n2343 , \unit_decode/n2342 , \unit_decode/n2341 ,
         \unit_decode/n2340 , \unit_decode/n2339 , \unit_decode/n2338 ,
         \unit_decode/n2337 , \unit_decode/n2336 , \unit_decode/n2335 ,
         \unit_decode/n2334 , \unit_decode/n2333 , \unit_decode/n2332 ,
         \unit_decode/n2331 , \unit_decode/n2330 , \unit_decode/n2329 ,
         \unit_decode/n2328 , \unit_decode/n2327 , \unit_decode/n2326 ,
         \unit_decode/n2325 , \unit_decode/n2324 , \unit_decode/n2323 ,
         \unit_decode/n2322 , \unit_decode/n2321 , \unit_decode/n2320 ,
         \unit_decode/n2319 , \unit_decode/n2318 , \unit_decode/n2317 ,
         \unit_decode/n2316 , \unit_decode/n2315 , \unit_decode/n2314 ,
         \unit_decode/n2313 , \unit_decode/n2312 , \unit_decode/n2311 ,
         \unit_decode/n2310 , \unit_decode/n2309 , \unit_decode/n2308 ,
         \unit_decode/n2307 , \unit_decode/n2306 , \unit_decode/n2305 ,
         \unit_decode/n2304 , \unit_decode/n2303 , \unit_decode/n2302 ,
         \unit_decode/n2301 , \unit_decode/n2300 , \unit_decode/n2299 ,
         \unit_decode/n2298 , \unit_decode/n2297 , \unit_decode/n2296 ,
         \unit_decode/n2295 , \unit_decode/n2294 , \unit_decode/n2293 ,
         \unit_decode/n2292 , \unit_decode/n2291 , \unit_decode/n2290 ,
         \unit_decode/n2289 , \unit_decode/n2288 , \unit_decode/n2287 ,
         \unit_decode/n2286 , \unit_decode/n2285 , \unit_decode/n2284 ,
         \unit_decode/n2283 , \unit_decode/n2282 , \unit_decode/n2281 ,
         \unit_decode/n2280 , \unit_decode/n2279 , \unit_decode/n2278 ,
         \unit_decode/n2277 , \unit_decode/n2276 , \unit_decode/n2275 ,
         \unit_decode/n2274 , \unit_decode/n2273 , \unit_decode/n2272 ,
         \unit_decode/n2271 , \unit_decode/n2270 , \unit_decode/n2269 ,
         \unit_decode/n2268 , \unit_decode/n2267 , \unit_decode/n2266 ,
         \unit_decode/n2265 , \unit_decode/n2264 , \unit_decode/n2263 ,
         \unit_decode/n2262 , \unit_decode/n2261 , \unit_decode/n2260 ,
         \unit_decode/n2259 , \unit_decode/n2258 , \unit_decode/n2257 ,
         \unit_decode/n2256 , \unit_decode/n2255 , \unit_decode/n2254 ,
         \unit_decode/n2253 , \unit_decode/n2252 , \unit_decode/n2251 ,
         \unit_decode/n2250 , \unit_decode/n2249 , \unit_decode/n2248 ,
         \unit_decode/n2247 , \unit_decode/n2246 , \unit_decode/n2245 ,
         \unit_decode/n2244 , \unit_decode/n2243 , \unit_decode/n2242 ,
         \unit_decode/n2241 , \unit_decode/n2240 , \unit_decode/n2239 ,
         \unit_decode/n2238 , \unit_decode/n2237 , \unit_decode/n2236 ,
         \unit_decode/n2235 , \unit_decode/n2234 , \unit_decode/n2233 ,
         \unit_decode/n2232 , \unit_decode/n2231 , \unit_decode/n2230 ,
         \unit_decode/n2229 , \unit_decode/n2228 , \unit_decode/n2227 ,
         \unit_decode/n2226 , \unit_decode/n2225 , \unit_decode/n2224 ,
         \unit_decode/n2223 , \unit_decode/n2222 , \unit_decode/n2221 ,
         \unit_decode/n2220 , \unit_decode/n2219 , \unit_decode/n2218 ,
         \unit_decode/n2217 , \unit_decode/n2216 , \unit_decode/n2215 ,
         \unit_decode/n2214 , \unit_decode/n2213 , \unit_decode/n2212 ,
         \unit_decode/n2211 , \unit_decode/n2210 , \unit_decode/n2209 ,
         \unit_decode/n2208 , \unit_decode/n2207 , \unit_decode/n2206 ,
         \unit_decode/n2205 , \unit_decode/n2204 , \unit_decode/n2203 ,
         \unit_decode/n2202 , \unit_decode/n2201 , \unit_decode/n2200 ,
         \unit_decode/n2199 , \unit_decode/n2198 , \unit_decode/n2197 ,
         \unit_decode/n2196 , \unit_decode/n2195 , \unit_decode/n2194 ,
         \unit_decode/n2193 , \unit_decode/n2192 , \unit_decode/n2191 ,
         \unit_decode/n2190 , \unit_decode/n2189 , \unit_decode/n2186 ,
         \unit_decode/n2185 , \unit_decode/n2184 , \unit_decode/n2183 ,
         \unit_decode/n2182 , \unit_decode/n2165 , \unit_decode/n2147 ,
         \unit_decode/n2146 , \unit_decode/n2145 , \unit_decode/n2144 ,
         \unit_decode/n2143 , \unit_decode/n2142 , \unit_decode/n2141 ,
         \unit_decode/n2140 , \unit_decode/n2139 , \unit_decode/n2138 ,
         \unit_decode/n2137 , \unit_decode/n2136 , \unit_decode/n2135 ,
         \unit_decode/n2134 , \unit_decode/n2133 , \unit_decode/n2132 ,
         \unit_decode/n2131 , \unit_decode/n2130 , \unit_decode/n2129 ,
         \unit_decode/n2128 , \unit_decode/n2127 , \unit_decode/n2126 ,
         \unit_decode/n2125 , \unit_decode/n2124 , \unit_decode/n2123 ,
         \unit_decode/n2122 , \unit_decode/n2121 , \unit_decode/n2120 ,
         \unit_decode/n2119 , \unit_decode/n2118 , \unit_decode/n2117 ,
         \unit_decode/n2116 , \unit_decode/n2115 , \unit_decode/n2114 ,
         \unit_decode/n2113 , \unit_decode/n2112 , \unit_decode/n2111 ,
         \unit_decode/n2110 , \unit_decode/n2109 , \unit_decode/n2108 ,
         \unit_decode/n2107 , \unit_decode/n2106 , \unit_decode/n2105 ,
         \unit_decode/n2104 , \unit_decode/n2103 , \unit_decode/n2102 ,
         \unit_decode/n2101 , \unit_decode/n2100 , \unit_decode/n2099 ,
         \unit_decode/n2098 , \unit_decode/n2097 , \unit_decode/n2096 ,
         \unit_decode/n2095 , \unit_decode/n2094 , \unit_decode/n2093 ,
         \unit_decode/n2092 , \unit_decode/n2091 , \unit_decode/n2090 ,
         \unit_decode/n2084 , \unit_decode/n2083 , \unit_decode/n2082 ,
         \unit_decode/n2081 , \unit_decode/n2080 , \unit_decode/n2079 ,
         \unit_decode/n2078 , \unit_decode/n2077 , \unit_decode/n2076 ,
         \unit_decode/n2075 , \unit_decode/n2074 , \unit_decode/n2073 ,
         \unit_decode/n2072 , \unit_decode/n2071 , \unit_decode/n2070 ,
         \unit_decode/n2069 , \unit_decode/n2068 , \unit_decode/n2067 ,
         \unit_decode/n2066 , \unit_decode/n2065 , \unit_decode/n2064 ,
         \unit_decode/n2063 , \unit_decode/n2062 , \unit_decode/n2061 ,
         \unit_decode/n2060 , \unit_decode/n2059 , \unit_decode/n2058 ,
         \unit_decode/n2057 , \unit_decode/n2056 , \unit_decode/n2055 ,
         \unit_decode/n2054 , \unit_decode/n2053 , \unit_decode/n2052 ,
         \unit_decode/n2051 , \unit_decode/n2050 , \unit_decode/n2049 ,
         \unit_decode/n2048 , \unit_decode/n2047 , \unit_decode/n2046 ,
         \unit_decode/n2045 , \unit_decode/n2044 , \unit_decode/n2043 ,
         \unit_decode/n2042 , \unit_decode/n2041 , \unit_decode/n2040 ,
         \unit_decode/n2039 , \unit_decode/n2038 , \unit_decode/n2037 ,
         \unit_decode/n2036 , \unit_decode/n2035 , \unit_decode/n2034 ,
         \unit_decode/n2033 , \unit_decode/n2032 , \unit_decode/n2031 ,
         \unit_decode/n2030 , \unit_decode/n2029 , \unit_decode/n2028 ,
         \unit_decode/n2027 , \unit_decode/n2026 , \unit_decode/n2025 ,
         \unit_decode/n2024 , \unit_decode/n2023 , \unit_decode/n2022 ,
         \unit_decode/n2021 , \unit_decode/n2020 , \unit_decode/n2019 ,
         \unit_decode/n2018 , \unit_decode/n2017 , \unit_decode/n2016 ,
         \unit_decode/n2015 , \unit_decode/n2014 , \unit_decode/n2013 ,
         \unit_decode/n2012 , \unit_decode/n2011 , \unit_decode/n2010 ,
         \unit_decode/n2009 , \unit_decode/n2008 , \unit_decode/n2007 ,
         \unit_decode/n2006 , \unit_decode/n2005 , \unit_decode/n2004 ,
         \unit_decode/n2003 , \unit_decode/n2002 , \unit_decode/n2001 ,
         \unit_decode/n2000 , \unit_decode/n1999 , \unit_decode/n1998 ,
         \unit_decode/n1997 , \unit_decode/n1996 , \unit_decode/n1995 ,
         \unit_decode/n1994 , \unit_decode/n1993 , \unit_decode/n1992 ,
         \unit_decode/n1991 , \unit_decode/n1990 , \unit_decode/n1989 ,
         \unit_decode/n1988 , \unit_decode/n1987 , \unit_decode/n1986 ,
         \unit_decode/n1985 , \unit_decode/n1984 , \unit_decode/n1983 ,
         \unit_decode/n1982 , \unit_decode/n1981 , \unit_decode/n1980 ,
         \unit_decode/n1979 , \unit_decode/n1978 , \unit_decode/n1977 ,
         \unit_decode/n1976 , \unit_decode/n1975 , \unit_decode/n1974 ,
         \unit_decode/n1973 , \unit_decode/n1972 , \unit_decode/n1971 ,
         \unit_decode/n1970 , \unit_decode/n1969 , \unit_decode/n1968 ,
         \unit_decode/n1967 , \unit_decode/n1966 , \unit_decode/n1965 ,
         \unit_decode/n1964 , \unit_decode/n1963 , \unit_decode/n1962 ,
         \unit_decode/n1961 , \unit_decode/n1960 , \unit_decode/n1959 ,
         \unit_decode/n1958 , \unit_decode/n1957 , \unit_decode/n1956 ,
         \unit_decode/n1955 , \unit_decode/n1954 , \unit_decode/n1953 ,
         \unit_decode/n1952 , \unit_decode/n1951 , \unit_decode/n1950 ,
         \unit_decode/n1949 , \unit_decode/n1948 , \unit_decode/n1947 ,
         \unit_decode/n1946 , \unit_decode/n1945 , \unit_decode/n1944 ,
         \unit_decode/n1943 , \unit_decode/n1942 , \unit_decode/n1941 ,
         \unit_decode/n1940 , \unit_decode/n1939 , \unit_decode/n1938 ,
         \unit_decode/n1937 , \unit_decode/n1936 , \unit_decode/n1935 ,
         \unit_decode/n1934 , \unit_decode/n1933 , \unit_decode/n1932 ,
         \unit_decode/n1931 , \unit_decode/n1930 , \unit_decode/n1929 ,
         \unit_decode/n1928 , \unit_decode/n1927 , \unit_decode/n1926 ,
         \unit_decode/n1925 , \unit_decode/n1924 , \unit_decode/n1923 ,
         \unit_decode/n1922 , \unit_decode/n1921 , \unit_decode/n1920 ,
         \unit_decode/n1919 , \unit_decode/n1918 , \unit_decode/n1917 ,
         \unit_decode/n1916 , \unit_decode/n1915 , \unit_decode/n1914 ,
         \unit_decode/n1913 , \unit_decode/n1912 , \unit_decode/n1911 ,
         \unit_decode/n1910 , \unit_decode/n1909 , \unit_decode/n1908 ,
         \unit_decode/n1907 , \unit_decode/n1906 , \unit_decode/n1905 ,
         \unit_decode/n1904 , \unit_decode/n1903 , \unit_decode/n1902 ,
         \unit_decode/n1901 , \unit_decode/n1900 , \unit_decode/n1899 ,
         \unit_decode/n1898 , \unit_decode/n1897 , \unit_decode/n1896 ,
         \unit_decode/n1895 , \unit_decode/n1894 , \unit_decode/n1893 ,
         \unit_decode/n1892 , \unit_decode/n1891 , \unit_decode/n1890 ,
         \unit_decode/n1889 , \unit_decode/n1888 , \unit_decode/n1887 ,
         \unit_decode/n1886 , \unit_decode/n1885 , \unit_decode/n1884 ,
         \unit_decode/n1883 , \unit_decode/n1882 , \unit_decode/n1881 ,
         \unit_decode/n1880 , \unit_decode/n1879 , \unit_decode/n1878 ,
         \unit_decode/n1877 , \unit_decode/n1876 , \unit_decode/n1875 ,
         \unit_decode/n1874 , \unit_decode/n1873 , \unit_decode/n1872 ,
         \unit_decode/n1871 , \unit_decode/n1870 , \unit_decode/n1869 ,
         \unit_decode/n1868 , \unit_decode/n1867 , \unit_decode/n1866 ,
         \unit_decode/n1865 , \unit_decode/n1864 , \unit_decode/n1863 ,
         \unit_decode/n1862 , \unit_decode/n1861 , \unit_decode/n1860 ,
         \unit_decode/n1859 , \unit_decode/n1858 , \unit_decode/n1857 ,
         \unit_decode/n1856 , \unit_decode/n1855 , \unit_decode/n1854 ,
         \unit_decode/n1853 , \unit_decode/n1852 , \unit_decode/n1851 ,
         \unit_decode/n1850 , \unit_decode/n1849 , \unit_decode/n1848 ,
         \unit_decode/n1847 , \unit_decode/n1846 , \unit_decode/n1845 ,
         \unit_decode/n1844 , \unit_decode/n1843 , \unit_decode/n1842 ,
         \unit_decode/n1841 , \unit_decode/n1840 , \unit_decode/n1839 ,
         \unit_decode/n1838 , \unit_decode/n1837 , \unit_decode/n1836 ,
         \unit_decode/n1835 , \unit_decode/n1834 , \unit_decode/n1833 ,
         \unit_decode/n1832 , \unit_decode/n1831 , \unit_decode/n1830 ,
         \unit_decode/n1829 , \unit_decode/n1828 , \unit_decode/n1827 ,
         \unit_decode/n1826 , \unit_decode/n1825 , \unit_decode/n1824 ,
         \unit_decode/n1823 , \unit_decode/n1822 , \unit_decode/n1821 ,
         \unit_decode/n1820 , \unit_decode/n1819 , \unit_decode/n1818 ,
         \unit_decode/n1817 , \unit_decode/n1816 , \unit_decode/n1815 ,
         \unit_decode/n1814 , \unit_decode/n1813 , \unit_decode/n1812 ,
         \unit_decode/n1811 , \unit_decode/n1810 , \unit_decode/n1809 ,
         \unit_decode/n1808 , \unit_decode/n1807 , \unit_decode/n1806 ,
         \unit_decode/n1805 , \unit_decode/n1804 , \unit_decode/n1803 ,
         \unit_decode/n1802 , \unit_decode/n1801 , \unit_decode/n1800 ,
         \unit_decode/n1799 , \unit_decode/n1798 , \unit_decode/n1797 ,
         \unit_decode/n1796 , \unit_decode/n1795 , \unit_decode/n1794 ,
         \unit_decode/n1793 , \unit_decode/n1792 , \unit_decode/n1791 ,
         \unit_decode/n1790 , \unit_decode/n1789 , \unit_decode/n1788 ,
         \unit_decode/n1787 , \unit_decode/n1786 , \unit_decode/n1785 ,
         \unit_decode/n1784 , \unit_decode/n1783 , \unit_decode/n1782 ,
         \unit_decode/n1781 , \unit_decode/n1780 , \unit_decode/n1779 ,
         \unit_decode/n1778 , \unit_decode/n1777 , \unit_decode/n1776 ,
         \unit_decode/n1775 , \unit_decode/n1774 , \unit_decode/n1773 ,
         \unit_decode/n1772 , \unit_decode/n1771 , \unit_decode/n1770 ,
         \unit_decode/n1769 , \unit_decode/n1768 , \unit_decode/n1767 ,
         \unit_decode/n1766 , \unit_decode/n1765 , \unit_decode/n1764 ,
         \unit_decode/n1763 , \unit_decode/n1762 , \unit_decode/n1761 ,
         \unit_decode/n1760 , \unit_decode/n1759 , \unit_decode/n1758 ,
         \unit_decode/n1757 , \unit_decode/n1756 , \unit_decode/n1755 ,
         \unit_decode/n1754 , \unit_decode/n1753 , \unit_decode/n1752 ,
         \unit_decode/n1751 , \unit_decode/n1750 , \unit_decode/n1749 ,
         \unit_decode/n1748 , \unit_decode/n1747 , \unit_decode/n1746 ,
         \unit_decode/n1745 , \unit_decode/n1744 , \unit_decode/n1743 ,
         \unit_decode/n1742 , \unit_decode/n1741 , \unit_decode/n1740 ,
         \unit_decode/n1739 , \unit_decode/n1738 , \unit_decode/n1737 ,
         \unit_decode/n1736 , \unit_decode/n1735 , \unit_decode/n1734 ,
         \unit_decode/n1733 , \unit_decode/n1732 , \unit_decode/n1731 ,
         \unit_decode/n1730 , \unit_decode/n1729 , \unit_decode/n1728 ,
         \unit_decode/n1727 , \unit_decode/n1726 , \unit_decode/n1725 ,
         \unit_decode/n1724 , \unit_decode/n1723 , \unit_decode/n1722 ,
         \unit_decode/n1721 , \unit_decode/n1720 , \unit_decode/n1719 ,
         \unit_decode/n1718 , \unit_decode/n1717 , \unit_decode/n1716 ,
         \unit_decode/n1715 , \unit_decode/n1714 , \unit_decode/n1713 ,
         \unit_decode/n1712 , \unit_decode/n1711 , \unit_decode/n1710 ,
         \unit_decode/n1709 , \unit_decode/n1708 , \unit_decode/n1707 ,
         \unit_decode/n1706 , \unit_decode/n1705 , \unit_decode/n1704 ,
         \unit_decode/n1703 , \unit_decode/n1702 , \unit_decode/n1701 ,
         \unit_decode/n1700 , \unit_decode/n1699 , \unit_decode/n1698 ,
         \unit_decode/n1697 , \unit_decode/n1696 , \unit_decode/n1695 ,
         \unit_decode/n1694 , \unit_decode/n1693 , \unit_decode/n1692 ,
         \unit_decode/n1691 , \unit_decode/n1690 , \unit_decode/n1689 ,
         \unit_decode/n1688 , \unit_decode/n1687 , \unit_decode/n1686 ,
         \unit_decode/n1685 , \unit_decode/n1684 , \unit_decode/n1683 ,
         \unit_decode/n1682 , \unit_decode/n1681 , \unit_decode/n1680 ,
         \unit_decode/n1679 , \unit_decode/n1678 , \unit_decode/n1677 ,
         \unit_decode/n1676 , \unit_decode/n1675 , \unit_decode/n1674 ,
         \unit_decode/n1673 , \unit_decode/n1672 , \unit_decode/n1671 ,
         \unit_decode/n1670 , \unit_decode/n1669 , \unit_decode/n1668 ,
         \unit_decode/n1667 , \unit_decode/n1666 , \unit_decode/n1665 ,
         \unit_decode/n1664 , \unit_decode/n1663 , \unit_decode/n1662 ,
         \unit_decode/n1661 , \unit_decode/n1660 , \unit_decode/n1659 ,
         \unit_decode/n1658 , \unit_decode/n1657 , \unit_decode/n1656 ,
         \unit_decode/n1655 , \unit_decode/n1654 , \unit_decode/n1653 ,
         \unit_decode/n1652 , \unit_decode/n1651 , \unit_decode/n1650 ,
         \unit_decode/n1649 , \unit_decode/n1648 , \unit_decode/n1647 ,
         \unit_decode/n1646 , \unit_decode/n1645 , \unit_decode/n1644 ,
         \unit_decode/n1643 , \unit_decode/n1642 , \unit_decode/n1641 ,
         \unit_decode/n1640 , \unit_decode/n1639 , \unit_decode/n1638 ,
         \unit_decode/n1637 , \unit_decode/n1636 , \unit_decode/n1635 ,
         \unit_decode/n1634 , \unit_decode/n1633 , \unit_decode/n1632 ,
         \unit_decode/n1631 , \unit_decode/n1630 , \unit_decode/n1629 ,
         \unit_decode/n1628 , \unit_decode/n1627 , \unit_decode/n1626 ,
         \unit_decode/n1625 , \unit_decode/n1624 , \unit_decode/n1623 ,
         \unit_decode/n1622 , \unit_decode/n1621 , \unit_decode/n1620 ,
         \unit_decode/n1619 , \unit_decode/n1618 , \unit_decode/n1617 ,
         \unit_decode/n1616 , \unit_decode/n1615 , \unit_decode/n1614 ,
         \unit_decode/n1613 , \unit_decode/n1612 , \unit_decode/n1611 ,
         \unit_decode/n1610 , \unit_decode/n1609 , \unit_decode/n1608 ,
         \unit_decode/n1607 , \unit_decode/n1606 , \unit_decode/n1605 ,
         \unit_decode/n1604 , \unit_decode/n1603 , \unit_decode/n1602 ,
         \unit_decode/n1601 , \unit_decode/n1600 , \unit_decode/n1599 ,
         \unit_decode/n1598 , \unit_decode/n1597 , \unit_decode/n1596 ,
         \unit_decode/n1595 , \unit_decode/n1594 , \unit_decode/n1593 ,
         \unit_decode/n1592 , \unit_decode/n1591 , \unit_decode/n1590 ,
         \unit_decode/n1589 , \unit_decode/n1588 , \unit_decode/n1587 ,
         \unit_decode/n1586 , \unit_decode/n1585 , \unit_decode/n1584 ,
         \unit_decode/n1583 , \unit_decode/n1582 , \unit_decode/n1581 ,
         \unit_decode/n1580 , \unit_decode/n1579 , \unit_decode/n1578 ,
         \unit_decode/n1577 , \unit_decode/n1576 , \unit_decode/n1575 ,
         \unit_decode/n1574 , \unit_decode/n1573 , \unit_decode/n1572 ,
         \unit_decode/n1571 , \unit_decode/n1570 , \unit_decode/n1569 ,
         \unit_decode/n1568 , \unit_decode/n1567 , \unit_decode/n1566 ,
         \unit_decode/n1565 , \unit_decode/n1564 , \unit_decode/n1563 ,
         \unit_decode/n1562 , \unit_decode/n1561 , \unit_decode/n1560 ,
         \unit_decode/n1559 , \unit_decode/n1558 , \unit_decode/n1557 ,
         \unit_decode/n1556 , \unit_decode/n1555 , \unit_decode/n1554 ,
         \unit_decode/n1553 , \unit_decode/n1552 , \unit_decode/n1551 ,
         \unit_decode/n1550 , \unit_decode/n1549 , \unit_decode/n1548 ,
         \unit_decode/n1547 , \unit_decode/n1546 , \unit_decode/n1545 ,
         \unit_decode/n1544 , \unit_decode/n1543 , \unit_decode/n1542 ,
         \unit_decode/n1541 , \unit_decode/n1540 , \unit_decode/n1539 ,
         \unit_decode/n1538 , \unit_decode/n1537 , \unit_decode/n1536 ,
         \unit_decode/n1535 , \unit_decode/n1534 , \unit_decode/n1533 ,
         \unit_decode/n1532 , \unit_decode/n1531 , \unit_decode/n1530 ,
         \unit_decode/n1529 , \unit_decode/n1528 , \unit_decode/n1527 ,
         \unit_decode/n1526 , \unit_decode/n1525 , \unit_decode/n1524 ,
         \unit_decode/n1523 , \unit_decode/n1522 , \unit_decode/n1521 ,
         \unit_decode/n1520 , \unit_decode/n1519 , \unit_decode/n1518 ,
         \unit_decode/n1517 , \unit_decode/n1516 , \unit_decode/n1515 ,
         \unit_decode/n1514 , \unit_decode/n1513 , \unit_decode/n1512 ,
         \unit_decode/n1511 , \unit_decode/n1510 , \unit_decode/n1509 ,
         \unit_decode/n1508 , \unit_decode/n1507 , \unit_decode/n1506 ,
         \unit_decode/n1505 , \unit_decode/n1504 , \unit_decode/n1503 ,
         \unit_decode/n1502 , \unit_decode/n1501 , \unit_decode/n1500 ,
         \unit_decode/n1499 , \unit_decode/n1498 , \unit_decode/n1497 ,
         \unit_decode/n1496 , \unit_decode/n1495 , \unit_decode/n1494 ,
         \unit_decode/n1493 , \unit_decode/n1492 , \unit_decode/n1491 ,
         \unit_decode/n1490 , \unit_decode/n1489 , \unit_decode/n1488 ,
         \unit_decode/n1487 , \unit_decode/n1486 , \unit_decode/n1485 ,
         \unit_decode/n1484 , \unit_decode/n1483 , \unit_decode/n1482 ,
         \unit_decode/n1481 , \unit_decode/n1480 , \unit_decode/n1479 ,
         \unit_decode/n1478 , \unit_decode/n1477 , \unit_decode/n1476 ,
         \unit_decode/n1475 , \unit_decode/n1474 , \unit_decode/n1473 ,
         \unit_decode/n1472 , \unit_decode/n1471 , \unit_decode/n1470 ,
         \unit_decode/n1469 , \unit_decode/n1468 , \unit_decode/n1467 ,
         \unit_decode/n1466 , \unit_decode/n1465 , \unit_decode/n1464 ,
         \unit_decode/n1463 , \unit_decode/n1462 , \unit_decode/n1461 ,
         \unit_decode/n1460 , \unit_decode/n1459 , \unit_decode/n1458 ,
         \unit_decode/n1457 , \unit_decode/n1456 , \unit_decode/n1455 ,
         \unit_decode/n1454 , \unit_decode/n1453 , \unit_decode/n1452 ,
         \unit_decode/n1451 , \unit_decode/n1450 , \unit_decode/n1449 ,
         \unit_decode/n1448 , \unit_decode/n1447 , \unit_decode/n1446 ,
         \unit_decode/n1445 , \unit_decode/n1444 , \unit_decode/n1443 ,
         \unit_decode/n1442 , \unit_decode/n1441 , \unit_decode/n1440 ,
         \unit_decode/n1439 , \unit_decode/n1438 , \unit_decode/n1437 ,
         \unit_decode/n1436 , \unit_decode/n1435 , \unit_decode/n1434 ,
         \unit_decode/n1433 , \unit_decode/n1432 , \unit_decode/n1431 ,
         \unit_decode/n1430 , \unit_decode/n1429 , \unit_decode/n1428 ,
         \unit_decode/n1427 , \unit_decode/n1426 , \unit_decode/n1425 ,
         \unit_decode/n1424 , \unit_decode/n1423 , \unit_decode/n1422 ,
         \unit_decode/n1421 , \unit_decode/n1420 , \unit_decode/n1419 ,
         \unit_decode/n1418 , \unit_decode/n1417 , \unit_decode/n1416 ,
         \unit_decode/n1415 , \unit_decode/n1414 , \unit_decode/n1413 ,
         \unit_decode/n1412 , \unit_decode/n1411 , \unit_decode/n1410 ,
         \unit_decode/n1409 , \unit_decode/n1408 , \unit_decode/n1407 ,
         \unit_decode/n1406 , \unit_decode/n1405 , \unit_decode/n1404 ,
         \unit_decode/n1403 , \unit_decode/n1402 , \unit_decode/n1401 ,
         \unit_decode/n1400 , \unit_decode/n1399 , \unit_decode/n1398 ,
         \unit_decode/n1397 , \unit_decode/n1396 , \unit_decode/n1395 ,
         \unit_decode/n1394 , \unit_decode/n1393 , \unit_decode/n1392 ,
         \unit_decode/n1391 , \unit_decode/n1390 , \unit_decode/n1389 ,
         \unit_decode/n1388 , \unit_decode/n1387 , \unit_decode/n1386 ,
         \unit_decode/n1385 , \unit_decode/n1384 , \unit_decode/n1383 ,
         \unit_decode/n1382 , \unit_decode/n1381 , \unit_decode/n1380 ,
         \unit_decode/n1379 , \unit_decode/n1378 , \unit_decode/n1377 ,
         \unit_decode/n1376 , \unit_decode/n1375 , \unit_decode/n1374 ,
         \unit_decode/n1373 , \unit_decode/n1372 , \unit_decode/n1371 ,
         \unit_decode/n1370 , \unit_decode/n1369 , \unit_decode/n1368 ,
         \unit_decode/n1367 , \unit_decode/n1366 , \unit_decode/n1365 ,
         \unit_decode/n1364 , \unit_decode/n1363 , \unit_decode/n1362 ,
         \unit_decode/n1361 , \unit_decode/n1360 , \unit_decode/n1359 ,
         \unit_decode/n1358 , \unit_decode/n1357 , \unit_decode/n1356 ,
         \unit_decode/n1355 , \unit_decode/n1354 , \unit_decode/n1353 ,
         \unit_decode/n1352 , \unit_decode/n1351 , \unit_decode/n1350 ,
         \unit_decode/n1349 , \unit_decode/n1348 , \unit_decode/n1347 ,
         \unit_decode/n1346 , \unit_decode/n1345 , \unit_decode/n1344 ,
         \unit_decode/n1343 , \unit_decode/n1342 , \unit_decode/n1341 ,
         \unit_decode/n1340 , \unit_decode/n1339 , \unit_decode/n1338 ,
         \unit_decode/n1337 , \unit_decode/n1336 , \unit_decode/n1335 ,
         \unit_decode/n1334 , \unit_decode/n1333 , \unit_decode/n1332 ,
         \unit_decode/n1331 , \unit_decode/n1330 , \unit_decode/n1329 ,
         \unit_decode/n1328 , \unit_decode/n1327 , \unit_decode/n1326 ,
         \unit_decode/n1325 , \unit_decode/n1324 , \unit_decode/n1323 ,
         \unit_decode/n1322 , \unit_decode/n1321 , \unit_decode/n1320 ,
         \unit_decode/n1319 , \unit_decode/n1318 , \unit_decode/n1317 ,
         \unit_decode/n1316 , \unit_decode/n1315 , \unit_decode/n1314 ,
         \unit_decode/n1313 , \unit_decode/n1312 , \unit_decode/n1311 ,
         \unit_decode/n1310 , \unit_decode/n1309 , \unit_decode/n1308 ,
         \unit_decode/n1307 , \unit_decode/n1306 , \unit_decode/n1305 ,
         \unit_decode/n1304 , \unit_decode/n1303 , \unit_decode/n1302 ,
         \unit_decode/n1301 , \unit_decode/n1300 , \unit_decode/n1299 ,
         \unit_decode/n1298 , \unit_decode/n1297 , \unit_decode/n1296 ,
         \unit_decode/n1295 , \unit_decode/n1294 , \unit_decode/n1293 ,
         \unit_decode/n1292 , \unit_decode/n1291 , \unit_decode/n1290 ,
         \unit_decode/n1289 , \unit_decode/n1288 , \unit_decode/n1287 ,
         \unit_decode/n1286 , \unit_decode/n1285 , \unit_decode/n1284 ,
         \unit_decode/n1283 , \unit_decode/n1282 , \unit_decode/n1281 ,
         \unit_decode/n1280 , \unit_decode/n1279 , \unit_decode/n1278 ,
         \unit_decode/n1277 , \unit_decode/n1276 , \unit_decode/n1275 ,
         \unit_decode/n1274 , \unit_decode/n1273 , \unit_decode/n1272 ,
         \unit_decode/n1271 , \unit_decode/n1270 , \unit_decode/n1269 ,
         \unit_decode/n1268 , \unit_decode/n1267 , \unit_decode/n1266 ,
         \unit_decode/n1265 , \unit_decode/n1264 , \unit_decode/n1263 ,
         \unit_decode/n1262 , \unit_decode/n1261 , \unit_decode/n1260 ,
         \unit_decode/n1259 , \unit_decode/n1258 , \unit_decode/n1257 ,
         \unit_decode/n1256 , \unit_decode/n1255 , \unit_decode/n1254 ,
         \unit_decode/n1253 , \unit_decode/n1252 , \unit_decode/n1251 ,
         \unit_decode/n1250 , \unit_decode/n1249 , \unit_decode/n1248 ,
         \unit_decode/n1247 , \unit_decode/n1246 , \unit_decode/n1245 ,
         \unit_decode/n1244 , \unit_decode/n1243 , \unit_decode/n1242 ,
         \unit_decode/n1241 , \unit_decode/n1240 , \unit_decode/n1239 ,
         \unit_decode/n1238 , \unit_decode/n1237 , \unit_decode/n1236 ,
         \unit_decode/n1235 , \unit_decode/n1234 , \unit_decode/n1233 ,
         \unit_decode/n1232 , \unit_decode/n1231 , \unit_decode/n1230 ,
         \unit_decode/n1229 , \unit_decode/n1228 , \unit_decode/n1227 ,
         \unit_decode/n1226 , \unit_decode/n1225 , \unit_decode/n1224 ,
         \unit_decode/n1223 , \unit_decode/n1222 , \unit_decode/n1221 ,
         \unit_decode/n1220 , \unit_decode/n1219 , \unit_decode/n1218 ,
         \unit_decode/n1217 , \unit_decode/n1216 , \unit_decode/n1215 ,
         \unit_decode/n1214 , \unit_decode/n1213 , \unit_decode/n1212 ,
         \unit_decode/n1211 , \unit_decode/n1210 , \unit_decode/n1209 ,
         \unit_decode/n1208 , \unit_decode/n1207 , \unit_decode/n1206 ,
         \unit_decode/n1205 , \unit_decode/n1204 , \unit_decode/n1203 ,
         \unit_decode/n1202 , \unit_decode/n1201 , \unit_decode/n1200 ,
         \unit_decode/n1199 , \unit_decode/n1198 , \unit_decode/n1197 ,
         \unit_decode/n1196 , \unit_decode/n1195 , \unit_decode/n1194 ,
         \unit_decode/n1193 , \unit_decode/n1192 , \unit_decode/n1191 ,
         \unit_decode/n1190 , \unit_decode/n1189 , \unit_decode/n1188 ,
         \unit_decode/n1187 , \unit_decode/n1186 , \unit_decode/n1185 ,
         \unit_decode/n1184 , \unit_decode/n1183 , \unit_decode/n1182 ,
         \unit_decode/n1181 , \unit_decode/n1180 , \unit_decode/n1179 ,
         \unit_decode/n1178 , \unit_decode/n1177 , \unit_decode/n1176 ,
         \unit_decode/n1175 , \unit_decode/n1174 , \unit_decode/n1173 ,
         \unit_decode/n1172 , \unit_decode/n1171 , \unit_decode/n1170 ,
         \unit_decode/n1169 , \unit_decode/n1168 , \unit_decode/n1167 ,
         \unit_decode/n1166 , \unit_decode/n1165 , \unit_decode/n1164 ,
         \unit_decode/n1163 , \unit_decode/n1162 , \unit_decode/n1161 ,
         \unit_decode/n1160 , \unit_decode/n1159 , \unit_decode/n1158 ,
         \unit_decode/n1157 , \unit_decode/n1156 , \unit_decode/n1155 ,
         \unit_decode/n1154 , \unit_decode/n1153 , \unit_decode/n1152 ,
         \unit_decode/n1151 , \unit_decode/n1150 , \unit_decode/n1149 ,
         \unit_decode/n1148 , \unit_decode/n1147 , \unit_decode/n1146 ,
         \unit_decode/n1145 , \unit_decode/n1144 , \unit_decode/n1143 ,
         \unit_decode/n1142 , \unit_decode/n1141 , \unit_decode/n1140 ,
         \unit_decode/n1139 , \unit_decode/n1138 , \unit_decode/n1137 ,
         \unit_decode/n1136 , \unit_decode/n1135 , \unit_decode/n1134 ,
         \unit_decode/n1133 , \unit_decode/n1132 , \unit_decode/n1131 ,
         \unit_decode/n1130 , \unit_decode/n1129 , \unit_decode/n1128 ,
         \unit_decode/n1127 , \unit_decode/n1126 , \unit_decode/n1125 ,
         \unit_decode/n1124 , \unit_decode/n1123 , \unit_decode/n1122 ,
         \unit_decode/n1121 , \unit_decode/n1120 , \unit_decode/n1119 ,
         \unit_decode/n1118 , \unit_decode/n1117 , \unit_decode/n1116 ,
         \unit_decode/n1115 , \unit_decode/n1114 , \unit_decode/n1113 ,
         \unit_decode/n1112 , \unit_decode/n1111 , \unit_decode/n1110 ,
         \unit_decode/n1109 , \unit_decode/n239 , \unit_decode/n237 ,
         \unit_decode/n235 , \unit_decode/n233 , \unit_decode/n231 ,
         \unit_decode/n229 , \unit_decode/n227 , \unit_decode/n225 ,
         \unit_decode/n223 , \unit_decode/n221 , \unit_decode/n219 ,
         \unit_decode/n217 , \unit_decode/n215 , \unit_decode/n213 ,
         \unit_decode/n211 , \unit_decode/n209 , \unit_decode/n207 ,
         \unit_decode/n205 , \unit_decode/n203 , \unit_decode/n201 ,
         \unit_decode/n199 , \unit_decode/n197 , \unit_decode/n195 ,
         \unit_decode/n193 , \unit_decode/n192 , \unit_decode/n191 ,
         \unit_decode/n190 , \unit_decode/n189 , \unit_decode/n188 ,
         \unit_decode/n187 , \unit_decode/n186 , \unit_decode/n185 ,
         \unit_decode/n184 , \unit_decode/n183 , \unit_decode/n182 ,
         \unit_decode/n181 , \unit_decode/n180 , \unit_decode/n179 ,
         \unit_decode/n178 , \unit_decode/n177 , \unit_decode/n176 ,
         \unit_decode/n175 , \unit_decode/n174 , \unit_decode/n173 ,
         \unit_decode/n172 , \unit_decode/n171 , \unit_decode/n170 ,
         \unit_decode/n169 , \unit_decode/n166 , \unit_decode/n163 ,
         \unit_decode/n160 , \unit_decode/n157 , \unit_decode/n154 ,
         \unit_decode/n151 , \unit_decode/n148 , \unit_decode/n145 ,
         \unit_decode/n142 , \unit_decode/n139 , \unit_decode/n136 ,
         \unit_decode/n133 , \unit_decode/n130 , \unit_decode/n127 ,
         \unit_decode/n124 , \unit_decode/n121 , \unit_decode/n118 ,
         \unit_decode/n115 , \unit_decode/n112 , \unit_decode/n109 ,
         \unit_decode/n106 , \unit_decode/n103 , \unit_decode/n100 ,
         \unit_decode/n97 , \unit_decode/n96 , \unit_decode/n94 ,
         \unit_decode/n92 , \unit_decode/n90 , \unit_decode/n88 ,
         \unit_decode/n86 , \unit_decode/n84 , \unit_decode/n82 ,
         \unit_decode/n80 , \unit_decode/n78 , \unit_decode/n76 ,
         \unit_decode/n74 , \unit_decode/n72 , \unit_decode/n70 ,
         \unit_decode/n68 , \unit_decode/n66 , \unit_decode/n64 ,
         \unit_decode/n62 , \unit_decode/n60 , \unit_decode/n58 ,
         \unit_decode/n56 , \unit_decode/n54 , \unit_decode/n52 ,
         \unit_decode/n50 , \unit_decode/n24 , \unit_decode/n23 ,
         \unit_decode/n22 , \unit_decode/n21 , \unit_decode/n20 ,
         \unit_decode/n19 , \unit_decode/n18 , \unit_decode/n17 ,
         \unit_decode/n16 , \unit_decode/n15 , \unit_decode/n14 ,
         \unit_decode/n13 , \unit_decode/n12 , \unit_decode/n11 ,
         \unit_decode/n10 , \unit_decode/n9 , \unit_decode/n8 ,
         \unit_decode/n7 , \unit_decode/n6 , \unit_decode/n5 ,
         \unit_decode/n4 , \unit_decode/n3 , \unit_decode/n2 ,
         \unit_decode/n1 , \unit_decode/NPC1reg/ffi_30/n5 ,
         \unit_decode/NPC1reg/ffi_29/n5 , \unit_decode/NPC1reg/ffi_28/n5 ,
         \unit_decode/NPC1reg/ffi_27/n5 , \unit_decode/NPC1reg/ffi_26/n5 ,
         \unit_decode/NPC1reg/ffi_25/n5 , \unit_decode/NPC1reg/ffi_24/n5 ,
         \unit_decode/NPC1reg/ffi_23/n5 , \unit_decode/NPC1reg/ffi_22/n5 ,
         \unit_decode/NPC1reg/ffi_21/n5 , \unit_decode/NPC1reg/ffi_20/n5 ,
         \unit_decode/NPC1reg/ffi_19/n5 , \unit_decode/NPC1reg/ffi_18/n5 ,
         \unit_decode/NPC1reg/ffi_17/n5 , \unit_decode/NPC1reg/ffi_16/n5 ,
         \unit_decode/NPC1reg/ffi_15/n5 , \unit_decode/NPC1reg/ffi_14/n5 ,
         \unit_decode/NPC1reg/ffi_13/n5 , \unit_decode/NPC1reg/ffi_12/n5 ,
         \unit_decode/NPC1reg/ffi_11/n5 , \unit_decode/NPC1reg/ffi_10/n5 ,
         \unit_decode/NPC1reg/ffi_9/n5 , \unit_decode/NPC1reg/ffi_8/n5 ,
         \unit_decode/NPC1reg/ffi_7/n5 , \unit_decode/NPC1reg/ffi_6/n5 ,
         \unit_decode/NPC1reg/ffi_5/n5 , \unit_decode/NPC1reg/ffi_4/n5 ,
         \unit_decode/NPC1reg/ffi_3/n5 , \unit_decode/NPC1reg/ffi_2/n5 ,
         \unit_decode/NPC1reg/ffi_1/n5 , \unit_decode/NPC1reg/ffi_0/n5 ,
         \unit_decode/Areg/ffi_31/n5 , \unit_decode/Areg/ffi_30/n5 ,
         \unit_decode/Areg/ffi_29/n5 , \unit_decode/Areg/ffi_28/n5 ,
         \unit_decode/Areg/ffi_27/n5 , \unit_decode/Areg/ffi_26/n5 ,
         \unit_decode/Areg/ffi_25/n5 , \unit_decode/Areg/ffi_24/n5 ,
         \unit_decode/Areg/ffi_23/n5 , \unit_decode/Areg/ffi_22/n5 ,
         \unit_decode/Areg/ffi_21/n5 , \unit_decode/Areg/ffi_20/n5 ,
         \unit_decode/Areg/ffi_19/n5 , \unit_decode/Areg/ffi_18/n5 ,
         \unit_decode/Areg/ffi_17/n5 , \unit_decode/Areg/ffi_16/n5 ,
         \unit_decode/Areg/ffi_15/n5 , \unit_decode/Areg/ffi_14/n5 ,
         \unit_decode/Areg/ffi_13/n5 , \unit_decode/Areg/ffi_12/n5 ,
         \unit_decode/Areg/ffi_11/n5 , \unit_decode/Areg/ffi_10/n5 ,
         \unit_decode/Areg/ffi_9/n5 , \unit_decode/Areg/ffi_8/n5 ,
         \unit_decode/Areg/ffi_7/n5 , \unit_decode/Areg/ffi_6/n5 ,
         \unit_decode/Areg/ffi_5/n5 , \unit_decode/Areg/ffi_4/n5 ,
         \unit_decode/Areg/ffi_3/n5 , \unit_decode/Areg/ffi_2/n5 ,
         \unit_decode/Areg/ffi_1/n5 , \unit_decode/Areg/ffi_0/n5 ,
         \unit_decode/Breg/ffi_31/n5 , \unit_decode/Breg/ffi_30/n5 ,
         \unit_decode/Breg/ffi_29/n5 , \unit_decode/Breg/ffi_28/n5 ,
         \unit_decode/Breg/ffi_27/n5 , \unit_decode/Breg/ffi_26/n5 ,
         \unit_decode/Breg/ffi_25/n5 , \unit_decode/Breg/ffi_24/n5 ,
         \unit_decode/Breg/ffi_23/n5 , \unit_decode/Breg/ffi_22/n5 ,
         \unit_decode/Breg/ffi_21/n5 , \unit_decode/Breg/ffi_20/n5 ,
         \unit_decode/Breg/ffi_19/n5 , \unit_decode/Breg/ffi_18/n5 ,
         \unit_decode/Breg/ffi_17/n5 , \unit_decode/Breg/ffi_16/n5 ,
         \unit_decode/Breg/ffi_15/n5 , \unit_decode/Breg/ffi_14/n5 ,
         \unit_decode/Breg/ffi_13/n5 , \unit_decode/Breg/ffi_12/n5 ,
         \unit_decode/Breg/ffi_11/n5 , \unit_decode/Breg/ffi_10/n5 ,
         \unit_decode/Breg/ffi_9/n5 , \unit_decode/Breg/ffi_8/n5 ,
         \unit_decode/Breg/ffi_7/n5 , \unit_decode/Breg/ffi_6/n5 ,
         \unit_decode/Breg/ffi_5/n5 , \unit_decode/Breg/ffi_4/n5 ,
         \unit_decode/Breg/ffi_3/n5 , \unit_decode/Breg/ffi_2/n5 ,
         \unit_decode/Breg/ffi_1/n5 , \unit_decode/Breg/ffi_0/n5 ,
         \unit_decode/IMMreg/ffi_31/n5 , \unit_decode/IMMreg/ffi_30/n5 ,
         \unit_decode/IMMreg/ffi_29/n5 , \unit_decode/IMMreg/ffi_28/n5 ,
         \unit_decode/IMMreg/ffi_27/n5 , \unit_decode/IMMreg/ffi_26/n5 ,
         \unit_decode/IMMreg/ffi_25/n5 , \unit_decode/IMMreg/ffi_24/n5 ,
         \unit_decode/IMMreg/ffi_23/n5 , \unit_decode/IMMreg/ffi_22/n5 ,
         \unit_decode/IMMreg/ffi_21/n5 , \unit_decode/IMMreg/ffi_20/n5 ,
         \unit_decode/IMMreg/ffi_19/n5 , \unit_decode/IMMreg/ffi_18/n5 ,
         \unit_decode/IMMreg/ffi_17/n5 , \unit_decode/IMMreg/ffi_16/n5 ,
         \unit_decode/IMMreg/ffi_15/n5 , \unit_decode/IMMreg/ffi_14/n5 ,
         \unit_decode/IMMreg/ffi_13/n5 , \unit_decode/IMMreg/ffi_12/n5 ,
         \unit_decode/IMMreg/ffi_11/n5 , \unit_decode/IMMreg/ffi_10/n5 ,
         \unit_decode/IMMreg/ffi_9/n5 , \unit_decode/IMMreg/ffi_8/n5 ,
         \unit_decode/IMMreg/ffi_7/n5 , \unit_decode/IMMreg/ffi_6/n5 ,
         \unit_decode/IMMreg/ffi_5/n5 , \unit_decode/IMMreg/ffi_4/n5 ,
         \unit_decode/IMMreg/ffi_3/n5 , \unit_decode/IMMreg/ffi_2/n5 ,
         \unit_decode/IMMreg/ffi_1/n5 , \unit_decode/IMMreg/ffi_0/n5 ,
         \unit_decode/RD1reg/ffi_4/n5 , \unit_decode/RD1reg/ffi_3/n5 ,
         \unit_decode/RD1reg/ffi_2/n5 , \unit_decode/RD1reg/ffi_1/n5 ,
         \unit_decode/RD1reg/ffi_0/n5 , \unit_decode/NPC1reg/ffi_31/n5 ,
         \unit_decode/RegisterFile/N379 , \unit_decode/RegisterFile/N380 ,
         \unit_decode/RegisterFile/N381 , \unit_decode/RegisterFile/N382 ,
         \unit_decode/RegisterFile/N383 , \unit_decode/RegisterFile/N384 ,
         \unit_decode/RegisterFile/N385 , \unit_decode/RegisterFile/N386 ,
         \unit_decode/RegisterFile/N387 , \unit_decode/RegisterFile/N388 ,
         \unit_decode/RegisterFile/N389 , \unit_decode/RegisterFile/N390 ,
         \unit_decode/RegisterFile/N391 , \unit_decode/RegisterFile/N392 ,
         \unit_decode/RegisterFile/N393 , \unit_decode/RegisterFile/N394 ,
         \unit_decode/RegisterFile/N395 , \unit_decode/RegisterFile/N396 ,
         \unit_decode/RegisterFile/N397 , \unit_decode/RegisterFile/N398 ,
         \unit_decode/RegisterFile/N399 , \unit_decode/RegisterFile/N400 ,
         \unit_decode/RegisterFile/N401 , \unit_decode/RegisterFile/N402 ,
         \unit_decode/RegisterFile/N403 , \unit_decode/RegisterFile/N404 ,
         \unit_decode/RegisterFile/N405 , \unit_decode/RegisterFile/N406 ,
         \unit_decode/RegisterFile/N407 , \unit_decode/RegisterFile/N408 ,
         \unit_decode/RegisterFile/N409 , \unit_decode/RegisterFile/N410 ,
         \unit_decode/RegisterFile/N412 , \unit_decode/RegisterFile/N413 ,
         \unit_decode/RegisterFile/N414 , \unit_decode/RegisterFile/N415 ,
         \unit_decode/RegisterFile/N416 , \unit_decode/RegisterFile/N417 ,
         \unit_decode/RegisterFile/N418 , \unit_decode/RegisterFile/N419 ,
         \unit_decode/RegisterFile/N420 , \unit_decode/RegisterFile/N421 ,
         \unit_decode/RegisterFile/N422 , \unit_decode/RegisterFile/N423 ,
         \unit_decode/RegisterFile/N424 , \unit_decode/RegisterFile/N425 ,
         \unit_decode/RegisterFile/N426 , \unit_decode/RegisterFile/N427 ,
         \unit_decode/RegisterFile/N428 , \unit_decode/RegisterFile/N429 ,
         \unit_decode/RegisterFile/N430 , \unit_decode/RegisterFile/N431 ,
         \unit_decode/RegisterFile/N432 , \unit_decode/RegisterFile/N433 ,
         \unit_decode/RegisterFile/N434 , \unit_decode/RegisterFile/N435 ,
         \unit_decode/RegisterFile/N436 , \unit_decode/RegisterFile/N437 ,
         \unit_decode/RegisterFile/N438 , \unit_decode/RegisterFile/N439 ,
         \unit_decode/RegisterFile/N440 , \unit_decode/RegisterFile/N441 ,
         \unit_decode/RegisterFile/N442 , \unit_decode/RegisterFile/N443 ,
         \unit_decode/RegisterFile/N444 , \unit_decode/RegisterFile/N445 ,
         \unit_decode/RegisterFile/n1140 , \unit_decode/RegisterFile/n1141 ,
         \unit_decode/RegisterFile/n1142 , \unit_decode/RegisterFile/n1143 ,
         \unit_decode/RegisterFile/n1144 , \unit_decode/RegisterFile/n1145 ,
         \unit_decode/RegisterFile/n1146 , \unit_decode/RegisterFile/n1147 ,
         \unit_decode/RegisterFile/n1148 , \unit_decode/RegisterFile/n1149 ,
         \unit_decode/RegisterFile/n1150 , \unit_decode/RegisterFile/n1151 ,
         \unit_decode/RegisterFile/n1152 , \unit_decode/RegisterFile/n1153 ,
         \unit_decode/RegisterFile/n1154 , \unit_decode/RegisterFile/n1155 ,
         \unit_decode/RegisterFile/n1156 , \unit_decode/RegisterFile/n1157 ,
         \unit_decode/RegisterFile/n1158 , \unit_decode/RegisterFile/n1159 ,
         \unit_decode/RegisterFile/n1160 , \unit_decode/RegisterFile/n1161 ,
         \unit_decode/RegisterFile/n1162 , \unit_decode/RegisterFile/n1163 ,
         \unit_decode/RegisterFile/n1164 , \unit_decode/RegisterFile/n1165 ,
         \unit_decode/RegisterFile/n1166 , \unit_decode/RegisterFile/n1167 ,
         \unit_decode/RegisterFile/n1168 , \unit_decode/RegisterFile/n1169 ,
         \unit_decode/RegisterFile/n1170 , \unit_decode/RegisterFile/n1171 ,
         \unit_decode/RegisterFile/n1172 , \unit_decode/RegisterFile/n1173 ,
         \unit_decode/RegisterFile/n1174 , \unit_decode/RegisterFile/n1175 ,
         \unit_decode/RegisterFile/n1176 , \unit_decode/RegisterFile/n1177 ,
         \unit_decode/RegisterFile/n1178 , \unit_decode/RegisterFile/n1179 ,
         \unit_decode/RegisterFile/n1180 , \unit_decode/RegisterFile/n1181 ,
         \unit_decode/RegisterFile/n1182 , \unit_decode/RegisterFile/n1183 ,
         \unit_decode/RegisterFile/n1184 , \unit_decode/RegisterFile/n1185 ,
         \unit_decode/RegisterFile/n1186 , \unit_decode/RegisterFile/n1187 ,
         \unit_decode/RegisterFile/n1188 , \unit_decode/RegisterFile/n1189 ,
         \unit_decode/RegisterFile/n1190 , \unit_decode/RegisterFile/n1191 ,
         \unit_decode/RegisterFile/n1192 , \unit_decode/RegisterFile/n1193 ,
         \unit_decode/RegisterFile/n1194 , \unit_decode/RegisterFile/n1195 ,
         \unit_decode/RegisterFile/n1196 , \unit_decode/RegisterFile/n1197 ,
         \unit_decode/RegisterFile/n1198 , \unit_decode/RegisterFile/n1199 ,
         \unit_decode/RegisterFile/n1200 , \unit_decode/RegisterFile/n1201 ,
         \unit_decode/RegisterFile/n1202 , \unit_decode/RegisterFile/n1203 ,
         \unit_decode/RegisterFile/n1204 , \unit_decode/RegisterFile/n1205 ,
         \unit_decode/RegisterFile/n1206 , \unit_decode/RegisterFile/n1207 ,
         \unit_decode/RegisterFile/n1208 , \unit_decode/RegisterFile/n1209 ,
         \unit_decode/RegisterFile/n1210 , \unit_decode/RegisterFile/n1211 ,
         \unit_decode/RegisterFile/n1212 , \unit_decode/RegisterFile/n1213 ,
         \unit_decode/RegisterFile/n1214 , \unit_decode/RegisterFile/n1215 ,
         \unit_decode/RegisterFile/n1216 , \unit_decode/RegisterFile/n1217 ,
         \unit_decode/RegisterFile/n1218 , \unit_decode/RegisterFile/n1219 ,
         \unit_decode/RegisterFile/n1220 , \unit_decode/RegisterFile/n1221 ,
         \unit_decode/RegisterFile/n1222 , \unit_decode/RegisterFile/n1223 ,
         \unit_decode/RegisterFile/n1224 , \unit_decode/RegisterFile/n1225 ,
         \unit_decode/RegisterFile/n1226 , \unit_decode/RegisterFile/n1227 ,
         \unit_decode/RegisterFile/n1228 , \unit_decode/RegisterFile/n1229 ,
         \unit_decode/RegisterFile/n1230 , \unit_decode/RegisterFile/n1231 ,
         \unit_decode/RegisterFile/n1232 , \unit_decode/RegisterFile/n1233 ,
         \unit_decode/RegisterFile/n1234 , \unit_decode/RegisterFile/n1235 ,
         \unit_decode/RegisterFile/n1236 , \unit_decode/RegisterFile/n1237 ,
         \unit_decode/RegisterFile/n1238 , \unit_decode/RegisterFile/n1239 ,
         \unit_decode/RegisterFile/n1240 , \unit_decode/RegisterFile/n1241 ,
         \unit_decode/RegisterFile/n1242 , \unit_decode/RegisterFile/n1243 ,
         \unit_decode/RegisterFile/n1244 , \unit_decode/RegisterFile/n1245 ,
         \unit_decode/RegisterFile/n1246 , \unit_decode/RegisterFile/n1247 ,
         \unit_decode/RegisterFile/n1248 , \unit_decode/RegisterFile/n1249 ,
         \unit_decode/RegisterFile/n1250 , \unit_decode/RegisterFile/n1251 ,
         \unit_decode/RegisterFile/n1252 , \unit_decode/RegisterFile/n1253 ,
         \unit_decode/RegisterFile/n1254 , \unit_decode/RegisterFile/n1255 ,
         \unit_decode/RegisterFile/n1256 , \unit_decode/RegisterFile/n1257 ,
         \unit_decode/RegisterFile/n1258 , \unit_decode/RegisterFile/n1259 ,
         \unit_decode/RegisterFile/n1260 , \unit_decode/RegisterFile/n1261 ,
         \unit_decode/RegisterFile/n1262 , \unit_decode/RegisterFile/n1263 ,
         \unit_decode/RegisterFile/n1264 , \unit_decode/RegisterFile/n1265 ,
         \unit_decode/RegisterFile/n1266 , \unit_decode/RegisterFile/n1267 ,
         \unit_decode/RegisterFile/n1268 , \unit_decode/RegisterFile/n1269 ,
         \unit_decode/RegisterFile/n1270 , \unit_decode/RegisterFile/n1271 ,
         \unit_decode/RegisterFile/n1272 , \unit_decode/RegisterFile/n1273 ,
         \unit_decode/RegisterFile/n1274 , \unit_decode/RegisterFile/n1275 ,
         \unit_decode/RegisterFile/n1276 , \unit_decode/RegisterFile/n1277 ,
         \unit_decode/RegisterFile/n1278 , \unit_decode/RegisterFile/n1279 ,
         \unit_decode/RegisterFile/n1280 , \unit_decode/RegisterFile/n1281 ,
         \unit_decode/RegisterFile/n1282 , \unit_decode/RegisterFile/n1283 ,
         \unit_decode/RegisterFile/n1284 , \unit_decode/RegisterFile/n1285 ,
         \unit_decode/RegisterFile/n1286 , \unit_decode/RegisterFile/n1287 ,
         \unit_decode/RegisterFile/n1288 , \unit_decode/RegisterFile/n1289 ,
         \unit_decode/RegisterFile/n1290 , \unit_decode/RegisterFile/n1291 ,
         \unit_decode/RegisterFile/n1292 , \unit_decode/RegisterFile/n1293 ,
         \unit_decode/RegisterFile/n1294 , \unit_decode/RegisterFile/n1295 ,
         \unit_decode/RegisterFile/n1296 , \unit_decode/RegisterFile/n1297 ,
         \unit_decode/RegisterFile/n1298 , \unit_decode/RegisterFile/n1299 ,
         \unit_decode/RegisterFile/n1300 , \unit_decode/RegisterFile/n1301 ,
         \unit_decode/RegisterFile/n1302 , \unit_decode/RegisterFile/n1303 ,
         \unit_decode/RegisterFile/n1304 , \unit_decode/RegisterFile/n1305 ,
         \unit_decode/RegisterFile/n1306 , \unit_decode/RegisterFile/n1307 ,
         \unit_decode/RegisterFile/n1308 , \unit_decode/RegisterFile/n1309 ,
         \unit_decode/RegisterFile/n1310 , \unit_decode/RegisterFile/n1311 ,
         \unit_decode/RegisterFile/n1312 , \unit_decode/RegisterFile/n1313 ,
         \unit_decode/RegisterFile/n1314 , \unit_decode/RegisterFile/n1315 ,
         \unit_decode/RegisterFile/n1316 , \unit_decode/RegisterFile/n1317 ,
         \unit_decode/RegisterFile/n1318 , \unit_decode/RegisterFile/n1319 ,
         \unit_decode/RegisterFile/n1320 , \unit_decode/RegisterFile/n1321 ,
         \unit_decode/RegisterFile/n1322 , \unit_decode/RegisterFile/n1323 ,
         \unit_decode/RegisterFile/n1324 , \unit_decode/RegisterFile/n1325 ,
         \unit_decode/RegisterFile/n1326 , \unit_decode/RegisterFile/n1327 ,
         \unit_decode/RegisterFile/n1328 , \unit_decode/RegisterFile/n1329 ,
         \unit_decode/RegisterFile/n1330 , \unit_decode/RegisterFile/n1331 ,
         \unit_decode/RegisterFile/n1332 , \unit_decode/RegisterFile/n1333 ,
         \unit_decode/RegisterFile/n1334 , \unit_decode/RegisterFile/n1335 ,
         \unit_decode/RegisterFile/n1336 , \unit_decode/RegisterFile/n1337 ,
         \unit_decode/RegisterFile/n1338 , \unit_decode/RegisterFile/n1339 ,
         \unit_decode/RegisterFile/n1340 , \unit_decode/RegisterFile/n1341 ,
         \unit_decode/RegisterFile/n1342 , \unit_decode/RegisterFile/n1343 ,
         \unit_decode/RegisterFile/n1344 , \unit_decode/RegisterFile/n1345 ,
         \unit_decode/RegisterFile/n1346 , \unit_decode/RegisterFile/n1347 ,
         \unit_decode/RegisterFile/n1348 , \unit_decode/RegisterFile/n1349 ,
         \unit_decode/RegisterFile/n1350 , \unit_decode/RegisterFile/n1351 ,
         \unit_decode/RegisterFile/n1352 , \unit_decode/RegisterFile/n1353 ,
         \unit_decode/RegisterFile/n1354 , \unit_decode/RegisterFile/n1355 ,
         \unit_decode/RegisterFile/n1356 , \unit_decode/RegisterFile/n1357 ,
         \unit_decode/RegisterFile/n1358 , \unit_decode/RegisterFile/n1359 ,
         \unit_decode/RegisterFile/n1360 , \unit_decode/RegisterFile/n1361 ,
         \unit_decode/RegisterFile/n1362 , \unit_decode/RegisterFile/n1363 ,
         \unit_decode/RegisterFile/n1364 , \unit_decode/RegisterFile/n1365 ,
         \unit_decode/RegisterFile/n1366 , \unit_decode/RegisterFile/n1367 ,
         \unit_decode/RegisterFile/n1368 , \unit_decode/RegisterFile/n1369 ,
         \unit_decode/RegisterFile/n1370 , \unit_decode/RegisterFile/n1371 ,
         \unit_decode/RegisterFile/n1372 , \unit_decode/RegisterFile/n1373 ,
         \unit_decode/RegisterFile/n1374 , \unit_decode/RegisterFile/n1375 ,
         \unit_decode/RegisterFile/n1376 , \unit_decode/RegisterFile/n1377 ,
         \unit_decode/RegisterFile/n1378 , \unit_decode/RegisterFile/n1379 ,
         \unit_decode/RegisterFile/n1380 , \unit_decode/RegisterFile/n1381 ,
         \unit_decode/RegisterFile/n1382 , \unit_decode/RegisterFile/n1383 ,
         \unit_decode/RegisterFile/n1384 , \unit_decode/RegisterFile/n1385 ,
         \unit_decode/RegisterFile/n1386 , \unit_decode/RegisterFile/n1387 ,
         \unit_decode/RegisterFile/n1388 , \unit_decode/RegisterFile/n1389 ,
         \unit_decode/RegisterFile/n1390 , \unit_decode/RegisterFile/n1391 ,
         \unit_decode/RegisterFile/n1392 , \unit_decode/RegisterFile/n1393 ,
         \unit_decode/RegisterFile/n1394 , \unit_decode/RegisterFile/n1395 ,
         \unit_decode/RegisterFile/n1396 , \unit_decode/RegisterFile/n1397 ,
         \unit_decode/RegisterFile/n1398 , \unit_decode/RegisterFile/n1399 ,
         \unit_decode/RegisterFile/n1400 , \unit_decode/RegisterFile/n1401 ,
         \unit_decode/RegisterFile/n1402 , \unit_decode/RegisterFile/n1403 ,
         \unit_decode/RegisterFile/n1404 , \unit_decode/RegisterFile/n1405 ,
         \unit_decode/RegisterFile/n1406 , \unit_decode/RegisterFile/n1407 ,
         \unit_decode/RegisterFile/n1408 , \unit_decode/RegisterFile/n1409 ,
         \unit_decode/RegisterFile/n1410 , \unit_decode/RegisterFile/n1411 ,
         \unit_decode/RegisterFile/n1412 , \unit_decode/RegisterFile/n1413 ,
         \unit_decode/RegisterFile/n1414 , \unit_decode/RegisterFile/n1415 ,
         \unit_decode/RegisterFile/n1416 , \unit_decode/RegisterFile/n1417 ,
         \unit_decode/RegisterFile/n1418 , \unit_decode/RegisterFile/n1419 ,
         \unit_decode/RegisterFile/n1420 , \unit_decode/RegisterFile/n1421 ,
         \unit_decode/RegisterFile/n1422 , \unit_decode/RegisterFile/n1423 ,
         \unit_decode/RegisterFile/n1424 , \unit_decode/RegisterFile/n1425 ,
         \unit_decode/RegisterFile/n1426 , \unit_decode/RegisterFile/n1427 ,
         \unit_decode/RegisterFile/n1428 , \unit_decode/RegisterFile/n1429 ,
         \unit_decode/RegisterFile/n1430 , \unit_decode/RegisterFile/n1431 ,
         \unit_decode/RegisterFile/n1432 , \unit_decode/RegisterFile/n1433 ,
         \unit_decode/RegisterFile/n1434 , \unit_decode/RegisterFile/n1435 ,
         \unit_decode/RegisterFile/n1436 , \unit_decode/RegisterFile/n1437 ,
         \unit_decode/RegisterFile/n1438 , \unit_decode/RegisterFile/n1439 ,
         \unit_decode/RegisterFile/n1440 , \unit_decode/RegisterFile/n1441 ,
         \unit_decode/RegisterFile/n1442 , \unit_decode/RegisterFile/n1443 ,
         \unit_decode/RegisterFile/n1444 , \unit_decode/RegisterFile/n1445 ,
         \unit_decode/RegisterFile/n1446 , \unit_decode/RegisterFile/n1447 ,
         \unit_decode/RegisterFile/n1448 , \unit_decode/RegisterFile/n1449 ,
         \unit_decode/RegisterFile/n1450 , \unit_decode/RegisterFile/n1451 ,
         \unit_decode/RegisterFile/n1452 , \unit_decode/RegisterFile/n1453 ,
         \unit_decode/RegisterFile/n1454 , \unit_decode/RegisterFile/n1455 ,
         \unit_decode/RegisterFile/n1456 , \unit_decode/RegisterFile/n1457 ,
         \unit_decode/RegisterFile/n1458 , \unit_decode/RegisterFile/n1459 ,
         \unit_decode/RegisterFile/n1460 , \unit_decode/RegisterFile/n1461 ,
         \unit_decode/RegisterFile/n1462 , \unit_decode/RegisterFile/n1463 ,
         \unit_decode/RegisterFile/n1464 , \unit_decode/RegisterFile/n1465 ,
         \unit_decode/RegisterFile/n1466 , \unit_decode/RegisterFile/n1467 ,
         \unit_decode/RegisterFile/n1468 , \unit_decode/RegisterFile/n1469 ,
         \unit_decode/RegisterFile/n1470 , \unit_decode/RegisterFile/n1471 ,
         \unit_decode/RegisterFile/n1472 , \unit_decode/RegisterFile/n1473 ,
         \unit_decode/RegisterFile/n1474 , \unit_decode/RegisterFile/n1475 ,
         \unit_decode/RegisterFile/n1476 , \unit_decode/RegisterFile/n1477 ,
         \unit_decode/RegisterFile/n1478 , \unit_decode/RegisterFile/n1479 ,
         \unit_decode/RegisterFile/n1480 , \unit_decode/RegisterFile/n1481 ,
         \unit_decode/RegisterFile/n1482 , \unit_decode/RegisterFile/n1483 ,
         \unit_decode/RegisterFile/n1484 , \unit_decode/RegisterFile/n1485 ,
         \unit_decode/RegisterFile/n1486 , \unit_decode/RegisterFile/n1487 ,
         \unit_decode/RegisterFile/n1488 , \unit_decode/RegisterFile/n1489 ,
         \unit_decode/RegisterFile/n1490 , \unit_decode/RegisterFile/n1491 ,
         \unit_decode/RegisterFile/n1492 , \unit_decode/RegisterFile/n1493 ,
         \unit_decode/RegisterFile/n1494 , \unit_decode/RegisterFile/n1495 ,
         \unit_decode/RegisterFile/n1496 , \unit_decode/RegisterFile/n1497 ,
         \unit_decode/RegisterFile/n1498 , \unit_decode/RegisterFile/n1499 ,
         \unit_decode/RegisterFile/n1500 , \unit_decode/RegisterFile/n1501 ,
         \unit_decode/RegisterFile/n1502 , \unit_decode/RegisterFile/n1503 ,
         \unit_decode/RegisterFile/n1504 , \unit_decode/RegisterFile/n1505 ,
         \unit_decode/RegisterFile/n1506 , \unit_decode/RegisterFile/n1507 ,
         \unit_decode/RegisterFile/n1508 , \unit_decode/RegisterFile/n1509 ,
         \unit_decode/RegisterFile/n1510 , \unit_decode/RegisterFile/n1511 ,
         \unit_decode/RegisterFile/n1512 , \unit_decode/RegisterFile/n1513 ,
         \unit_decode/RegisterFile/n1514 , \unit_decode/RegisterFile/n1515 ,
         \unit_decode/RegisterFile/n1516 , \unit_decode/RegisterFile/n1517 ,
         \unit_decode/RegisterFile/n1518 , \unit_decode/RegisterFile/n1519 ,
         \unit_decode/RegisterFile/n1520 , \unit_decode/RegisterFile/n1521 ,
         \unit_decode/RegisterFile/n1522 , \unit_decode/RegisterFile/n1523 ,
         \unit_decode/RegisterFile/n1524 , \unit_decode/RegisterFile/n1525 ,
         \unit_decode/RegisterFile/n1526 , \unit_decode/RegisterFile/n1527 ,
         \unit_decode/RegisterFile/n1528 , \unit_decode/RegisterFile/n1529 ,
         \unit_decode/RegisterFile/n1530 , \unit_decode/RegisterFile/n1531 ,
         \unit_decode/RegisterFile/n1532 , \unit_decode/RegisterFile/n1533 ,
         \unit_decode/RegisterFile/n1534 , \unit_decode/RegisterFile/n1535 ,
         \unit_decode/RegisterFile/n1536 , \unit_decode/RegisterFile/n1537 ,
         \unit_decode/RegisterFile/n1538 , \unit_decode/RegisterFile/n1539 ,
         \unit_decode/RegisterFile/n1540 , \unit_decode/RegisterFile/n1541 ,
         \unit_decode/RegisterFile/n1542 , \unit_decode/RegisterFile/n1543 ,
         \unit_decode/RegisterFile/n1544 , \unit_decode/RegisterFile/n1545 ,
         \unit_decode/RegisterFile/n1546 , \unit_decode/RegisterFile/n1547 ,
         \unit_decode/RegisterFile/n1548 , \unit_decode/RegisterFile/n1549 ,
         \unit_decode/RegisterFile/n1550 , \unit_decode/RegisterFile/n1551 ,
         \unit_decode/RegisterFile/n1552 , \unit_decode/RegisterFile/n1553 ,
         \unit_decode/RegisterFile/n1554 , \unit_decode/RegisterFile/n1555 ,
         \unit_decode/RegisterFile/n1556 , \unit_decode/RegisterFile/n1557 ,
         \unit_decode/RegisterFile/n1558 , \unit_decode/RegisterFile/n1559 ,
         \unit_decode/RegisterFile/n1560 , \unit_decode/RegisterFile/n1561 ,
         \unit_decode/RegisterFile/n1562 , \unit_decode/RegisterFile/n1563 ,
         \unit_decode/RegisterFile/n1564 , \unit_decode/RegisterFile/n1565 ,
         \unit_decode/RegisterFile/n1566 , \unit_decode/RegisterFile/n1567 ,
         \unit_decode/RegisterFile/n1568 , \unit_decode/RegisterFile/n1569 ,
         \unit_decode/RegisterFile/n1570 , \unit_decode/RegisterFile/n1571 ,
         \unit_decode/RegisterFile/n1572 , \unit_decode/RegisterFile/n1573 ,
         \unit_decode/RegisterFile/n1574 , \unit_decode/RegisterFile/n1575 ,
         \unit_decode/RegisterFile/n1576 , \unit_decode/RegisterFile/n1577 ,
         \unit_decode/RegisterFile/n1578 , \unit_decode/RegisterFile/n1579 ,
         \unit_decode/RegisterFile/n1580 , \unit_decode/RegisterFile/n1581 ,
         \unit_decode/RegisterFile/n1582 , \unit_decode/RegisterFile/n1583 ,
         \unit_decode/RegisterFile/n1584 , \unit_decode/RegisterFile/n1585 ,
         \unit_decode/RegisterFile/n1586 , \unit_decode/RegisterFile/n1587 ,
         \unit_decode/RegisterFile/n1588 , \unit_decode/RegisterFile/n1589 ,
         \unit_decode/RegisterFile/n1590 , \unit_decode/RegisterFile/n1591 ,
         \unit_decode/RegisterFile/n1592 , \unit_decode/RegisterFile/n1593 ,
         \unit_decode/RegisterFile/n1594 , \unit_decode/RegisterFile/n1595 ,
         \unit_decode/RegisterFile/n1596 , \unit_decode/RegisterFile/n1597 ,
         \unit_decode/RegisterFile/n1598 , \unit_decode/RegisterFile/n1599 ,
         \unit_decode/RegisterFile/n1600 , \unit_decode/RegisterFile/n1601 ,
         \unit_decode/RegisterFile/n1602 , \unit_decode/RegisterFile/n1603 ,
         \unit_decode/RegisterFile/n1604 , \unit_decode/RegisterFile/n1605 ,
         \unit_decode/RegisterFile/n1606 , \unit_decode/RegisterFile/n1607 ,
         \unit_decode/RegisterFile/n1608 , \unit_decode/RegisterFile/n1609 ,
         \unit_decode/RegisterFile/n1610 , \unit_decode/RegisterFile/n1611 ,
         \unit_decode/RegisterFile/n1612 , \unit_decode/RegisterFile/n1613 ,
         \unit_decode/RegisterFile/n1614 , \unit_decode/RegisterFile/n1615 ,
         \unit_decode/RegisterFile/n1616 , \unit_decode/RegisterFile/n1617 ,
         \unit_decode/RegisterFile/n1618 , \unit_decode/RegisterFile/n1619 ,
         \unit_decode/RegisterFile/n1620 , \unit_decode/RegisterFile/n1621 ,
         \unit_decode/RegisterFile/n1622 , \unit_decode/RegisterFile/n1623 ,
         \unit_decode/RegisterFile/n1624 , \unit_decode/RegisterFile/n1625 ,
         \unit_decode/RegisterFile/n1626 , \unit_decode/RegisterFile/n1627 ,
         \unit_decode/RegisterFile/n1628 , \unit_decode/RegisterFile/n1629 ,
         \unit_decode/RegisterFile/n1630 , \unit_decode/RegisterFile/n1631 ,
         \unit_decode/RegisterFile/n1632 , \unit_decode/RegisterFile/n1633 ,
         \unit_decode/RegisterFile/n1634 , \unit_decode/RegisterFile/n1635 ,
         \unit_decode/RegisterFile/n1636 , \unit_decode/RegisterFile/n1637 ,
         \unit_decode/RegisterFile/n1638 , \unit_decode/RegisterFile/n1639 ,
         \unit_decode/RegisterFile/n1640 , \unit_decode/RegisterFile/n1641 ,
         \unit_decode/RegisterFile/n1642 , \unit_decode/RegisterFile/n1643 ,
         \unit_decode/RegisterFile/n1644 , \unit_decode/RegisterFile/n1645 ,
         \unit_decode/RegisterFile/n1646 , \unit_decode/RegisterFile/n1647 ,
         \unit_decode/RegisterFile/n1648 , \unit_decode/RegisterFile/n1649 ,
         \unit_decode/RegisterFile/n1650 , \unit_decode/RegisterFile/n1651 ,
         \unit_decode/RegisterFile/n1652 , \unit_decode/RegisterFile/n1653 ,
         \unit_decode/RegisterFile/n1654 , \unit_decode/RegisterFile/n1655 ,
         \unit_decode/RegisterFile/n1656 , \unit_decode/RegisterFile/n1657 ,
         \unit_decode/RegisterFile/n1658 , \unit_decode/RegisterFile/n1659 ,
         \unit_decode/RegisterFile/n1660 , \unit_decode/RegisterFile/n1661 ,
         \unit_decode/RegisterFile/n1662 , \unit_decode/RegisterFile/n1663 ,
         \unit_decode/RegisterFile/n1664 , \unit_decode/RegisterFile/n1665 ,
         \unit_decode/RegisterFile/n1666 , \unit_decode/RegisterFile/n1667 ,
         \unit_decode/RegisterFile/n1668 , \unit_decode/RegisterFile/n1669 ,
         \unit_decode/RegisterFile/n1670 , \unit_decode/RegisterFile/n1671 ,
         \unit_decode/RegisterFile/n1672 , \unit_decode/RegisterFile/n1673 ,
         \unit_decode/RegisterFile/n1674 , \unit_decode/RegisterFile/n1675 ,
         \unit_decode/RegisterFile/n1676 , \unit_decode/RegisterFile/n1677 ,
         \unit_decode/RegisterFile/n1678 , \unit_decode/RegisterFile/n1679 ,
         \unit_decode/RegisterFile/n1680 , \unit_decode/RegisterFile/n1681 ,
         \unit_decode/RegisterFile/n1682 , \unit_decode/RegisterFile/n1683 ,
         \unit_decode/RegisterFile/n1684 , \unit_decode/RegisterFile/n1685 ,
         \unit_decode/RegisterFile/n1686 , \unit_decode/RegisterFile/n1687 ,
         \unit_decode/RegisterFile/n1688 , \unit_decode/RegisterFile/n1689 ,
         \unit_decode/RegisterFile/n1690 , \unit_decode/RegisterFile/n1691 ,
         \unit_decode/RegisterFile/n1692 , \unit_decode/RegisterFile/n1693 ,
         \unit_decode/RegisterFile/n1694 , \unit_decode/RegisterFile/n1695 ,
         \unit_decode/RegisterFile/n1696 , \unit_decode/RegisterFile/n1697 ,
         \unit_decode/RegisterFile/n1698 , \unit_decode/RegisterFile/n1699 ,
         \unit_decode/RegisterFile/n1700 , \unit_decode/RegisterFile/n1701 ,
         \unit_decode/RegisterFile/n1702 , \unit_decode/RegisterFile/n1703 ,
         \unit_decode/RegisterFile/n1704 , \unit_decode/RegisterFile/n1705 ,
         \unit_decode/RegisterFile/n1706 , \unit_decode/RegisterFile/n1707 ,
         \unit_decode/RegisterFile/n1708 , \unit_decode/RegisterFile/n1709 ,
         \unit_decode/RegisterFile/n1710 , \unit_decode/RegisterFile/n1711 ,
         \unit_decode/RegisterFile/n1712 , \unit_decode/RegisterFile/n1713 ,
         \unit_decode/RegisterFile/n1714 , \unit_decode/RegisterFile/n1715 ,
         \unit_decode/RegisterFile/n1716 , \unit_decode/RegisterFile/n1717 ,
         \unit_decode/RegisterFile/n1718 , \unit_decode/RegisterFile/n1719 ,
         \unit_decode/RegisterFile/n1720 , \unit_decode/RegisterFile/n1721 ,
         \unit_decode/RegisterFile/n1722 , \unit_decode/RegisterFile/n1723 ,
         \unit_decode/RegisterFile/n1724 , \unit_decode/RegisterFile/n1725 ,
         \unit_decode/RegisterFile/n1726 , \unit_decode/RegisterFile/n1727 ,
         \unit_decode/RegisterFile/n1728 , \unit_decode/RegisterFile/n1729 ,
         \unit_decode/RegisterFile/n1730 , \unit_decode/RegisterFile/n1731 ,
         \unit_decode/RegisterFile/n1732 , \unit_decode/RegisterFile/n1733 ,
         \unit_decode/RegisterFile/n1734 , \unit_decode/RegisterFile/n1735 ,
         \unit_decode/RegisterFile/n1736 , \unit_decode/RegisterFile/n1737 ,
         \unit_decode/RegisterFile/n1738 , \unit_decode/RegisterFile/n1739 ,
         \unit_decode/RegisterFile/n1740 , \unit_decode/RegisterFile/n1741 ,
         \unit_decode/RegisterFile/n1742 , \unit_decode/RegisterFile/n1743 ,
         \unit_decode/RegisterFile/n1744 , \unit_decode/RegisterFile/n1745 ,
         \unit_decode/RegisterFile/n1746 , \unit_decode/RegisterFile/n1747 ,
         \unit_decode/RegisterFile/n1748 , \unit_decode/RegisterFile/n1749 ,
         \unit_decode/RegisterFile/n1750 , \unit_decode/RegisterFile/n1751 ,
         \unit_decode/RegisterFile/n1752 , \unit_decode/RegisterFile/n1753 ,
         \unit_decode/RegisterFile/n1754 , \unit_decode/RegisterFile/n1755 ,
         \unit_decode/RegisterFile/n1756 , \unit_decode/RegisterFile/n1757 ,
         \unit_decode/RegisterFile/n1758 , \unit_decode/RegisterFile/n1759 ,
         \unit_decode/RegisterFile/n1760 , \unit_decode/RegisterFile/n1761 ,
         \unit_decode/RegisterFile/n1762 , \unit_decode/RegisterFile/n1763 ,
         \unit_decode/RegisterFile/n1764 , \unit_decode/RegisterFile/n1765 ,
         \unit_decode/RegisterFile/n1766 , \unit_decode/RegisterFile/n1767 ,
         \unit_decode/RegisterFile/n1768 , \unit_decode/RegisterFile/n1769 ,
         \unit_decode/RegisterFile/n1770 , \unit_decode/RegisterFile/n1771 ,
         \unit_decode/RegisterFile/n1772 , \unit_decode/RegisterFile/n1773 ,
         \unit_decode/RegisterFile/n1774 , \unit_decode/RegisterFile/n1775 ,
         \unit_decode/RegisterFile/n1776 , \unit_decode/RegisterFile/n1777 ,
         \unit_decode/RegisterFile/n1778 , \unit_decode/RegisterFile/n1779 ,
         \unit_decode/RegisterFile/n1780 , \unit_decode/RegisterFile/n1781 ,
         \unit_decode/RegisterFile/n1782 , \unit_decode/RegisterFile/n1783 ,
         \unit_decode/RegisterFile/n1784 , \unit_decode/RegisterFile/n1785 ,
         \unit_decode/RegisterFile/n1786 , \unit_decode/RegisterFile/n1787 ,
         \unit_decode/RegisterFile/n1788 , \unit_decode/RegisterFile/n1789 ,
         \unit_decode/RegisterFile/n1790 , \unit_decode/RegisterFile/n1791 ,
         \unit_decode/RegisterFile/n1792 , \unit_decode/RegisterFile/n1793 ,
         \unit_decode/RegisterFile/n1794 , \unit_decode/RegisterFile/n1795 ,
         \unit_decode/RegisterFile/n1796 , \unit_decode/RegisterFile/n1797 ,
         \unit_decode/RegisterFile/n1798 , \unit_decode/RegisterFile/n1799 ,
         \unit_decode/RegisterFile/n1800 , \unit_decode/RegisterFile/n1801 ,
         \unit_decode/RegisterFile/n1802 , \unit_decode/RegisterFile/n1803 ,
         \unit_decode/RegisterFile/n1804 , \unit_decode/RegisterFile/n1805 ,
         \unit_decode/RegisterFile/n1806 , \unit_decode/RegisterFile/n1807 ,
         \unit_decode/RegisterFile/n1808 , \unit_decode/RegisterFile/n1809 ,
         \unit_decode/RegisterFile/n1810 , \unit_decode/RegisterFile/n1811 ,
         \unit_decode/RegisterFile/n1812 , \unit_decode/RegisterFile/n1813 ,
         \unit_decode/RegisterFile/n1814 , \unit_decode/RegisterFile/n1815 ,
         \unit_decode/RegisterFile/n1816 , \unit_decode/RegisterFile/n1817 ,
         \unit_decode/RegisterFile/n1818 , \unit_decode/RegisterFile/n1819 ,
         \unit_decode/RegisterFile/n1820 , \unit_decode/RegisterFile/n1821 ,
         \unit_decode/RegisterFile/n1822 , \unit_decode/RegisterFile/n1823 ,
         \unit_decode/RegisterFile/n1824 , \unit_decode/RegisterFile/n1825 ,
         \unit_decode/RegisterFile/n1826 , \unit_decode/RegisterFile/n1827 ,
         \unit_decode/RegisterFile/n1828 , \unit_decode/RegisterFile/n1829 ,
         \unit_decode/RegisterFile/n1830 , \unit_decode/RegisterFile/n1831 ,
         \unit_decode/RegisterFile/n1832 , \unit_decode/RegisterFile/n1833 ,
         \unit_decode/RegisterFile/n1834 , \unit_decode/RegisterFile/n1835 ,
         \unit_decode/RegisterFile/n1836 , \unit_decode/RegisterFile/n1837 ,
         \unit_decode/RegisterFile/n1838 , \unit_decode/RegisterFile/n1839 ,
         \unit_decode/RegisterFile/n1840 , \unit_decode/RegisterFile/n1841 ,
         \unit_decode/RegisterFile/n1842 , \unit_decode/RegisterFile/n1843 ,
         \unit_decode/RegisterFile/n1844 , \unit_decode/RegisterFile/n1845 ,
         \unit_decode/RegisterFile/n1846 , \unit_decode/RegisterFile/n1847 ,
         \unit_decode/RegisterFile/n1848 , \unit_decode/RegisterFile/n1849 ,
         \unit_decode/RegisterFile/n1850 , \unit_decode/RegisterFile/n1851 ,
         \unit_decode/RegisterFile/n1852 , \unit_decode/RegisterFile/n1853 ,
         \unit_decode/RegisterFile/n1854 , \unit_decode/RegisterFile/n1855 ,
         \unit_decode/RegisterFile/n1856 , \unit_decode/RegisterFile/n1857 ,
         \unit_decode/RegisterFile/n1858 , \unit_decode/RegisterFile/n1859 ,
         \unit_decode/RegisterFile/n1860 , \unit_decode/RegisterFile/n1861 ,
         \unit_decode/RegisterFile/n1862 , \unit_decode/RegisterFile/n1863 ,
         \unit_decode/RegisterFile/n1864 , \unit_decode/RegisterFile/n1865 ,
         \unit_decode/RegisterFile/n1866 , \unit_decode/RegisterFile/n1867 ,
         \unit_decode/RegisterFile/n1868 , \unit_decode/RegisterFile/n1869 ,
         \unit_decode/RegisterFile/n1870 , \unit_decode/RegisterFile/n1871 ,
         \unit_decode/RegisterFile/n1872 , \unit_decode/RegisterFile/n1873 ,
         \unit_decode/RegisterFile/n1874 , \unit_decode/RegisterFile/n1875 ,
         \unit_decode/RegisterFile/n1876 , \unit_decode/RegisterFile/n1877 ,
         \unit_decode/RegisterFile/n1878 , \unit_decode/RegisterFile/n1879 ,
         \unit_decode/RegisterFile/n1880 , \unit_decode/RegisterFile/n1881 ,
         \unit_decode/RegisterFile/n1882 , \unit_decode/RegisterFile/n1883 ,
         \unit_decode/RegisterFile/n1884 , \unit_decode/RegisterFile/n1885 ,
         \unit_decode/RegisterFile/n1886 , \unit_decode/RegisterFile/n1887 ,
         \unit_decode/RegisterFile/n1888 , \unit_decode/RegisterFile/n1889 ,
         \unit_decode/RegisterFile/n1890 , \unit_decode/RegisterFile/n1891 ,
         \unit_decode/RegisterFile/n1892 , \unit_decode/RegisterFile/n1893 ,
         \unit_decode/RegisterFile/n1894 , \unit_decode/RegisterFile/n1895 ,
         \unit_decode/RegisterFile/n1896 , \unit_decode/RegisterFile/n1897 ,
         \unit_decode/RegisterFile/n1898 , \unit_decode/RegisterFile/n1899 ,
         \unit_decode/RegisterFile/n1900 , \unit_decode/RegisterFile/n1901 ,
         \unit_decode/RegisterFile/n1902 , \unit_decode/RegisterFile/n1903 ,
         \unit_decode/RegisterFile/n1904 , \unit_decode/RegisterFile/n1905 ,
         \unit_decode/RegisterFile/n1906 , \unit_decode/RegisterFile/n1907 ,
         \unit_decode/RegisterFile/n1908 , \unit_decode/RegisterFile/n1909 ,
         \unit_decode/RegisterFile/n1910 , \unit_decode/RegisterFile/n1911 ,
         \unit_decode/RegisterFile/n1912 , \unit_decode/RegisterFile/n1913 ,
         \unit_decode/RegisterFile/n1914 , \unit_decode/RegisterFile/n1915 ,
         \unit_decode/RegisterFile/n1916 , \unit_decode/RegisterFile/n1917 ,
         \unit_decode/RegisterFile/n1918 , \unit_decode/RegisterFile/n1919 ,
         \unit_decode/RegisterFile/n1920 , \unit_decode/RegisterFile/n1921 ,
         \unit_decode/RegisterFile/n1922 , \unit_decode/RegisterFile/n1923 ,
         \unit_decode/RegisterFile/n1924 , \unit_decode/RegisterFile/n1925 ,
         \unit_decode/RegisterFile/n1926 , \unit_decode/RegisterFile/n1927 ,
         \unit_decode/RegisterFile/n1928 , \unit_decode/RegisterFile/n1929 ,
         \unit_decode/RegisterFile/n1930 , \unit_decode/RegisterFile/n1931 ,
         \unit_decode/RegisterFile/n1932 , \unit_decode/RegisterFile/n1933 ,
         \unit_decode/RegisterFile/n1934 , \unit_decode/RegisterFile/n1935 ,
         \unit_decode/RegisterFile/n1936 , \unit_decode/RegisterFile/n1937 ,
         \unit_decode/RegisterFile/n1938 , \unit_decode/RegisterFile/n1939 ,
         \unit_decode/RegisterFile/n1940 , \unit_decode/RegisterFile/n1941 ,
         \unit_decode/RegisterFile/n1942 , \unit_decode/RegisterFile/n1943 ,
         \unit_decode/RegisterFile/n1944 , \unit_decode/RegisterFile/n1945 ,
         \unit_decode/RegisterFile/n1946 , \unit_decode/RegisterFile/n1947 ,
         \unit_decode/RegisterFile/n1948 , \unit_decode/RegisterFile/n1949 ,
         \unit_decode/RegisterFile/n1950 , \unit_decode/RegisterFile/n1951 ,
         \unit_decode/RegisterFile/n1952 , \unit_decode/RegisterFile/n1953 ,
         \unit_decode/RegisterFile/n1954 , \unit_decode/RegisterFile/n1955 ,
         \unit_decode/RegisterFile/n1956 , \unit_decode/RegisterFile/n1957 ,
         \unit_decode/RegisterFile/n1958 , \unit_decode/RegisterFile/n1959 ,
         \unit_decode/RegisterFile/n1960 , \unit_decode/RegisterFile/n1961 ,
         \unit_decode/RegisterFile/n1962 , \unit_decode/RegisterFile/n1963 ,
         \unit_decode/RegisterFile/n1964 , \unit_decode/RegisterFile/n1965 ,
         \unit_decode/RegisterFile/n1966 , \unit_decode/RegisterFile/n1967 ,
         \unit_decode/RegisterFile/n1968 , \unit_decode/RegisterFile/n1969 ,
         \unit_decode/RegisterFile/n1970 , \unit_decode/RegisterFile/n1971 ,
         \unit_decode/RegisterFile/n1972 , \unit_decode/RegisterFile/n1973 ,
         \unit_decode/RegisterFile/n1974 , \unit_decode/RegisterFile/n1975 ,
         \unit_decode/RegisterFile/n1976 , \unit_decode/RegisterFile/n1977 ,
         \unit_decode/RegisterFile/n1978 , \unit_decode/RegisterFile/n1979 ,
         \unit_decode/RegisterFile/n1980 , \unit_decode/RegisterFile/n1981 ,
         \unit_decode/RegisterFile/n1982 , \unit_decode/RegisterFile/n1983 ,
         \unit_decode/RegisterFile/n1984 , \unit_decode/RegisterFile/n1985 ,
         \unit_decode/RegisterFile/n1986 , \unit_decode/RegisterFile/n1987 ,
         \unit_decode/RegisterFile/n1988 , \unit_decode/RegisterFile/n1989 ,
         \unit_decode/RegisterFile/n1990 , \unit_decode/RegisterFile/n1991 ,
         \unit_decode/RegisterFile/n1992 , \unit_decode/RegisterFile/n1993 ,
         \unit_decode/RegisterFile/n1994 , \unit_decode/RegisterFile/n1995 ,
         \unit_decode/RegisterFile/n1996 , \unit_decode/RegisterFile/n1997 ,
         \unit_decode/RegisterFile/n1998 , \unit_decode/RegisterFile/n1999 ,
         \unit_decode/RegisterFile/n2000 , \unit_decode/RegisterFile/n2001 ,
         \unit_decode/RegisterFile/n2002 , \unit_decode/RegisterFile/n2003 ,
         \unit_decode/RegisterFile/n2004 , \unit_decode/RegisterFile/n2005 ,
         \unit_decode/RegisterFile/n2006 , \unit_decode/RegisterFile/n2007 ,
         \unit_decode/RegisterFile/n2008 , \unit_decode/RegisterFile/n2009 ,
         \unit_decode/RegisterFile/n2010 , \unit_decode/RegisterFile/n2011 ,
         \unit_decode/RegisterFile/n2012 , \unit_decode/RegisterFile/n2013 ,
         \unit_decode/RegisterFile/n2014 , \unit_decode/RegisterFile/n2015 ,
         \unit_decode/RegisterFile/n2016 , \unit_decode/RegisterFile/n2017 ,
         \unit_decode/RegisterFile/n2018 , \unit_decode/RegisterFile/n2019 ,
         \unit_decode/RegisterFile/n2020 , \unit_decode/RegisterFile/n2021 ,
         \unit_decode/RegisterFile/n2022 , \unit_decode/RegisterFile/n2023 ,
         \unit_decode/RegisterFile/n2024 , \unit_decode/RegisterFile/n2025 ,
         \unit_decode/RegisterFile/n2026 , \unit_decode/RegisterFile/n2027 ,
         \unit_decode/RegisterFile/n2028 , \unit_decode/RegisterFile/n2029 ,
         \unit_decode/RegisterFile/n2030 , \unit_decode/RegisterFile/n2031 ,
         \unit_decode/RegisterFile/n2032 , \unit_decode/RegisterFile/n2033 ,
         \unit_decode/RegisterFile/n2034 , \unit_decode/RegisterFile/n2035 ,
         \unit_decode/RegisterFile/n2036 , \unit_decode/RegisterFile/n2037 ,
         \unit_decode/RegisterFile/n2038 , \unit_decode/RegisterFile/n2039 ,
         \unit_decode/RegisterFile/n2040 , \unit_decode/RegisterFile/n2041 ,
         \unit_decode/RegisterFile/n2042 , \unit_decode/RegisterFile/n2043 ,
         \unit_decode/RegisterFile/n2044 , \unit_decode/RegisterFile/n2045 ,
         \unit_decode/RegisterFile/n2046 , \unit_decode/RegisterFile/n2047 ,
         \unit_decode/RegisterFile/n2048 , \unit_decode/RegisterFile/n2049 ,
         \unit_decode/RegisterFile/n2050 , \unit_decode/RegisterFile/n2051 ,
         \unit_decode/RegisterFile/n2052 , \unit_decode/RegisterFile/n2053 ,
         \unit_decode/RegisterFile/n2054 , \unit_decode/RegisterFile/n2055 ,
         \unit_decode/RegisterFile/n2056 , \unit_decode/RegisterFile/n2057 ,
         \unit_decode/RegisterFile/n2058 , \unit_decode/RegisterFile/n2059 ,
         \unit_decode/RegisterFile/n2060 , \unit_decode/RegisterFile/n2061 ,
         \unit_decode/RegisterFile/n2062 , \unit_decode/RegisterFile/n2063 ,
         \unit_decode/RegisterFile/n2064 , \unit_decode/RegisterFile/n2065 ,
         \unit_decode/RegisterFile/n2066 , \unit_decode/RegisterFile/n2067 ,
         \unit_decode/RegisterFile/n2068 , \unit_decode/RegisterFile/n2069 ,
         \unit_decode/RegisterFile/n2070 , \unit_decode/RegisterFile/n2071 ,
         \unit_decode/RegisterFile/n2072 , \unit_decode/RegisterFile/n2073 ,
         \unit_decode/RegisterFile/n2074 , \unit_decode/RegisterFile/n2075 ,
         \unit_decode/RegisterFile/n2076 , \unit_decode/RegisterFile/n2077 ,
         \unit_decode/RegisterFile/n2078 , \unit_decode/RegisterFile/n2079 ,
         \unit_decode/RegisterFile/n2080 , \unit_decode/RegisterFile/n2081 ,
         \unit_decode/RegisterFile/n2082 , \unit_decode/RegisterFile/n2083 ,
         \unit_decode/RegisterFile/n2084 , \unit_decode/RegisterFile/n2085 ,
         \unit_decode/RegisterFile/n2086 , \unit_decode/RegisterFile/n2087 ,
         \unit_decode/RegisterFile/n2088 , \unit_decode/RegisterFile/n2089 ,
         \unit_decode/RegisterFile/n2090 , \unit_decode/RegisterFile/n2091 ,
         \unit_decode/RegisterFile/n2092 , \unit_decode/RegisterFile/n2093 ,
         \unit_decode/RegisterFile/n2094 , \unit_decode/RegisterFile/n2095 ,
         \unit_decode/RegisterFile/n2096 , \unit_decode/RegisterFile/n2097 ,
         \unit_decode/RegisterFile/n2098 , \unit_decode/RegisterFile/n2099 ,
         \unit_decode/RegisterFile/n2100 , \unit_decode/RegisterFile/n2101 ,
         \unit_decode/RegisterFile/n2102 , \unit_decode/RegisterFile/n2103 ,
         \unit_decode/RegisterFile/n2104 , \unit_decode/RegisterFile/n2105 ,
         \unit_decode/RegisterFile/n2106 , \unit_decode/RegisterFile/n2107 ,
         \unit_decode/RegisterFile/n2108 , \unit_decode/RegisterFile/n2109 ,
         \unit_decode/RegisterFile/n2110 , \unit_decode/RegisterFile/n2111 ,
         \unit_decode/RegisterFile/n2112 , \unit_decode/RegisterFile/n2113 ,
         \unit_decode/RegisterFile/n2114 , \unit_decode/RegisterFile/n2115 ,
         \unit_decode/RegisterFile/n2116 , \unit_decode/RegisterFile/n2117 ,
         \unit_decode/RegisterFile/n2118 , \unit_decode/RegisterFile/n2119 ,
         \unit_decode/RegisterFile/n2120 , \unit_decode/RegisterFile/n2121 ,
         \unit_decode/RegisterFile/n2122 , \unit_decode/RegisterFile/n2123 ,
         \unit_decode/RegisterFile/n2124 , \unit_decode/RegisterFile/n2125 ,
         \unit_decode/RegisterFile/n2126 , \unit_decode/RegisterFile/n2127 ,
         \unit_decode/RegisterFile/n2128 , \unit_decode/RegisterFile/n2129 ,
         \unit_decode/RegisterFile/n2130 , \unit_decode/RegisterFile/n2131 ,
         \unit_decode/RegisterFile/n2132 , \unit_decode/RegisterFile/n2133 ,
         \unit_decode/RegisterFile/n2134 , \unit_decode/RegisterFile/n2135 ,
         \unit_decode/RegisterFile/n2136 , \unit_decode/RegisterFile/n2137 ,
         \unit_decode/RegisterFile/n2138 , \unit_decode/RegisterFile/n2139 ,
         \unit_decode/RegisterFile/n2140 , \unit_decode/RegisterFile/n2141 ,
         \unit_decode/RegisterFile/n2142 , \unit_decode/RegisterFile/n2143 ,
         \unit_decode/RegisterFile/n2144 , \unit_decode/RegisterFile/n2145 ,
         \unit_decode/RegisterFile/n2146 , \unit_decode/RegisterFile/n2147 ,
         \unit_decode/RegisterFile/n2148 , \unit_decode/RegisterFile/n2149 ,
         \unit_decode/RegisterFile/n2150 , \unit_decode/RegisterFile/n2151 ,
         \unit_decode/RegisterFile/n2152 , \unit_decode/RegisterFile/n2153 ,
         \unit_decode/RegisterFile/n2154 , \unit_decode/RegisterFile/n2155 ,
         \unit_decode/RegisterFile/n2156 , \unit_decode/RegisterFile/n2157 ,
         \unit_decode/RegisterFile/n2158 , \unit_decode/RegisterFile/n2159 ,
         \unit_decode/RegisterFile/n2160 , \unit_decode/RegisterFile/n2161 ,
         \unit_decode/RegisterFile/n2162 , \unit_decode/RegisterFile/n2163 ,
         \unit_decode/RegisterFile/n4 , \unit_decode/RegisterFile/n5 ,
         \unit_decode/RegisterFile/n6 , \unit_decode/RegisterFile/n7 ,
         \unit_decode/RegisterFile/n8 , \unit_decode/RegisterFile/n9 ,
         \unit_decode/RegisterFile/n36 , \unit_decode/RegisterFile/n37 ,
         \unit_decode/RegisterFile/n38 , \unit_decode/RegisterFile/n39 ,
         \unit_decode/RegisterFile/n40 , \unit_decode/RegisterFile/n41 ,
         \unit_decode/RegisterFile/n42 , \unit_decode/RegisterFile/n43 ,
         \unit_decode/RegisterFile/n44 , \unit_decode/RegisterFile/n45 ,
         \unit_decode/RegisterFile/n46 , \unit_decode/RegisterFile/n47 ,
         \unit_decode/RegisterFile/n48 , \unit_decode/RegisterFile/n49 ,
         \unit_decode/RegisterFile/n50 , \unit_decode/RegisterFile/n51 ,
         \unit_decode/RegisterFile/n52 , \unit_decode/RegisterFile/n53 ,
         \unit_decode/RegisterFile/n54 , \unit_decode/RegisterFile/n55 ,
         \unit_decode/RegisterFile/n56 , \unit_decode/RegisterFile/n57 ,
         \unit_decode/RegisterFile/n58 , \unit_decode/RegisterFile/n59 ,
         \unit_decode/RegisterFile/n60 , \unit_decode/RegisterFile/n61 ,
         \unit_decode/RegisterFile/n62 , \unit_decode/RegisterFile/n63 ,
         \unit_decode/RegisterFile/n64 , \unit_decode/RegisterFile/n449 ,
         \unit_decode/RegisterFile/n450 , \unit_decode/RegisterFile/n451 ,
         \unit_decode/RegisterFile/n452 , \unit_decode/RegisterFile/n453 ,
         \unit_decode/RegisterFile/n454 , \unit_decode/RegisterFile/n455 ,
         \unit_decode/RegisterFile/n456 , \unit_decode/RegisterFile/n505 ,
         \unit_decode/RegisterFile/n506 , \unit_decode/RegisterFile/n507 ,
         \unit_decode/RegisterFile/n508 , \unit_decode/RegisterFile/n509 ,
         \unit_decode/RegisterFile/n510 , \unit_decode/RegisterFile/n511 ,
         \unit_decode/RegisterFile/n512 , \unit_decode/RegisterFile/n3484 ,
         \unit_decode/RegisterFile/n3485 , \unit_decode/RegisterFile/n3486 ,
         \unit_decode/RegisterFile/n3493 , \unit_decode/RegisterFile/n3494 ,
         \unit_decode/RegisterFile/n3495 , \unit_decode/RegisterFile/n3496 ,
         \unit_decode/RegisterFile/n3497 , \unit_decode/RegisterFile/n3498 ,
         \unit_decode/RegisterFile/n3499 , \unit_decode/RegisterFile/n3500 ,
         \unit_decode/RegisterFile/n3501 , \unit_decode/RegisterFile/n3502 ,
         \unit_decode/RegisterFile/n3503 , \unit_decode/RegisterFile/n3504 ,
         \unit_decode/RegisterFile/n3505 , \unit_decode/RegisterFile/n3506 ,
         \unit_decode/RegisterFile/n3507 , \unit_decode/RegisterFile/n3508 ,
         \unit_decode/RegisterFile/n3509 , \unit_decode/RegisterFile/n3510 ,
         \unit_decode/RegisterFile/n3511 , \unit_decode/RegisterFile/n3512 ,
         \unit_decode/RegisterFile/n3513 , \unit_decode/RegisterFile/n3514 ,
         \unit_decode/RegisterFile/n3515 , \unit_decode/RegisterFile/n3516 ,
         \unit_decode/RegisterFile/n3517 , \unit_decode/RegisterFile/n3518 ,
         \unit_decode/RegisterFile/n3583 , \unit_decode/RegisterFile/n3584 ,
         \unit_decode/RegisterFile/n3585 , \unit_decode/RegisterFile/n3586 ,
         \unit_decode/RegisterFile/n3587 , \unit_decode/RegisterFile/n3588 ,
         \unit_decode/RegisterFile/n3589 , \unit_decode/RegisterFile/n3590 ,
         \unit_decode/RegisterFile/n3591 , \unit_decode/RegisterFile/n3592 ,
         \unit_decode/RegisterFile/n3593 , \unit_decode/RegisterFile/n3594 ,
         \unit_decode/RegisterFile/n3595 , \unit_decode/RegisterFile/n3596 ,
         \unit_decode/RegisterFile/n3597 , \unit_decode/RegisterFile/n3598 ,
         \unit_decode/RegisterFile/n3599 , \unit_decode/RegisterFile/n3600 ,
         \unit_decode/RegisterFile/n3601 , \unit_decode/RegisterFile/n3602 ,
         \unit_decode/RegisterFile/n3603 , \unit_decode/RegisterFile/n3604 ,
         \unit_decode/RegisterFile/n3605 , \unit_decode/RegisterFile/n3606 ,
         \unit_decode/RegisterFile/n3607 , \unit_decode/RegisterFile/n3608 ,
         \unit_decode/RegisterFile/n3609 , \unit_decode/RegisterFile/n3610 ,
         \unit_decode/RegisterFile/n3611 , \unit_decode/RegisterFile/n3612 ,
         \unit_decode/RegisterFile/n3613 , \unit_decode/RegisterFile/n3614 ,
         \unit_decode/RegisterFile/n3615 , \unit_decode/RegisterFile/n3616 ,
         \unit_decode/RegisterFile/n3617 , \unit_decode/RegisterFile/n3618 ,
         \unit_decode/RegisterFile/n3619 , \unit_decode/RegisterFile/n3620 ,
         \unit_decode/RegisterFile/n3621 , \unit_decode/RegisterFile/n3622 ,
         \unit_decode/RegisterFile/n3623 , \unit_decode/RegisterFile/n3624 ,
         \unit_decode/RegisterFile/n3625 , \unit_decode/RegisterFile/n3626 ,
         \unit_decode/RegisterFile/n3627 , \unit_decode/RegisterFile/n3628 ,
         \unit_decode/RegisterFile/n3629 , \unit_decode/RegisterFile/n3630 ,
         \unit_decode/RegisterFile/n3631 , \unit_decode/RegisterFile/n3632 ,
         \unit_decode/RegisterFile/n3633 , \unit_decode/RegisterFile/n3634 ,
         \unit_decode/RegisterFile/n3635 , \unit_decode/RegisterFile/n3636 ,
         \unit_decode/RegisterFile/n3637 , \unit_decode/RegisterFile/n3638 ,
         \unit_decode/RegisterFile/n3639 , \unit_decode/RegisterFile/n3640 ,
         \unit_decode/RegisterFile/n3641 , \unit_decode/RegisterFile/n3642 ,
         \unit_decode/RegisterFile/n3643 , \unit_decode/RegisterFile/n3644 ,
         \unit_decode/RegisterFile/n3645 , \unit_decode/RegisterFile/n3646 ,
         \unit_decode/RegisterFile/n3647 , \unit_decode/RegisterFile/n3648 ,
         \unit_decode/RegisterFile/n3649 , \unit_decode/RegisterFile/n3650 ,
         \unit_decode/RegisterFile/n3651 , \unit_decode/RegisterFile/n3652 ,
         \unit_decode/RegisterFile/n3653 , \unit_decode/RegisterFile/n3654 ,
         \unit_decode/RegisterFile/n3655 , \unit_decode/RegisterFile/n3656 ,
         \unit_decode/RegisterFile/n3657 , \unit_decode/RegisterFile/n3658 ,
         \unit_decode/RegisterFile/n3659 , \unit_decode/RegisterFile/n3660 ,
         \unit_decode/RegisterFile/n3661 , \unit_decode/RegisterFile/n3662 ,
         \unit_decode/RegisterFile/n3663 , \unit_decode/RegisterFile/n3664 ,
         \unit_decode/RegisterFile/n3665 , \unit_decode/RegisterFile/n3666 ,
         \unit_decode/RegisterFile/n3667 , \unit_decode/RegisterFile/n3668 ,
         \unit_decode/RegisterFile/n3669 , \unit_decode/RegisterFile/n3670 ,
         \unit_decode/RegisterFile/n3671 , \unit_decode/RegisterFile/n3672 ,
         \unit_decode/RegisterFile/n3673 , \unit_decode/RegisterFile/n3674 ,
         \unit_decode/RegisterFile/n3675 , \unit_decode/RegisterFile/n3676 ,
         \unit_decode/RegisterFile/n3677 , \unit_decode/RegisterFile/n3678 ,
         \unit_decode/RegisterFile/n3679 , \unit_decode/RegisterFile/n3680 ,
         \unit_decode/RegisterFile/n3681 , \unit_decode/RegisterFile/n3682 ,
         \unit_decode/RegisterFile/n3683 , \unit_decode/RegisterFile/n3684 ,
         \unit_decode/RegisterFile/n3685 , \unit_decode/RegisterFile/n3686 ,
         \unit_decode/RegisterFile/n3687 , \unit_decode/RegisterFile/n3688 ,
         \unit_decode/RegisterFile/n3689 , \unit_decode/RegisterFile/n3690 ,
         \unit_decode/RegisterFile/n3691 , \unit_decode/RegisterFile/n3692 ,
         \unit_decode/RegisterFile/n3693 , \unit_decode/RegisterFile/n3694 ,
         \unit_decode/RegisterFile/n3695 , \unit_decode/RegisterFile/n3696 ,
         \unit_decode/RegisterFile/n3697 , \unit_decode/RegisterFile/n3698 ,
         \unit_decode/RegisterFile/n3699 , \unit_decode/RegisterFile/n3700 ,
         \unit_decode/RegisterFile/n3701 , \unit_decode/RegisterFile/n3702 ,
         \unit_decode/RegisterFile/n3703 , \unit_decode/RegisterFile/n3704 ,
         \unit_decode/RegisterFile/n3705 , \unit_decode/RegisterFile/n3706 ,
         \unit_decode/RegisterFile/n3707 , \unit_decode/RegisterFile/n3708 ,
         \unit_decode/RegisterFile/n3709 , \unit_decode/RegisterFile/n3710 ,
         \unit_decode/RegisterFile/n3711 , \unit_decode/RegisterFile/n3712 ,
         \unit_decode/RegisterFile/n3713 , \unit_decode/RegisterFile/n3714 ,
         \unit_decode/RegisterFile/n3715 , \unit_decode/RegisterFile/n3716 ,
         \unit_decode/RegisterFile/n3717 , \unit_decode/RegisterFile/n3718 ,
         \unit_decode/RegisterFile/n3719 , \unit_decode/RegisterFile/n3720 ,
         \unit_decode/RegisterFile/n3721 , \unit_decode/RegisterFile/n3722 ,
         \unit_decode/RegisterFile/n3723 , \unit_decode/RegisterFile/n3724 ,
         \unit_decode/RegisterFile/n3725 , \unit_decode/RegisterFile/n3726 ,
         \unit_decode/RegisterFile/n3727 , \unit_decode/RegisterFile/n3728 ,
         \unit_decode/RegisterFile/n3729 , \unit_decode/RegisterFile/n3730 ,
         \unit_decode/RegisterFile/n3731 , \unit_decode/RegisterFile/n3732 ,
         \unit_decode/RegisterFile/n3733 , \unit_decode/RegisterFile/n3734 ,
         \unit_decode/RegisterFile/n3735 , \unit_decode/RegisterFile/n3736 ,
         \unit_decode/RegisterFile/n3737 , \unit_decode/RegisterFile/n3738 ,
         \unit_decode/RegisterFile/n3739 , \unit_decode/RegisterFile/n3740 ,
         \unit_decode/RegisterFile/n3741 , \unit_decode/RegisterFile/n3742 ,
         \unit_decode/RegisterFile/n3743 , \unit_decode/RegisterFile/n3744 ,
         \unit_decode/RegisterFile/n3745 , \unit_decode/RegisterFile/n3746 ,
         \unit_decode/RegisterFile/n3747 , \unit_decode/RegisterFile/n3772 ,
         \unit_decode/RegisterFile/n3773 , \unit_decode/RegisterFile/n3774 ,
         \unit_decode/RegisterFile/n3775 , \unit_decode/RegisterFile/n3776 ,
         \unit_decode/RegisterFile/n3777 , \unit_decode/RegisterFile/n3778 ,
         \unit_decode/RegisterFile/n3779 , \unit_decode/RegisterFile/n3804 ,
         \unit_decode/RegisterFile/n3805 , \unit_decode/RegisterFile/n3806 ,
         \unit_decode/RegisterFile/n3807 , \unit_decode/RegisterFile/n3808 ,
         \unit_decode/RegisterFile/n3809 , \unit_decode/RegisterFile/n3810 ,
         \unit_decode/RegisterFile/n3811 , \unit_decode/RegisterFile/n3836 ,
         \unit_decode/RegisterFile/n3837 , \unit_decode/RegisterFile/n3838 ,
         \unit_decode/RegisterFile/n3839 , \unit_decode/RegisterFile/n3840 ,
         \unit_decode/RegisterFile/n3841 , \unit_decode/RegisterFile/n3842 ,
         \unit_decode/RegisterFile/n3843 , \unit_decode/RegisterFile/n3868 ,
         \unit_decode/RegisterFile/n3869 , \unit_decode/RegisterFile/n3870 ,
         \unit_decode/registerB[31] , \unit_decode/registerB[30] ,
         \unit_decode/registerB[29] , \unit_decode/registerB[28] ,
         \unit_decode/registerB[27] , \unit_decode/registerB[26] ,
         \unit_decode/registerB[25] , \unit_decode/registerB[24] ,
         \unit_decode/registerB[23] , \unit_decode/registerB[22] ,
         \unit_decode/registerB[21] , \unit_decode/registerB[20] ,
         \unit_decode/registerB[19] , \unit_decode/registerB[18] ,
         \unit_decode/registerB[17] , \unit_decode/registerB[16] ,
         \unit_decode/registerB[15] , \unit_decode/registerB[14] ,
         \unit_decode/registerB[13] , \unit_decode/registerB[12] ,
         \unit_decode/registerB[11] , \unit_decode/registerB[10] ,
         \unit_decode/registerB[9] , \unit_decode/registerB[8] ,
         \unit_decode/registerB[7] , \unit_decode/registerB[6] ,
         \unit_decode/registerB[5] , \unit_decode/registerB[4] ,
         \unit_decode/registerB[3] , \unit_decode/registerB[2] ,
         \unit_decode/registerB[1] , \unit_decode/registerB[0] ,
         \unit_decode/registerA[31] , \unit_decode/registerA[30] ,
         \unit_decode/registerA[29] , \unit_decode/registerA[28] ,
         \unit_decode/registerA[27] , \unit_decode/registerA[26] ,
         \unit_decode/registerA[25] , \unit_decode/registerA[24] ,
         \unit_decode/registerA[23] , \unit_decode/registerA[22] ,
         \unit_decode/registerA[21] , \unit_decode/registerA[20] ,
         \unit_decode/registerA[19] , \unit_decode/registerA[18] ,
         \unit_decode/registerA[17] , \unit_decode/registerA[16] ,
         \unit_decode/registerA[15] , \unit_decode/registerA[14] ,
         \unit_decode/registerA[13] , \unit_decode/registerA[12] ,
         \unit_decode/registerA[11] , \unit_decode/registerA[10] ,
         \unit_decode/registerA[9] , \unit_decode/registerA[8] ,
         \unit_decode/registerA[7] , \unit_decode/registerA[6] ,
         \unit_decode/registerA[5] , \unit_decode/registerA[4] ,
         \unit_decode/registerA[3] , \unit_decode/registerA[2] ,
         \unit_decode/registerA[1] , \unit_decode/registerA[0] ,
         \unit_memory/wb_prime[31] , \unit_memory/wb_prime[30] ,
         \unit_memory/wb_prime[29] , \unit_memory/wb_prime[28] ,
         \unit_memory/wb_prime[27] , \unit_memory/wb_prime[26] ,
         \unit_memory/wb_prime[25] , \unit_memory/wb_prime[24] ,
         \unit_memory/wb_prime[23] , \unit_memory/wb_prime[22] ,
         \unit_memory/wb_prime[21] , \unit_memory/wb_prime[20] ,
         \unit_memory/wb_prime[19] , \unit_memory/wb_prime[18] ,
         \unit_memory/wb_prime[17] , \unit_memory/wb_prime[16] ,
         \unit_memory/wb_prime[15] , \unit_memory/wb_prime[14] ,
         \unit_memory/wb_prime[13] , \unit_memory/wb_prime[12] ,
         \unit_memory/wb_prime[11] , \unit_memory/wb_prime[10] ,
         \unit_memory/wb_prime[9] , \unit_memory/wb_prime[8] ,
         \unit_memory/wb_prime[7] , \unit_memory/wb_prime[6] ,
         \unit_memory/wb_prime[5] , \unit_memory/wb_prime[4] ,
         \unit_memory/wb_prime[3] , \unit_memory/wb_prime[2] ,
         \unit_memory/wb_prime[1] , \unit_memory/wb_prime[0] ,
         \unit_memory/DataMemOut[31] , \unit_memory/DataMemOut[30] ,
         \unit_memory/DataMemOut[29] , \unit_memory/DataMemOut[28] ,
         \unit_memory/DataMemOut[27] , \unit_memory/DataMemOut[26] ,
         \unit_memory/DataMemOut[25] , \unit_memory/DataMemOut[24] ,
         \unit_memory/DataMemOut[23] , \unit_memory/DataMemOut[22] ,
         \unit_memory/DataMemOut[21] , \unit_memory/DataMemOut[20] ,
         \unit_memory/DataMemOut[19] , \unit_memory/DataMemOut[18] ,
         \unit_memory/DataMemOut[17] , \unit_memory/DataMemOut[16] ,
         \unit_memory/DataMemOut[15] , \unit_memory/DataMemOut[14] ,
         \unit_memory/DataMemOut[13] , \unit_memory/DataMemOut[12] ,
         \unit_memory/DataMemOut[11] , \unit_memory/DataMemOut[10] ,
         \unit_memory/DataMemOut[9] , \unit_memory/DataMemOut[8] ,
         \unit_memory/DataMemOut[7] , \unit_memory/DataMemOut[6] ,
         \unit_memory/DataMemOut[5] , \unit_memory/DataMemOut[4] ,
         \unit_memory/DataMemOut[3] , \unit_memory/DataMemOut[2] ,
         \unit_memory/DataMemOut[1] , \unit_memory/DataMemOut[0] ,
         \unit_memory/DRAM/n3398 , \unit_memory/DRAM/n3397 ,
         \unit_memory/DRAM/n3396 , \unit_memory/DRAM/n3395 ,
         \unit_memory/DRAM/n3394 , \unit_memory/DRAM/n3393 ,
         \unit_memory/DRAM/n3392 , \unit_memory/DRAM/n3391 ,
         \unit_memory/DRAM/n3390 , \unit_memory/DRAM/n3389 ,
         \unit_memory/DRAM/n3388 , \unit_memory/DRAM/n3387 ,
         \unit_memory/DRAM/n3386 , \unit_memory/DRAM/n3385 ,
         \unit_memory/DRAM/n3384 , \unit_memory/DRAM/n3383 ,
         \unit_memory/DRAM/n3382 , \unit_memory/DRAM/n3381 ,
         \unit_memory/DRAM/n3380 , \unit_memory/DRAM/n3379 ,
         \unit_memory/DRAM/n3378 , \unit_memory/DRAM/n3377 ,
         \unit_memory/DRAM/n3376 , \unit_memory/DRAM/n3375 ,
         \unit_memory/DRAM/n3374 , \unit_memory/DRAM/n3373 ,
         \unit_memory/DRAM/n3372 , \unit_memory/DRAM/n3371 ,
         \unit_memory/DRAM/n3370 , \unit_memory/DRAM/n3369 ,
         \unit_memory/DRAM/n3368 , \unit_memory/DRAM/n3367 ,
         \unit_memory/DRAM/n3366 , \unit_memory/DRAM/n3365 ,
         \unit_memory/DRAM/n3364 , \unit_memory/DRAM/n3363 ,
         \unit_memory/DRAM/n3362 , \unit_memory/DRAM/n3361 ,
         \unit_memory/DRAM/n3360 , \unit_memory/DRAM/n3359 ,
         \unit_memory/DRAM/n3358 , \unit_memory/DRAM/n3357 ,
         \unit_memory/DRAM/n3356 , \unit_memory/DRAM/n3355 ,
         \unit_memory/DRAM/n3354 , \unit_memory/DRAM/n3353 ,
         \unit_memory/DRAM/n3352 , \unit_memory/DRAM/n3351 ,
         \unit_memory/DRAM/n3350 , \unit_memory/DRAM/n3349 ,
         \unit_memory/DRAM/n3348 , \unit_memory/DRAM/n3347 ,
         \unit_memory/DRAM/n3346 , \unit_memory/DRAM/n3345 ,
         \unit_memory/DRAM/n3344 , \unit_memory/DRAM/n3343 ,
         \unit_memory/DRAM/n3342 , \unit_memory/DRAM/n3341 ,
         \unit_memory/DRAM/n3340 , \unit_memory/DRAM/n3339 ,
         \unit_memory/DRAM/n3338 , \unit_memory/DRAM/n3337 ,
         \unit_memory/DRAM/n3336 , \unit_memory/DRAM/n3335 ,
         \unit_memory/DRAM/n3334 , \unit_memory/DRAM/n3333 ,
         \unit_memory/DRAM/n3332 , \unit_memory/DRAM/n3331 ,
         \unit_memory/DRAM/n3330 , \unit_memory/DRAM/n3329 ,
         \unit_memory/DRAM/n3328 , \unit_memory/DRAM/n3327 ,
         \unit_memory/DRAM/n3326 , \unit_memory/DRAM/n3325 ,
         \unit_memory/DRAM/n3324 , \unit_memory/DRAM/n3323 ,
         \unit_memory/DRAM/n3322 , \unit_memory/DRAM/n3321 ,
         \unit_memory/DRAM/n3320 , \unit_memory/DRAM/n3319 ,
         \unit_memory/DRAM/n3318 , \unit_memory/DRAM/n3317 ,
         \unit_memory/DRAM/n3316 , \unit_memory/DRAM/n3315 ,
         \unit_memory/DRAM/n3314 , \unit_memory/DRAM/n3313 ,
         \unit_memory/DRAM/n3312 , \unit_memory/DRAM/n3311 ,
         \unit_memory/DRAM/n3310 , \unit_memory/DRAM/n3309 ,
         \unit_memory/DRAM/n3308 , \unit_memory/DRAM/n3307 ,
         \unit_memory/DRAM/n3306 , \unit_memory/DRAM/n3305 ,
         \unit_memory/DRAM/n3304 , \unit_memory/DRAM/n3303 ,
         \unit_memory/DRAM/n3302 , \unit_memory/DRAM/n3301 ,
         \unit_memory/DRAM/n3300 , \unit_memory/DRAM/n3299 ,
         \unit_memory/DRAM/n3298 , \unit_memory/DRAM/n3297 ,
         \unit_memory/DRAM/n3296 , \unit_memory/DRAM/n3295 ,
         \unit_memory/DRAM/n3294 , \unit_memory/DRAM/n3293 ,
         \unit_memory/DRAM/n3292 , \unit_memory/DRAM/n3291 ,
         \unit_memory/DRAM/n3290 , \unit_memory/DRAM/n3289 ,
         \unit_memory/DRAM/n3288 , \unit_memory/DRAM/n3287 ,
         \unit_memory/DRAM/n3286 , \unit_memory/DRAM/n3285 ,
         \unit_memory/DRAM/n3284 , \unit_memory/DRAM/n3283 ,
         \unit_memory/DRAM/n3282 , \unit_memory/DRAM/n3281 ,
         \unit_memory/DRAM/n3280 , \unit_memory/DRAM/n3279 ,
         \unit_memory/DRAM/n3278 , \unit_memory/DRAM/n3277 ,
         \unit_memory/DRAM/n3276 , \unit_memory/DRAM/n3275 ,
         \unit_memory/DRAM/n3274 , \unit_memory/DRAM/n3273 ,
         \unit_memory/DRAM/n3272 , \unit_memory/DRAM/n3271 ,
         \unit_memory/DRAM/n3270 , \unit_memory/DRAM/n3269 ,
         \unit_memory/DRAM/n3268 , \unit_memory/DRAM/n3267 ,
         \unit_memory/DRAM/n3266 , \unit_memory/DRAM/n3265 ,
         \unit_memory/DRAM/n3264 , \unit_memory/DRAM/n3263 ,
         \unit_memory/DRAM/n3262 , \unit_memory/DRAM/n3261 ,
         \unit_memory/DRAM/n3260 , \unit_memory/DRAM/n3259 ,
         \unit_memory/DRAM/n3258 , \unit_memory/DRAM/n3257 ,
         \unit_memory/DRAM/n3256 , \unit_memory/DRAM/n3255 ,
         \unit_memory/DRAM/n3254 , \unit_memory/DRAM/n3253 ,
         \unit_memory/DRAM/n3252 , \unit_memory/DRAM/n3251 ,
         \unit_memory/DRAM/n3250 , \unit_memory/DRAM/n3249 ,
         \unit_memory/DRAM/n3248 , \unit_memory/DRAM/n3247 ,
         \unit_memory/DRAM/n3246 , \unit_memory/DRAM/n3245 ,
         \unit_memory/DRAM/n3244 , \unit_memory/DRAM/n3243 ,
         \unit_memory/DRAM/n3242 , \unit_memory/DRAM/n3241 ,
         \unit_memory/DRAM/n3240 , \unit_memory/DRAM/n3239 ,
         \unit_memory/DRAM/n3238 , \unit_memory/DRAM/n3237 ,
         \unit_memory/DRAM/n3236 , \unit_memory/DRAM/n3235 ,
         \unit_memory/DRAM/n3234 , \unit_memory/DRAM/n3233 ,
         \unit_memory/DRAM/n3232 , \unit_memory/DRAM/n3231 ,
         \unit_memory/DRAM/n3230 , \unit_memory/DRAM/n3229 ,
         \unit_memory/DRAM/n3228 , \unit_memory/DRAM/n3227 ,
         \unit_memory/DRAM/n3226 , \unit_memory/DRAM/n3225 ,
         \unit_memory/DRAM/n3224 , \unit_memory/DRAM/n3223 ,
         \unit_memory/DRAM/n3222 , \unit_memory/DRAM/n3221 ,
         \unit_memory/DRAM/n3220 , \unit_memory/DRAM/n3219 ,
         \unit_memory/DRAM/n3218 , \unit_memory/DRAM/n3217 ,
         \unit_memory/DRAM/n3216 , \unit_memory/DRAM/n3215 ,
         \unit_memory/DRAM/n3214 , \unit_memory/DRAM/n3213 ,
         \unit_memory/DRAM/n3212 , \unit_memory/DRAM/n3211 ,
         \unit_memory/DRAM/n3210 , \unit_memory/DRAM/n3209 ,
         \unit_memory/DRAM/n3208 , \unit_memory/DRAM/n3207 ,
         \unit_memory/DRAM/n3206 , \unit_memory/DRAM/n3205 ,
         \unit_memory/DRAM/n3204 , \unit_memory/DRAM/n3203 ,
         \unit_memory/DRAM/n3202 , \unit_memory/DRAM/n3201 ,
         \unit_memory/DRAM/n3200 , \unit_memory/DRAM/n3199 ,
         \unit_memory/DRAM/n3198 , \unit_memory/DRAM/n3197 ,
         \unit_memory/DRAM/n3196 , \unit_memory/DRAM/n3195 ,
         \unit_memory/DRAM/n3194 , \unit_memory/DRAM/n3193 ,
         \unit_memory/DRAM/n3192 , \unit_memory/DRAM/n3191 ,
         \unit_memory/DRAM/n3190 , \unit_memory/DRAM/n3189 ,
         \unit_memory/DRAM/n3188 , \unit_memory/DRAM/n3187 ,
         \unit_memory/DRAM/n3186 , \unit_memory/DRAM/n3185 ,
         \unit_memory/DRAM/n3184 , \unit_memory/DRAM/n3183 ,
         \unit_memory/DRAM/n3182 , \unit_memory/DRAM/n3181 ,
         \unit_memory/DRAM/n3180 , \unit_memory/DRAM/n3179 ,
         \unit_memory/DRAM/n3178 , \unit_memory/DRAM/n3177 ,
         \unit_memory/DRAM/n3176 , \unit_memory/DRAM/n3175 ,
         \unit_memory/DRAM/n3174 , \unit_memory/DRAM/n3173 ,
         \unit_memory/DRAM/n3172 , \unit_memory/DRAM/n3171 ,
         \unit_memory/DRAM/n3170 , \unit_memory/DRAM/n3169 ,
         \unit_memory/DRAM/n3168 , \unit_memory/DRAM/n3167 ,
         \unit_memory/DRAM/n3166 , \unit_memory/DRAM/n3165 ,
         \unit_memory/DRAM/n3164 , \unit_memory/DRAM/n3163 ,
         \unit_memory/DRAM/n3162 , \unit_memory/DRAM/n3161 ,
         \unit_memory/DRAM/n3160 , \unit_memory/DRAM/n3159 ,
         \unit_memory/DRAM/n3158 , \unit_memory/DRAM/n3157 ,
         \unit_memory/DRAM/n3156 , \unit_memory/DRAM/n3155 ,
         \unit_memory/DRAM/n3154 , \unit_memory/DRAM/n3153 ,
         \unit_memory/DRAM/n3152 , \unit_memory/DRAM/n3151 ,
         \unit_memory/DRAM/n3150 , \unit_memory/DRAM/n3149 ,
         \unit_memory/DRAM/n3148 , \unit_memory/DRAM/n3147 ,
         \unit_memory/DRAM/n3146 , \unit_memory/DRAM/n3145 ,
         \unit_memory/DRAM/n3144 , \unit_memory/DRAM/n3143 ,
         \unit_memory/DRAM/n3142 , \unit_memory/DRAM/n3141 ,
         \unit_memory/DRAM/n3140 , \unit_memory/DRAM/n3139 ,
         \unit_memory/DRAM/n3138 , \unit_memory/DRAM/n3137 ,
         \unit_memory/DRAM/n3136 , \unit_memory/DRAM/n3135 ,
         \unit_memory/DRAM/n3134 , \unit_memory/DRAM/n3133 ,
         \unit_memory/DRAM/n3132 , \unit_memory/DRAM/n3131 ,
         \unit_memory/DRAM/n3130 , \unit_memory/DRAM/n3129 ,
         \unit_memory/DRAM/n3128 , \unit_memory/DRAM/n3127 ,
         \unit_memory/DRAM/n3126 , \unit_memory/DRAM/n3125 ,
         \unit_memory/DRAM/n3124 , \unit_memory/DRAM/n3123 ,
         \unit_memory/DRAM/n3122 , \unit_memory/DRAM/n3121 ,
         \unit_memory/DRAM/n3120 , \unit_memory/DRAM/n3119 ,
         \unit_memory/DRAM/n3118 , \unit_memory/DRAM/n3117 ,
         \unit_memory/DRAM/n3116 , \unit_memory/DRAM/n3115 ,
         \unit_memory/DRAM/n3114 , \unit_memory/DRAM/n3113 ,
         \unit_memory/DRAM/n3112 , \unit_memory/DRAM/n3111 ,
         \unit_memory/DRAM/n3110 , \unit_memory/DRAM/n3109 ,
         \unit_memory/DRAM/n3108 , \unit_memory/DRAM/n3107 ,
         \unit_memory/DRAM/n3106 , \unit_memory/DRAM/n3105 ,
         \unit_memory/DRAM/n3104 , \unit_memory/DRAM/n3103 ,
         \unit_memory/DRAM/n3102 , \unit_memory/DRAM/n3101 ,
         \unit_memory/DRAM/n3100 , \unit_memory/DRAM/n3099 ,
         \unit_memory/DRAM/n3098 , \unit_memory/DRAM/n3097 ,
         \unit_memory/DRAM/n3096 , \unit_memory/DRAM/n3095 ,
         \unit_memory/DRAM/n3094 , \unit_memory/DRAM/n3093 ,
         \unit_memory/DRAM/n3092 , \unit_memory/DRAM/n3091 ,
         \unit_memory/DRAM/n3090 , \unit_memory/DRAM/n3089 ,
         \unit_memory/DRAM/n3088 , \unit_memory/DRAM/n3087 ,
         \unit_memory/DRAM/n3086 , \unit_memory/DRAM/n3085 ,
         \unit_memory/DRAM/n3084 , \unit_memory/DRAM/n3083 ,
         \unit_memory/DRAM/n3082 , \unit_memory/DRAM/n3081 ,
         \unit_memory/DRAM/n3080 , \unit_memory/DRAM/n3079 ,
         \unit_memory/DRAM/n3078 , \unit_memory/DRAM/n3077 ,
         \unit_memory/DRAM/n3076 , \unit_memory/DRAM/n3075 ,
         \unit_memory/DRAM/n3074 , \unit_memory/DRAM/n3073 ,
         \unit_memory/DRAM/n3072 , \unit_memory/DRAM/n3071 ,
         \unit_memory/DRAM/n3070 , \unit_memory/DRAM/n3069 ,
         \unit_memory/DRAM/n3068 , \unit_memory/DRAM/n3067 ,
         \unit_memory/DRAM/n3066 , \unit_memory/DRAM/n3065 ,
         \unit_memory/DRAM/n3064 , \unit_memory/DRAM/n3063 ,
         \unit_memory/DRAM/n3062 , \unit_memory/DRAM/n3061 ,
         \unit_memory/DRAM/n3060 , \unit_memory/DRAM/n3059 ,
         \unit_memory/DRAM/n3058 , \unit_memory/DRAM/n3057 ,
         \unit_memory/DRAM/n3056 , \unit_memory/DRAM/n3055 ,
         \unit_memory/DRAM/n3054 , \unit_memory/DRAM/n3053 ,
         \unit_memory/DRAM/n3052 , \unit_memory/DRAM/n3051 ,
         \unit_memory/DRAM/n3050 , \unit_memory/DRAM/n3049 ,
         \unit_memory/DRAM/n3048 , \unit_memory/DRAM/n3047 ,
         \unit_memory/DRAM/n3046 , \unit_memory/DRAM/n3045 ,
         \unit_memory/DRAM/n3044 , \unit_memory/DRAM/n3043 ,
         \unit_memory/DRAM/n3042 , \unit_memory/DRAM/n3041 ,
         \unit_memory/DRAM/n3040 , \unit_memory/DRAM/n3039 ,
         \unit_memory/DRAM/n3038 , \unit_memory/DRAM/n3037 ,
         \unit_memory/DRAM/n3036 , \unit_memory/DRAM/n3035 ,
         \unit_memory/DRAM/n3034 , \unit_memory/DRAM/n3033 ,
         \unit_memory/DRAM/n3032 , \unit_memory/DRAM/n3031 ,
         \unit_memory/DRAM/n3030 , \unit_memory/DRAM/n3029 ,
         \unit_memory/DRAM/n3028 , \unit_memory/DRAM/n3027 ,
         \unit_memory/DRAM/n3026 , \unit_memory/DRAM/n3025 ,
         \unit_memory/DRAM/n3024 , \unit_memory/DRAM/n3023 ,
         \unit_memory/DRAM/n3022 , \unit_memory/DRAM/n3021 ,
         \unit_memory/DRAM/n3020 , \unit_memory/DRAM/n3019 ,
         \unit_memory/DRAM/n3018 , \unit_memory/DRAM/n3017 ,
         \unit_memory/DRAM/n3016 , \unit_memory/DRAM/n3015 ,
         \unit_memory/DRAM/n3014 , \unit_memory/DRAM/n3013 ,
         \unit_memory/DRAM/n3012 , \unit_memory/DRAM/n3011 ,
         \unit_memory/DRAM/n3010 , \unit_memory/DRAM/n3009 ,
         \unit_memory/DRAM/n3008 , \unit_memory/DRAM/n3007 ,
         \unit_memory/DRAM/n3006 , \unit_memory/DRAM/n3005 ,
         \unit_memory/DRAM/n3004 , \unit_memory/DRAM/n3003 ,
         \unit_memory/DRAM/n3002 , \unit_memory/DRAM/n3001 ,
         \unit_memory/DRAM/n3000 , \unit_memory/DRAM/n2999 ,
         \unit_memory/DRAM/n2998 , \unit_memory/DRAM/n2997 ,
         \unit_memory/DRAM/n2996 , \unit_memory/DRAM/n2995 ,
         \unit_memory/DRAM/n2994 , \unit_memory/DRAM/n2993 ,
         \unit_memory/DRAM/n2992 , \unit_memory/DRAM/n2991 ,
         \unit_memory/DRAM/n2990 , \unit_memory/DRAM/n2989 ,
         \unit_memory/DRAM/n2988 , \unit_memory/DRAM/n2987 ,
         \unit_memory/DRAM/n2986 , \unit_memory/DRAM/n2985 ,
         \unit_memory/DRAM/n2984 , \unit_memory/DRAM/n2983 ,
         \unit_memory/DRAM/n2982 , \unit_memory/DRAM/n2981 ,
         \unit_memory/DRAM/n2980 , \unit_memory/DRAM/n2979 ,
         \unit_memory/DRAM/n2978 , \unit_memory/DRAM/n2977 ,
         \unit_memory/DRAM/n2976 , \unit_memory/DRAM/n2975 ,
         \unit_memory/DRAM/n2974 , \unit_memory/DRAM/n2973 ,
         \unit_memory/DRAM/n2972 , \unit_memory/DRAM/n2971 ,
         \unit_memory/DRAM/n2970 , \unit_memory/DRAM/n2969 ,
         \unit_memory/DRAM/n2968 , \unit_memory/DRAM/n2967 ,
         \unit_memory/DRAM/n2966 , \unit_memory/DRAM/n2965 ,
         \unit_memory/DRAM/n2964 , \unit_memory/DRAM/n2963 ,
         \unit_memory/DRAM/n2962 , \unit_memory/DRAM/n2961 ,
         \unit_memory/DRAM/n2960 , \unit_memory/DRAM/n2959 ,
         \unit_memory/DRAM/n2958 , \unit_memory/DRAM/n2957 ,
         \unit_memory/DRAM/n2956 , \unit_memory/DRAM/n2955 ,
         \unit_memory/DRAM/n2954 , \unit_memory/DRAM/n2953 ,
         \unit_memory/DRAM/n2952 , \unit_memory/DRAM/n2951 ,
         \unit_memory/DRAM/n2950 , \unit_memory/DRAM/n2949 ,
         \unit_memory/DRAM/n2948 , \unit_memory/DRAM/n2947 ,
         \unit_memory/DRAM/n2946 , \unit_memory/DRAM/n2945 ,
         \unit_memory/DRAM/n2944 , \unit_memory/DRAM/n2943 ,
         \unit_memory/DRAM/n2942 , \unit_memory/DRAM/n2941 ,
         \unit_memory/DRAM/n2940 , \unit_memory/DRAM/n2939 ,
         \unit_memory/DRAM/n2938 , \unit_memory/DRAM/n2937 ,
         \unit_memory/DRAM/n2936 , \unit_memory/DRAM/n2935 ,
         \unit_memory/DRAM/n2934 , \unit_memory/DRAM/n2933 ,
         \unit_memory/DRAM/n2932 , \unit_memory/DRAM/n2931 ,
         \unit_memory/DRAM/n2930 , \unit_memory/DRAM/n2929 ,
         \unit_memory/DRAM/n2928 , \unit_memory/DRAM/n2927 ,
         \unit_memory/DRAM/n2926 , \unit_memory/DRAM/n2925 ,
         \unit_memory/DRAM/n2924 , \unit_memory/DRAM/n2923 ,
         \unit_memory/DRAM/n2922 , \unit_memory/DRAM/n2921 ,
         \unit_memory/DRAM/n2920 , \unit_memory/DRAM/n2919 ,
         \unit_memory/DRAM/n2918 , \unit_memory/DRAM/n2917 ,
         \unit_memory/DRAM/n2916 , \unit_memory/DRAM/n2915 ,
         \unit_memory/DRAM/n2914 , \unit_memory/DRAM/n2913 ,
         \unit_memory/DRAM/n2912 , \unit_memory/DRAM/n2911 ,
         \unit_memory/DRAM/n2910 , \unit_memory/DRAM/n2909 ,
         \unit_memory/DRAM/n2908 , \unit_memory/DRAM/n2907 ,
         \unit_memory/DRAM/n2906 , \unit_memory/DRAM/n2905 ,
         \unit_memory/DRAM/n2904 , \unit_memory/DRAM/n2903 ,
         \unit_memory/DRAM/n2902 , \unit_memory/DRAM/n2901 ,
         \unit_memory/DRAM/n2900 , \unit_memory/DRAM/n2899 ,
         \unit_memory/DRAM/n2898 , \unit_memory/DRAM/n2897 ,
         \unit_memory/DRAM/n2896 , \unit_memory/DRAM/n2895 ,
         \unit_memory/DRAM/n2894 , \unit_memory/DRAM/n2893 ,
         \unit_memory/DRAM/n2892 , \unit_memory/DRAM/n2891 ,
         \unit_memory/DRAM/n2890 , \unit_memory/DRAM/n2889 ,
         \unit_memory/DRAM/n2888 , \unit_memory/DRAM/n2887 ,
         \unit_memory/DRAM/n2886 , \unit_memory/DRAM/n2885 ,
         \unit_memory/DRAM/n2884 , \unit_memory/DRAM/n2883 ,
         \unit_memory/DRAM/n2882 , \unit_memory/DRAM/n2881 ,
         \unit_memory/DRAM/n2880 , \unit_memory/DRAM/n2879 ,
         \unit_memory/DRAM/n2878 , \unit_memory/DRAM/n2877 ,
         \unit_memory/DRAM/n2876 , \unit_memory/DRAM/n2875 ,
         \unit_memory/DRAM/n2874 , \unit_memory/DRAM/n2873 ,
         \unit_memory/DRAM/n2872 , \unit_memory/DRAM/n2871 ,
         \unit_memory/DRAM/n2870 , \unit_memory/DRAM/n2869 ,
         \unit_memory/DRAM/n2868 , \unit_memory/DRAM/n2867 ,
         \unit_memory/DRAM/n2866 , \unit_memory/DRAM/n2865 ,
         \unit_memory/DRAM/n2864 , \unit_memory/DRAM/n2863 ,
         \unit_memory/DRAM/n2862 , \unit_memory/DRAM/n2861 ,
         \unit_memory/DRAM/n2860 , \unit_memory/DRAM/n2859 ,
         \unit_memory/DRAM/n2858 , \unit_memory/DRAM/n2857 ,
         \unit_memory/DRAM/n2856 , \unit_memory/DRAM/n2855 ,
         \unit_memory/DRAM/n2854 , \unit_memory/DRAM/n2853 ,
         \unit_memory/DRAM/n2852 , \unit_memory/DRAM/n2851 ,
         \unit_memory/DRAM/n2850 , \unit_memory/DRAM/n2849 ,
         \unit_memory/DRAM/n2848 , \unit_memory/DRAM/n2847 ,
         \unit_memory/DRAM/n2846 , \unit_memory/DRAM/n2845 ,
         \unit_memory/DRAM/n2844 , \unit_memory/DRAM/n2843 ,
         \unit_memory/DRAM/n2842 , \unit_memory/DRAM/n2841 ,
         \unit_memory/DRAM/n2840 , \unit_memory/DRAM/n2839 ,
         \unit_memory/DRAM/n2838 , \unit_memory/DRAM/n2837 ,
         \unit_memory/DRAM/n2836 , \unit_memory/DRAM/n2835 ,
         \unit_memory/DRAM/n2834 , \unit_memory/DRAM/n2833 ,
         \unit_memory/DRAM/n2832 , \unit_memory/DRAM/n2831 ,
         \unit_memory/DRAM/n2830 , \unit_memory/DRAM/n2829 ,
         \unit_memory/DRAM/n2828 , \unit_memory/DRAM/n2827 ,
         \unit_memory/DRAM/n2826 , \unit_memory/DRAM/n2825 ,
         \unit_memory/DRAM/n2824 , \unit_memory/DRAM/n2823 ,
         \unit_memory/DRAM/n2822 , \unit_memory/DRAM/n2821 ,
         \unit_memory/DRAM/n2820 , \unit_memory/DRAM/n2819 ,
         \unit_memory/DRAM/n2818 , \unit_memory/DRAM/n2817 ,
         \unit_memory/DRAM/n2816 , \unit_memory/DRAM/n2815 ,
         \unit_memory/DRAM/n2814 , \unit_memory/DRAM/n2813 ,
         \unit_memory/DRAM/n2812 , \unit_memory/DRAM/n2811 ,
         \unit_memory/DRAM/n2810 , \unit_memory/DRAM/n2809 ,
         \unit_memory/DRAM/n2808 , \unit_memory/DRAM/n2807 ,
         \unit_memory/DRAM/n2806 , \unit_memory/DRAM/n2805 ,
         \unit_memory/DRAM/n2804 , \unit_memory/DRAM/n2803 ,
         \unit_memory/DRAM/n2802 , \unit_memory/DRAM/n2801 ,
         \unit_memory/DRAM/n2800 , \unit_memory/DRAM/n2799 ,
         \unit_memory/DRAM/n2798 , \unit_memory/DRAM/n2797 ,
         \unit_memory/DRAM/n2796 , \unit_memory/DRAM/n2795 ,
         \unit_memory/DRAM/n2794 , \unit_memory/DRAM/n2793 ,
         \unit_memory/DRAM/n2792 , \unit_memory/DRAM/n2791 ,
         \unit_memory/DRAM/n2790 , \unit_memory/DRAM/n2789 ,
         \unit_memory/DRAM/n2788 , \unit_memory/DRAM/n2787 ,
         \unit_memory/DRAM/n2786 , \unit_memory/DRAM/n2785 ,
         \unit_memory/DRAM/n2784 , \unit_memory/DRAM/n2783 ,
         \unit_memory/DRAM/n2782 , \unit_memory/DRAM/n2781 ,
         \unit_memory/DRAM/n2780 , \unit_memory/DRAM/n2779 ,
         \unit_memory/DRAM/n2778 , \unit_memory/DRAM/n2777 ,
         \unit_memory/DRAM/n2776 , \unit_memory/DRAM/n2775 ,
         \unit_memory/DRAM/n2774 , \unit_memory/DRAM/n2773 ,
         \unit_memory/DRAM/n2772 , \unit_memory/DRAM/n2771 ,
         \unit_memory/DRAM/n2770 , \unit_memory/DRAM/n2769 ,
         \unit_memory/DRAM/n2768 , \unit_memory/DRAM/n2767 ,
         \unit_memory/DRAM/n2766 , \unit_memory/DRAM/n2765 ,
         \unit_memory/DRAM/n2764 , \unit_memory/DRAM/n2763 ,
         \unit_memory/DRAM/n2762 , \unit_memory/DRAM/n2761 ,
         \unit_memory/DRAM/n2760 , \unit_memory/DRAM/n2759 ,
         \unit_memory/DRAM/n2758 , \unit_memory/DRAM/n2757 ,
         \unit_memory/DRAM/n2756 , \unit_memory/DRAM/n2755 ,
         \unit_memory/DRAM/n2754 , \unit_memory/DRAM/n2753 ,
         \unit_memory/DRAM/n2752 , \unit_memory/DRAM/n2751 ,
         \unit_memory/DRAM/n2750 , \unit_memory/DRAM/n2749 ,
         \unit_memory/DRAM/n2748 , \unit_memory/DRAM/n2747 ,
         \unit_memory/DRAM/n2746 , \unit_memory/DRAM/n2745 ,
         \unit_memory/DRAM/n2744 , \unit_memory/DRAM/n2743 ,
         \unit_memory/DRAM/n2742 , \unit_memory/DRAM/n2741 ,
         \unit_memory/DRAM/n2740 , \unit_memory/DRAM/n2739 ,
         \unit_memory/DRAM/n2738 , \unit_memory/DRAM/n2737 ,
         \unit_memory/DRAM/n2736 , \unit_memory/DRAM/n2735 ,
         \unit_memory/DRAM/n2734 , \unit_memory/DRAM/n2733 ,
         \unit_memory/DRAM/n2732 , \unit_memory/DRAM/n2731 ,
         \unit_memory/DRAM/n2730 , \unit_memory/DRAM/n2729 ,
         \unit_memory/DRAM/n2728 , \unit_memory/DRAM/n2727 ,
         \unit_memory/DRAM/n2726 , \unit_memory/DRAM/n2725 ,
         \unit_memory/DRAM/n2724 , \unit_memory/DRAM/n2723 ,
         \unit_memory/DRAM/n2722 , \unit_memory/DRAM/n2721 ,
         \unit_memory/DRAM/n2720 , \unit_memory/DRAM/n2719 ,
         \unit_memory/DRAM/n2718 , \unit_memory/DRAM/n2717 ,
         \unit_memory/DRAM/n2716 , \unit_memory/DRAM/n2715 ,
         \unit_memory/DRAM/n2714 , \unit_memory/DRAM/n2713 ,
         \unit_memory/DRAM/n2712 , \unit_memory/DRAM/n2711 ,
         \unit_memory/DRAM/n2710 , \unit_memory/DRAM/n2709 ,
         \unit_memory/DRAM/n2708 , \unit_memory/DRAM/n2707 ,
         \unit_memory/DRAM/n2706 , \unit_memory/DRAM/n2705 ,
         \unit_memory/DRAM/n2704 , \unit_memory/DRAM/n2703 ,
         \unit_memory/DRAM/n2702 , \unit_memory/DRAM/n2701 ,
         \unit_memory/DRAM/n2700 , \unit_memory/DRAM/n2699 ,
         \unit_memory/DRAM/n2698 , \unit_memory/DRAM/n2697 ,
         \unit_memory/DRAM/n2696 , \unit_memory/DRAM/n2695 ,
         \unit_memory/DRAM/n2694 , \unit_memory/DRAM/n2693 ,
         \unit_memory/DRAM/n2692 , \unit_memory/DRAM/n2691 ,
         \unit_memory/DRAM/n2690 , \unit_memory/DRAM/n2689 ,
         \unit_memory/DRAM/n2688 , \unit_memory/DRAM/n2687 ,
         \unit_memory/DRAM/n2686 , \unit_memory/DRAM/n2685 ,
         \unit_memory/DRAM/n2684 , \unit_memory/DRAM/n2683 ,
         \unit_memory/DRAM/n2682 , \unit_memory/DRAM/n2681 ,
         \unit_memory/DRAM/n2680 , \unit_memory/DRAM/n2679 ,
         \unit_memory/DRAM/n2678 , \unit_memory/DRAM/n2677 ,
         \unit_memory/DRAM/n2676 , \unit_memory/DRAM/n2675 ,
         \unit_memory/DRAM/n2674 , \unit_memory/DRAM/n2673 ,
         \unit_memory/DRAM/n2672 , \unit_memory/DRAM/n2671 ,
         \unit_memory/DRAM/n2670 , \unit_memory/DRAM/n2669 ,
         \unit_memory/DRAM/n2668 , \unit_memory/DRAM/n2667 ,
         \unit_memory/DRAM/n2666 , \unit_memory/DRAM/n2665 ,
         \unit_memory/DRAM/n2664 , \unit_memory/DRAM/n2663 ,
         \unit_memory/DRAM/n2662 , \unit_memory/DRAM/n2661 ,
         \unit_memory/DRAM/n2660 , \unit_memory/DRAM/n2659 ,
         \unit_memory/DRAM/n2658 , \unit_memory/DRAM/n2657 ,
         \unit_memory/DRAM/n2656 , \unit_memory/DRAM/n2655 ,
         \unit_memory/DRAM/n2654 , \unit_memory/DRAM/n2653 ,
         \unit_memory/DRAM/n2652 , \unit_memory/DRAM/n2651 ,
         \unit_memory/DRAM/n2650 , \unit_memory/DRAM/n2649 ,
         \unit_memory/DRAM/n2648 , \unit_memory/DRAM/n2647 ,
         \unit_memory/DRAM/n2646 , \unit_memory/DRAM/n2645 ,
         \unit_memory/DRAM/n2644 , \unit_memory/DRAM/n2643 ,
         \unit_memory/DRAM/n2642 , \unit_memory/DRAM/n2641 ,
         \unit_memory/DRAM/n2640 , \unit_memory/DRAM/n2639 ,
         \unit_memory/DRAM/n2638 , \unit_memory/DRAM/n2637 ,
         \unit_memory/DRAM/n2636 , \unit_memory/DRAM/n2635 ,
         \unit_memory/DRAM/n2634 , \unit_memory/DRAM/n2633 ,
         \unit_memory/DRAM/n2632 , \unit_memory/DRAM/n2631 ,
         \unit_memory/DRAM/n2630 , \unit_memory/DRAM/n2629 ,
         \unit_memory/DRAM/n2628 , \unit_memory/DRAM/n2627 ,
         \unit_memory/DRAM/n2626 , \unit_memory/DRAM/n2625 ,
         \unit_memory/DRAM/n2624 , \unit_memory/DRAM/n2623 ,
         \unit_memory/DRAM/n2622 , \unit_memory/DRAM/n2621 ,
         \unit_memory/DRAM/n2620 , \unit_memory/DRAM/n2619 ,
         \unit_memory/DRAM/n2618 , \unit_memory/DRAM/n2617 ,
         \unit_memory/DRAM/n2616 , \unit_memory/DRAM/n2615 ,
         \unit_memory/DRAM/n2614 , \unit_memory/DRAM/n2613 ,
         \unit_memory/DRAM/n2612 , \unit_memory/DRAM/n2611 ,
         \unit_memory/DRAM/n2610 , \unit_memory/DRAM/n2609 ,
         \unit_memory/DRAM/n2608 , \unit_memory/DRAM/n2607 ,
         \unit_memory/DRAM/n2606 , \unit_memory/DRAM/n2605 ,
         \unit_memory/DRAM/n2604 , \unit_memory/DRAM/n2603 ,
         \unit_memory/DRAM/n2602 , \unit_memory/DRAM/n2601 ,
         \unit_memory/DRAM/n2600 , \unit_memory/DRAM/n2599 ,
         \unit_memory/DRAM/n2598 , \unit_memory/DRAM/n2597 ,
         \unit_memory/DRAM/n2596 , \unit_memory/DRAM/n2595 ,
         \unit_memory/DRAM/n2594 , \unit_memory/DRAM/n2593 ,
         \unit_memory/DRAM/n2592 , \unit_memory/DRAM/n2591 ,
         \unit_memory/DRAM/n2590 , \unit_memory/DRAM/n2589 ,
         \unit_memory/DRAM/n2588 , \unit_memory/DRAM/n2587 ,
         \unit_memory/DRAM/n2586 , \unit_memory/DRAM/n2585 ,
         \unit_memory/DRAM/n2584 , \unit_memory/DRAM/n2583 ,
         \unit_memory/DRAM/n2582 , \unit_memory/DRAM/n2581 ,
         \unit_memory/DRAM/n2580 , \unit_memory/DRAM/n2579 ,
         \unit_memory/DRAM/n2578 , \unit_memory/DRAM/n2577 ,
         \unit_memory/DRAM/n2576 , \unit_memory/DRAM/n2575 ,
         \unit_memory/DRAM/n2574 , \unit_memory/DRAM/n2573 ,
         \unit_memory/DRAM/n2572 , \unit_memory/DRAM/n2571 ,
         \unit_memory/DRAM/n2570 , \unit_memory/DRAM/n2569 ,
         \unit_memory/DRAM/n2568 , \unit_memory/DRAM/n2567 ,
         \unit_memory/DRAM/n2566 , \unit_memory/DRAM/n2565 ,
         \unit_memory/DRAM/n2564 , \unit_memory/DRAM/n2563 ,
         \unit_memory/DRAM/n2562 , \unit_memory/DRAM/n2561 ,
         \unit_memory/DRAM/n2560 , \unit_memory/DRAM/n2559 ,
         \unit_memory/DRAM/n2558 , \unit_memory/DRAM/n2557 ,
         \unit_memory/DRAM/n2556 , \unit_memory/DRAM/n2555 ,
         \unit_memory/DRAM/n2554 , \unit_memory/DRAM/n2553 ,
         \unit_memory/DRAM/n2552 , \unit_memory/DRAM/n2551 ,
         \unit_memory/DRAM/n2550 , \unit_memory/DRAM/n2549 ,
         \unit_memory/DRAM/n2548 , \unit_memory/DRAM/n2547 ,
         \unit_memory/DRAM/n2546 , \unit_memory/DRAM/n2545 ,
         \unit_memory/DRAM/n2544 , \unit_memory/DRAM/n2543 ,
         \unit_memory/DRAM/n2542 , \unit_memory/DRAM/n2541 ,
         \unit_memory/DRAM/n2540 , \unit_memory/DRAM/n2539 ,
         \unit_memory/DRAM/n2538 , \unit_memory/DRAM/n2537 ,
         \unit_memory/DRAM/n2536 , \unit_memory/DRAM/n2535 ,
         \unit_memory/DRAM/n2534 , \unit_memory/DRAM/n2533 ,
         \unit_memory/DRAM/n2532 , \unit_memory/DRAM/n2531 ,
         \unit_memory/DRAM/n2530 , \unit_memory/DRAM/n2529 ,
         \unit_memory/DRAM/n2528 , \unit_memory/DRAM/n2527 ,
         \unit_memory/DRAM/n2526 , \unit_memory/DRAM/n2525 ,
         \unit_memory/DRAM/n2524 , \unit_memory/DRAM/n2523 ,
         \unit_memory/DRAM/n2522 , \unit_memory/DRAM/n2521 ,
         \unit_memory/DRAM/n2520 , \unit_memory/DRAM/n2519 ,
         \unit_memory/DRAM/n2518 , \unit_memory/DRAM/n2517 ,
         \unit_memory/DRAM/n2516 , \unit_memory/DRAM/n2515 ,
         \unit_memory/DRAM/n2514 , \unit_memory/DRAM/n2513 ,
         \unit_memory/DRAM/n2512 , \unit_memory/DRAM/n2511 ,
         \unit_memory/DRAM/n2510 , \unit_memory/DRAM/n2509 ,
         \unit_memory/DRAM/n2508 , \unit_memory/DRAM/n2507 ,
         \unit_memory/DRAM/n2506 , \unit_memory/DRAM/n2505 ,
         \unit_memory/DRAM/n2504 , \unit_memory/DRAM/n2503 ,
         \unit_memory/DRAM/n2502 , \unit_memory/DRAM/n2501 ,
         \unit_memory/DRAM/n2500 , \unit_memory/DRAM/n2499 ,
         \unit_memory/DRAM/n2498 , \unit_memory/DRAM/n2497 ,
         \unit_memory/DRAM/n2496 , \unit_memory/DRAM/n2495 ,
         \unit_memory/DRAM/n2494 , \unit_memory/DRAM/n2493 ,
         \unit_memory/DRAM/n2492 , \unit_memory/DRAM/n2491 ,
         \unit_memory/DRAM/n2490 , \unit_memory/DRAM/n2489 ,
         \unit_memory/DRAM/n2488 , \unit_memory/DRAM/n2487 ,
         \unit_memory/DRAM/n2486 , \unit_memory/DRAM/n2485 ,
         \unit_memory/DRAM/n2484 , \unit_memory/DRAM/n2483 ,
         \unit_memory/DRAM/n2482 , \unit_memory/DRAM/n2481 ,
         \unit_memory/DRAM/n2480 , \unit_memory/DRAM/n2479 ,
         \unit_memory/DRAM/n2478 , \unit_memory/DRAM/n2477 ,
         \unit_memory/DRAM/n2476 , \unit_memory/DRAM/n2475 ,
         \unit_memory/DRAM/n2474 , \unit_memory/DRAM/n2473 ,
         \unit_memory/DRAM/n2472 , \unit_memory/DRAM/n2471 ,
         \unit_memory/DRAM/n2470 , \unit_memory/DRAM/n2469 ,
         \unit_memory/DRAM/n2468 , \unit_memory/DRAM/n2467 ,
         \unit_memory/DRAM/n2466 , \unit_memory/DRAM/n2465 ,
         \unit_memory/DRAM/n2464 , \unit_memory/DRAM/n2463 ,
         \unit_memory/DRAM/n2462 , \unit_memory/DRAM/n2461 ,
         \unit_memory/DRAM/n2460 , \unit_memory/DRAM/n2459 ,
         \unit_memory/DRAM/n2458 , \unit_memory/DRAM/n2457 ,
         \unit_memory/DRAM/n2456 , \unit_memory/DRAM/n2455 ,
         \unit_memory/DRAM/n2454 , \unit_memory/DRAM/n2453 ,
         \unit_memory/DRAM/n2452 , \unit_memory/DRAM/n2451 ,
         \unit_memory/DRAM/n2450 , \unit_memory/DRAM/n2449 ,
         \unit_memory/DRAM/n2448 , \unit_memory/DRAM/n2447 ,
         \unit_memory/DRAM/n2446 , \unit_memory/DRAM/n2445 ,
         \unit_memory/DRAM/n2444 , \unit_memory/DRAM/n2443 ,
         \unit_memory/DRAM/n2442 , \unit_memory/DRAM/n2441 ,
         \unit_memory/DRAM/n2440 , \unit_memory/DRAM/n2439 ,
         \unit_memory/DRAM/n2438 , \unit_memory/DRAM/n2437 ,
         \unit_memory/DRAM/n2436 , \unit_memory/DRAM/n2435 ,
         \unit_memory/DRAM/n2434 , \unit_memory/DRAM/n2433 ,
         \unit_memory/DRAM/n2432 , \unit_memory/DRAM/n2431 ,
         \unit_memory/DRAM/n2430 , \unit_memory/DRAM/n2429 ,
         \unit_memory/DRAM/n2428 , \unit_memory/DRAM/n2427 ,
         \unit_memory/DRAM/n2426 , \unit_memory/DRAM/n2425 ,
         \unit_memory/DRAM/n2424 , \unit_memory/DRAM/n2423 ,
         \unit_memory/DRAM/n2422 , \unit_memory/DRAM/n2421 ,
         \unit_memory/DRAM/n2420 , \unit_memory/DRAM/n2419 ,
         \unit_memory/DRAM/n2418 , \unit_memory/DRAM/n2417 ,
         \unit_memory/DRAM/n2416 , \unit_memory/DRAM/n2415 ,
         \unit_memory/DRAM/n2414 , \unit_memory/DRAM/n2413 ,
         \unit_memory/DRAM/n2412 , \unit_memory/DRAM/n2411 ,
         \unit_memory/DRAM/n2410 , \unit_memory/DRAM/n2409 ,
         \unit_memory/DRAM/n2408 , \unit_memory/DRAM/n2407 ,
         \unit_memory/DRAM/n2406 , \unit_memory/DRAM/n2405 ,
         \unit_memory/DRAM/n2404 , \unit_memory/DRAM/n2403 ,
         \unit_memory/DRAM/n2402 , \unit_memory/DRAM/n2401 ,
         \unit_memory/DRAM/n2400 , \unit_memory/DRAM/n2399 ,
         \unit_memory/DRAM/n2398 , \unit_memory/DRAM/n2397 ,
         \unit_memory/DRAM/n2396 , \unit_memory/DRAM/n2395 ,
         \unit_memory/DRAM/n2394 , \unit_memory/DRAM/n2393 ,
         \unit_memory/DRAM/n2392 , \unit_memory/DRAM/n2391 ,
         \unit_memory/DRAM/n2390 , \unit_memory/DRAM/n2389 ,
         \unit_memory/DRAM/n2388 , \unit_memory/DRAM/n2387 ,
         \unit_memory/DRAM/n2386 , \unit_memory/DRAM/n2385 ,
         \unit_memory/DRAM/n2384 , \unit_memory/DRAM/n2383 ,
         \unit_memory/DRAM/n2382 , \unit_memory/DRAM/n2381 ,
         \unit_memory/DRAM/n2380 , \unit_memory/DRAM/n2379 ,
         \unit_memory/DRAM/n2378 , \unit_memory/DRAM/n2377 ,
         \unit_memory/DRAM/n2376 , \unit_memory/DRAM/n2375 ,
         \unit_memory/DRAM/n2374 , \unit_memory/DRAM/n2373 ,
         \unit_memory/DRAM/n2372 , \unit_memory/DRAM/n2371 ,
         \unit_memory/DRAM/n2370 , \unit_memory/DRAM/n2369 ,
         \unit_memory/DRAM/n2368 , \unit_memory/DRAM/n2367 ,
         \unit_memory/DRAM/n2366 , \unit_memory/DRAM/n2365 ,
         \unit_memory/DRAM/n2364 , \unit_memory/DRAM/n2363 ,
         \unit_memory/DRAM/n2362 , \unit_memory/DRAM/n2361 ,
         \unit_memory/DRAM/n2360 , \unit_memory/DRAM/n2359 ,
         \unit_memory/DRAM/n2358 , \unit_memory/DRAM/n2357 ,
         \unit_memory/DRAM/n2356 , \unit_memory/DRAM/n2355 ,
         \unit_memory/DRAM/n2354 , \unit_memory/DRAM/n2353 ,
         \unit_memory/DRAM/n2352 , \unit_memory/DRAM/n2351 ,
         \unit_memory/DRAM/n2350 , \unit_memory/DRAM/n2349 ,
         \unit_memory/DRAM/n2348 , \unit_memory/DRAM/n2347 ,
         \unit_memory/DRAM/n2346 , \unit_memory/DRAM/n2345 ,
         \unit_memory/DRAM/n2344 , \unit_memory/DRAM/n2343 ,
         \unit_memory/DRAM/n2342 , \unit_memory/DRAM/n2341 ,
         \unit_memory/DRAM/n2340 , \unit_memory/DRAM/n2339 ,
         \unit_memory/DRAM/n2338 , \unit_memory/DRAM/n2337 ,
         \unit_memory/DRAM/n2336 , \unit_memory/DRAM/n2335 ,
         \unit_memory/DRAM/n2334 , \unit_memory/DRAM/n2333 ,
         \unit_memory/DRAM/n2332 , \unit_memory/DRAM/n2331 ,
         \unit_memory/DRAM/n2330 , \unit_memory/DRAM/n2329 ,
         \unit_memory/DRAM/n2328 , \unit_memory/DRAM/n2327 ,
         \unit_memory/DRAM/n2326 , \unit_memory/DRAM/n2325 ,
         \unit_memory/DRAM/n2324 , \unit_memory/DRAM/n2323 ,
         \unit_memory/DRAM/n2322 , \unit_memory/DRAM/n2321 ,
         \unit_memory/DRAM/n2320 , \unit_memory/DRAM/n2319 ,
         \unit_memory/DRAM/n2318 , \unit_memory/DRAM/n2317 ,
         \unit_memory/DRAM/n2316 , \unit_memory/DRAM/n2315 ,
         \unit_memory/DRAM/n2314 , \unit_memory/DRAM/n2313 ,
         \unit_memory/DRAM/n2312 , \unit_memory/DRAM/n2311 ,
         \unit_memory/DRAM/n2310 , \unit_memory/DRAM/n2309 ,
         \unit_memory/DRAM/n2308 , \unit_memory/DRAM/n2307 ,
         \unit_memory/DRAM/n2306 , \unit_memory/DRAM/n2305 ,
         \unit_memory/DRAM/n2304 , \unit_memory/DRAM/n2303 ,
         \unit_memory/DRAM/n2302 , \unit_memory/DRAM/n2301 ,
         \unit_memory/DRAM/n2300 , \unit_memory/DRAM/n2299 ,
         \unit_memory/DRAM/n2298 , \unit_memory/DRAM/n2297 ,
         \unit_memory/DRAM/n2296 , \unit_memory/DRAM/n2295 ,
         \unit_memory/DRAM/n2294 , \unit_memory/DRAM/n2293 ,
         \unit_memory/DRAM/n2292 , \unit_memory/DRAM/n2291 ,
         \unit_memory/DRAM/n2290 , \unit_memory/DRAM/n2289 ,
         \unit_memory/DRAM/n2288 , \unit_memory/DRAM/n2287 ,
         \unit_memory/DRAM/n2286 , \unit_memory/DRAM/n2285 ,
         \unit_memory/DRAM/n2284 , \unit_memory/DRAM/n2283 ,
         \unit_memory/DRAM/n2282 , \unit_memory/DRAM/n2281 ,
         \unit_memory/DRAM/n2280 , \unit_memory/DRAM/n2279 ,
         \unit_memory/DRAM/n2278 , \unit_memory/DRAM/n2277 ,
         \unit_memory/DRAM/n2276 , \unit_memory/DRAM/n2275 ,
         \unit_memory/DRAM/n2274 , \unit_memory/DRAM/n2273 ,
         \unit_memory/DRAM/n2272 , \unit_memory/DRAM/n2271 ,
         \unit_memory/DRAM/n2270 , \unit_memory/DRAM/n2269 ,
         \unit_memory/DRAM/n2268 , \unit_memory/DRAM/n2267 ,
         \unit_memory/DRAM/n2266 , \unit_memory/DRAM/n2265 ,
         \unit_memory/DRAM/n2264 , \unit_memory/DRAM/n2263 ,
         \unit_memory/DRAM/n2262 , \unit_memory/DRAM/n2261 ,
         \unit_memory/DRAM/n2260 , \unit_memory/DRAM/n2259 ,
         \unit_memory/DRAM/n2258 , \unit_memory/DRAM/n2257 ,
         \unit_memory/DRAM/n2256 , \unit_memory/DRAM/n2255 ,
         \unit_memory/DRAM/n2254 , \unit_memory/DRAM/n2253 ,
         \unit_memory/DRAM/n2252 , \unit_memory/DRAM/n2251 ,
         \unit_memory/DRAM/n2250 , \unit_memory/DRAM/n2249 ,
         \unit_memory/DRAM/n2248 , \unit_memory/DRAM/n2247 ,
         \unit_memory/DRAM/n2246 , \unit_memory/DRAM/n2245 ,
         \unit_memory/DRAM/n2244 , \unit_memory/DRAM/n2243 ,
         \unit_memory/DRAM/n2242 , \unit_memory/DRAM/n2241 ,
         \unit_memory/DRAM/n2240 , \unit_memory/DRAM/n2239 ,
         \unit_memory/DRAM/n2238 , \unit_memory/DRAM/n2237 ,
         \unit_memory/DRAM/n2236 , \unit_memory/DRAM/n2235 ,
         \unit_memory/DRAM/n2234 , \unit_memory/DRAM/n2233 ,
         \unit_memory/DRAM/n2232 , \unit_memory/DRAM/n2231 ,
         \unit_memory/DRAM/n2230 , \unit_memory/DRAM/n2229 ,
         \unit_memory/DRAM/n2228 , \unit_memory/DRAM/n2227 ,
         \unit_memory/DRAM/n2226 , \unit_memory/DRAM/n2225 ,
         \unit_memory/DRAM/n2224 , \unit_memory/DRAM/n2223 ,
         \unit_memory/DRAM/n2222 , \unit_memory/DRAM/n2221 ,
         \unit_memory/DRAM/n2220 , \unit_memory/DRAM/n2219 ,
         \unit_memory/DRAM/n2218 , \unit_memory/DRAM/n2217 ,
         \unit_memory/DRAM/n2216 , \unit_memory/DRAM/n2215 ,
         \unit_memory/DRAM/n2214 , \unit_memory/DRAM/n2213 ,
         \unit_memory/DRAM/n2212 , \unit_memory/DRAM/n2211 ,
         \unit_memory/DRAM/n2210 , \unit_memory/DRAM/n2209 ,
         \unit_memory/DRAM/n2208 , \unit_memory/DRAM/n2207 ,
         \unit_memory/DRAM/n2206 , \unit_memory/DRAM/n2205 ,
         \unit_memory/DRAM/n2204 , \unit_memory/DRAM/n2203 ,
         \unit_memory/DRAM/n2202 , \unit_memory/DRAM/n2201 ,
         \unit_memory/DRAM/n2200 , \unit_memory/DRAM/n2198 ,
         \unit_memory/DRAM/n2197 , \unit_memory/DRAM/n2196 ,
         \unit_memory/DRAM/n2195 , \unit_memory/DRAM/n2194 ,
         \unit_memory/DRAM/n2193 , \unit_memory/DRAM/n2192 ,
         \unit_memory/DRAM/n2191 , \unit_memory/DRAM/n2190 ,
         \unit_memory/DRAM/n2189 , \unit_memory/DRAM/n2188 ,
         \unit_memory/DRAM/n2187 , \unit_memory/DRAM/n2186 ,
         \unit_memory/DRAM/n2185 , \unit_memory/DRAM/n2184 ,
         \unit_memory/DRAM/n2183 , \unit_memory/DRAM/n2182 ,
         \unit_memory/DRAM/n2181 , \unit_memory/DRAM/n1156 ,
         \unit_memory/DRAM/n1155 , \unit_memory/DRAM/n1154 ,
         \unit_memory/DRAM/n1153 , \unit_memory/DRAM/n1152 ,
         \unit_memory/DRAM/n1151 , \unit_memory/DRAM/n1150 ,
         \unit_memory/DRAM/n1149 , \unit_memory/DRAM/n1148 ,
         \unit_memory/DRAM/n1147 , \unit_memory/DRAM/n1146 ,
         \unit_memory/DRAM/n1145 , \unit_memory/DRAM/n1144 ,
         \unit_memory/DRAM/n1143 , \unit_memory/DRAM/n1142 ,
         \unit_memory/DRAM/n1141 , \unit_memory/DRAM/n1140 ,
         \unit_memory/DRAM/n1139 , \unit_memory/DRAM/n1138 ,
         \unit_memory/DRAM/n1137 , \unit_memory/DRAM/n1135 ,
         \unit_memory/DRAM/n1134 , \unit_memory/DRAM/n1133 ,
         \unit_memory/DRAM/n1132 , \unit_memory/DRAM/n1131 ,
         \unit_memory/DRAM/n1130 , \unit_memory/DRAM/n1129 ,
         \unit_memory/DRAM/n1128 , \unit_memory/DRAM/n1127 ,
         \unit_memory/DRAM/n1126 , \unit_memory/DRAM/n1125 ,
         \unit_memory/DRAM/n1124 , \unit_memory/DRAM/n1123 ,
         \unit_memory/DRAM/n1122 , \unit_memory/DRAM/n1121 ,
         \unit_memory/DRAM/n1120 , \unit_memory/DRAM/n1119 ,
         \unit_memory/DRAM/n1118 , \unit_memory/DRAM/n1117 ,
         \unit_memory/DRAM/n1116 , \unit_memory/DRAM/n1115 ,
         \unit_memory/DRAM/n1114 , \unit_memory/DRAM/n1113 ,
         \unit_memory/DRAM/n1112 , \unit_memory/DRAM/n1111 ,
         \unit_memory/DRAM/n1110 , \unit_memory/DRAM/n1109 ,
         \unit_memory/DRAM/n1108 , \unit_memory/DRAM/n1107 ,
         \unit_memory/DRAM/n1106 , \unit_memory/DRAM/n1105 ,
         \unit_memory/DRAM/n1104 , \unit_memory/DRAM/n1103 ,
         \unit_memory/DRAM/n1102 , \unit_memory/DRAM/n1101 ,
         \unit_memory/DRAM/n1100 , \unit_memory/DRAM/n1099 ,
         \unit_memory/DRAM/n1098 , \unit_memory/DRAM/n1097 ,
         \unit_memory/DRAM/n1096 , \unit_memory/DRAM/n1095 ,
         \unit_memory/DRAM/n1094 , \unit_memory/DRAM/n1093 ,
         \unit_memory/DRAM/n1092 , \unit_memory/DRAM/n1091 ,
         \unit_memory/DRAM/n1090 , \unit_memory/DRAM/n1089 ,
         \unit_memory/DRAM/n1088 , \unit_memory/DRAM/n1087 ,
         \unit_memory/DRAM/n1086 , \unit_memory/DRAM/n1085 ,
         \unit_memory/DRAM/n1084 , \unit_memory/DRAM/n1083 ,
         \unit_memory/DRAM/n1082 , \unit_memory/DRAM/n1081 ,
         \unit_memory/DRAM/n1080 , \unit_memory/DRAM/n1079 ,
         \unit_memory/DRAM/n1078 , \unit_memory/DRAM/n1077 ,
         \unit_memory/DRAM/n1076 , \unit_memory/DRAM/n1075 ,
         \unit_memory/DRAM/n1074 , \unit_memory/DRAM/n1073 ,
         \unit_memory/DRAM/n1072 , \unit_memory/DRAM/n1071 ,
         \unit_memory/DRAM/n1070 , \unit_memory/DRAM/n1069 ,
         \unit_memory/DRAM/n1068 , \unit_memory/DRAM/n1067 ,
         \unit_memory/DRAM/n1066 , \unit_memory/DRAM/n1065 ,
         \unit_memory/DRAM/n1064 , \unit_memory/DRAM/n1063 ,
         \unit_memory/DRAM/n1062 , \unit_memory/DRAM/n1061 ,
         \unit_memory/DRAM/n1060 , \unit_memory/DRAM/n1059 ,
         \unit_memory/DRAM/n1058 , \unit_memory/DRAM/n1057 ,
         \unit_memory/DRAM/n1056 , \unit_memory/DRAM/n1055 ,
         \unit_memory/DRAM/n1054 , \unit_memory/DRAM/n1053 ,
         \unit_memory/DRAM/n1052 , \unit_memory/DRAM/n1051 ,
         \unit_memory/DRAM/n1050 , \unit_memory/DRAM/n1049 ,
         \unit_memory/DRAM/n1048 , \unit_memory/DRAM/n1047 ,
         \unit_memory/DRAM/n1046 , \unit_memory/DRAM/n1045 ,
         \unit_memory/DRAM/n1044 , \unit_memory/DRAM/n1043 ,
         \unit_memory/DRAM/n1042 , \unit_memory/DRAM/n1041 ,
         \unit_memory/DRAM/n1040 , \unit_memory/DRAM/n1039 ,
         \unit_memory/DRAM/n1038 , \unit_memory/DRAM/n1037 ,
         \unit_memory/DRAM/n1036 , \unit_memory/DRAM/n1035 ,
         \unit_memory/DRAM/n1034 , \unit_memory/DRAM/n1033 ,
         \unit_memory/DRAM/n1032 , \unit_memory/DRAM/n1031 ,
         \unit_memory/DRAM/n1030 , \unit_memory/DRAM/n1029 ,
         \unit_memory/DRAM/n1028 , \unit_memory/DRAM/n1027 ,
         \unit_memory/DRAM/n1026 , \unit_memory/DRAM/n1025 ,
         \unit_memory/DRAM/n1024 , \unit_memory/DRAM/n1023 ,
         \unit_memory/DRAM/n1022 , \unit_memory/DRAM/n1021 ,
         \unit_memory/DRAM/n1020 , \unit_memory/DRAM/n1019 ,
         \unit_memory/DRAM/n1018 , \unit_memory/DRAM/n1017 ,
         \unit_memory/DRAM/n1016 , \unit_memory/DRAM/n1015 ,
         \unit_memory/DRAM/n1014 , \unit_memory/DRAM/n1013 ,
         \unit_memory/DRAM/n1012 , \unit_memory/DRAM/n1011 ,
         \unit_memory/DRAM/n1010 , \unit_memory/DRAM/n1009 ,
         \unit_memory/DRAM/n1008 , \unit_memory/DRAM/n1007 ,
         \unit_memory/DRAM/n1006 , \unit_memory/DRAM/n1005 ,
         \unit_memory/DRAM/n1004 , \unit_memory/DRAM/n1003 ,
         \unit_memory/DRAM/n1002 , \unit_memory/DRAM/n1001 ,
         \unit_memory/DRAM/n1000 , \unit_memory/DRAM/n999 ,
         \unit_memory/DRAM/n998 , \unit_memory/DRAM/n997 ,
         \unit_memory/DRAM/n996 , \unit_memory/DRAM/n995 ,
         \unit_memory/DRAM/n994 , \unit_memory/DRAM/n993 ,
         \unit_memory/DRAM/n992 , \unit_memory/DRAM/n991 ,
         \unit_memory/DRAM/n990 , \unit_memory/DRAM/n989 ,
         \unit_memory/DRAM/n988 , \unit_memory/DRAM/n987 ,
         \unit_memory/DRAM/n986 , \unit_memory/DRAM/n985 ,
         \unit_memory/DRAM/n984 , \unit_memory/DRAM/n983 ,
         \unit_memory/DRAM/n982 , \unit_memory/DRAM/n981 ,
         \unit_memory/DRAM/n980 , \unit_memory/DRAM/n979 ,
         \unit_memory/DRAM/n978 , \unit_memory/DRAM/n977 ,
         \unit_memory/DRAM/n976 , \unit_memory/DRAM/n975 ,
         \unit_memory/DRAM/n974 , \unit_memory/DRAM/n973 ,
         \unit_memory/DRAM/n972 , \unit_memory/DRAM/n971 ,
         \unit_memory/DRAM/n970 , \unit_memory/DRAM/n969 ,
         \unit_memory/DRAM/n968 , \unit_memory/DRAM/n967 ,
         \unit_memory/DRAM/n966 , \unit_memory/DRAM/n965 ,
         \unit_memory/DRAM/n964 , \unit_memory/DRAM/n963 ,
         \unit_memory/DRAM/n962 , \unit_memory/DRAM/n961 ,
         \unit_memory/DRAM/n960 , \unit_memory/DRAM/n959 ,
         \unit_memory/DRAM/n958 , \unit_memory/DRAM/n957 ,
         \unit_memory/DRAM/n956 , \unit_memory/DRAM/n955 ,
         \unit_memory/DRAM/n954 , \unit_memory/DRAM/n953 ,
         \unit_memory/DRAM/n952 , \unit_memory/DRAM/n951 ,
         \unit_memory/DRAM/n950 , \unit_memory/DRAM/n949 ,
         \unit_memory/DRAM/n948 , \unit_memory/DRAM/n947 ,
         \unit_memory/DRAM/n946 , \unit_memory/DRAM/n945 ,
         \unit_memory/DRAM/n944 , \unit_memory/DRAM/n943 ,
         \unit_memory/DRAM/n942 , \unit_memory/DRAM/n941 ,
         \unit_memory/DRAM/n940 , \unit_memory/DRAM/n939 ,
         \unit_memory/DRAM/n938 , \unit_memory/DRAM/n937 ,
         \unit_memory/DRAM/n936 , \unit_memory/DRAM/n935 ,
         \unit_memory/DRAM/n934 , \unit_memory/DRAM/n933 ,
         \unit_memory/DRAM/n932 , \unit_memory/DRAM/n931 ,
         \unit_memory/DRAM/n930 , \unit_memory/DRAM/n929 ,
         \unit_memory/DRAM/n928 , \unit_memory/DRAM/n927 ,
         \unit_memory/DRAM/n926 , \unit_memory/DRAM/n925 ,
         \unit_memory/DRAM/n924 , \unit_memory/DRAM/n923 ,
         \unit_memory/DRAM/n922 , \unit_memory/DRAM/n921 ,
         \unit_memory/DRAM/n920 , \unit_memory/DRAM/n919 ,
         \unit_memory/DRAM/n918 , \unit_memory/DRAM/n917 ,
         \unit_memory/DRAM/n916 , \unit_memory/DRAM/n915 ,
         \unit_memory/DRAM/n914 , \unit_memory/DRAM/n913 ,
         \unit_memory/DRAM/n912 , \unit_memory/DRAM/n911 ,
         \unit_memory/DRAM/n910 , \unit_memory/DRAM/n909 ,
         \unit_memory/DRAM/n908 , \unit_memory/DRAM/n907 ,
         \unit_memory/DRAM/n906 , \unit_memory/DRAM/n905 ,
         \unit_memory/DRAM/n904 , \unit_memory/DRAM/n903 ,
         \unit_memory/DRAM/n902 , \unit_memory/DRAM/n901 ,
         \unit_memory/DRAM/n900 , \unit_memory/DRAM/n899 ,
         \unit_memory/DRAM/n898 , \unit_memory/DRAM/n897 ,
         \unit_memory/DRAM/n896 , \unit_memory/DRAM/n895 ,
         \unit_memory/DRAM/n894 , \unit_memory/DRAM/n893 ,
         \unit_memory/DRAM/n892 , \unit_memory/DRAM/n891 ,
         \unit_memory/DRAM/n890 , \unit_memory/DRAM/n889 ,
         \unit_memory/DRAM/n888 , \unit_memory/DRAM/n887 ,
         \unit_memory/DRAM/n886 , \unit_memory/DRAM/n885 ,
         \unit_memory/DRAM/n884 , \unit_memory/DRAM/n883 ,
         \unit_memory/DRAM/n882 , \unit_memory/DRAM/n881 ,
         \unit_memory/DRAM/n880 , \unit_memory/DRAM/n879 ,
         \unit_memory/DRAM/n878 , \unit_memory/DRAM/n877 ,
         \unit_memory/DRAM/n876 , \unit_memory/DRAM/n875 ,
         \unit_memory/DRAM/n874 , \unit_memory/DRAM/n873 ,
         \unit_memory/DRAM/n872 , \unit_memory/DRAM/n871 ,
         \unit_memory/DRAM/n870 , \unit_memory/DRAM/n869 ,
         \unit_memory/DRAM/n868 , \unit_memory/DRAM/n867 ,
         \unit_memory/DRAM/n866 , \unit_memory/DRAM/n865 ,
         \unit_memory/DRAM/n864 , \unit_memory/DRAM/n863 ,
         \unit_memory/DRAM/n862 , \unit_memory/DRAM/n861 ,
         \unit_memory/DRAM/n860 , \unit_memory/DRAM/n859 ,
         \unit_memory/DRAM/n858 , \unit_memory/DRAM/n857 ,
         \unit_memory/DRAM/n856 , \unit_memory/DRAM/n855 ,
         \unit_memory/DRAM/n854 , \unit_memory/DRAM/n853 ,
         \unit_memory/DRAM/n852 , \unit_memory/DRAM/n851 ,
         \unit_memory/DRAM/n850 , \unit_memory/DRAM/n849 ,
         \unit_memory/DRAM/n848 , \unit_memory/DRAM/n847 ,
         \unit_memory/DRAM/n846 , \unit_memory/DRAM/n845 ,
         \unit_memory/DRAM/n844 , \unit_memory/DRAM/n843 ,
         \unit_memory/DRAM/n842 , \unit_memory/DRAM/n841 ,
         \unit_memory/DRAM/n840 , \unit_memory/DRAM/n839 ,
         \unit_memory/DRAM/n838 , \unit_memory/DRAM/n837 ,
         \unit_memory/DRAM/n836 , \unit_memory/DRAM/n835 ,
         \unit_memory/DRAM/n834 , \unit_memory/DRAM/n833 ,
         \unit_memory/DRAM/n832 , \unit_memory/DRAM/n831 ,
         \unit_memory/DRAM/n830 , \unit_memory/DRAM/n829 ,
         \unit_memory/DRAM/n828 , \unit_memory/DRAM/n827 ,
         \unit_memory/DRAM/n826 , \unit_memory/DRAM/n825 ,
         \unit_memory/DRAM/n824 , \unit_memory/DRAM/n823 ,
         \unit_memory/DRAM/n822 , \unit_memory/DRAM/n821 ,
         \unit_memory/DRAM/n820 , \unit_memory/DRAM/n819 ,
         \unit_memory/DRAM/n818 , \unit_memory/DRAM/n817 ,
         \unit_memory/DRAM/n815 , \unit_memory/DRAM/n814 ,
         \unit_memory/DRAM/n813 , \unit_memory/DRAM/n812 ,
         \unit_memory/DRAM/n811 , \unit_memory/DRAM/n809 ,
         \unit_memory/DRAM/n801 , \unit_memory/DRAM/n794 ,
         \unit_memory/DRAM/n792 , \unit_memory/DRAM/n784 ,
         \unit_memory/DRAM/n782 , \unit_memory/DRAM/n774 ,
         \unit_memory/DRAM/n772 , \unit_memory/DRAM/n771 ,
         \unit_memory/DRAM/n770 , \unit_memory/DRAM/n768 ,
         \unit_memory/DRAM/n766 , \unit_memory/DRAM/n764 ,
         \unit_memory/DRAM/n762 , \unit_memory/DRAM/n760 ,
         \unit_memory/DRAM/n758 , \unit_memory/DRAM/n756 ,
         \unit_memory/DRAM/n755 , \unit_memory/DRAM/n754 ,
         \unit_memory/DRAM/n753 , \unit_memory/DRAM/n752 ,
         \unit_memory/DRAM/n751 , \unit_memory/DRAM/n750 ,
         \unit_memory/DRAM/n749 , \unit_memory/DRAM/n748 ,
         \unit_memory/DRAM/n747 , \unit_memory/DRAM/n746 ,
         \unit_memory/DRAM/n745 , \unit_memory/DRAM/n744 ,
         \unit_memory/DRAM/n743 , \unit_memory/DRAM/n742 ,
         \unit_memory/DRAM/n741 , \unit_memory/DRAM/n740 ,
         \unit_memory/DRAM/n739 , \unit_memory/DRAM/n738 ,
         \unit_memory/DRAM/n737 , \unit_memory/DRAM/n736 ,
         \unit_memory/DRAM/n735 , \unit_memory/DRAM/n734 ,
         \unit_memory/DRAM/n733 , \unit_memory/DRAM/n732 ,
         \unit_memory/DRAM/n731 , \unit_memory/DRAM/n730 ,
         \unit_memory/DRAM/n729 , \unit_memory/DRAM/n728 ,
         \unit_memory/DRAM/n727 , \unit_memory/DRAM/n726 ,
         \unit_memory/DRAM/n725 , \unit_memory/DRAM/n724 ,
         \unit_memory/DRAM/n723 , \unit_memory/DRAM/n722 ,
         \unit_memory/DRAM/n719 , \unit_memory/DRAM/n718 ,
         \unit_memory/DRAM/n717 , \unit_memory/DRAM/n716 ,
         \unit_memory/DRAM/n715 , \unit_memory/DRAM/n714 ,
         \unit_memory/DRAM/n713 , \unit_memory/DRAM/n712 ,
         \unit_memory/DRAM/n711 , \unit_memory/DRAM/n710 ,
         \unit_memory/DRAM/n709 , \unit_memory/DRAM/n708 ,
         \unit_memory/DRAM/n707 , \unit_memory/DRAM/n706 ,
         \unit_memory/DRAM/n705 , \unit_memory/DRAM/n704 ,
         \unit_memory/DRAM/n703 , \unit_memory/DRAM/n702 ,
         \unit_memory/DRAM/n701 , \unit_memory/DRAM/n700 ,
         \unit_memory/DRAM/n699 , \unit_memory/DRAM/n698 ,
         \unit_memory/DRAM/n697 , \unit_memory/DRAM/n696 ,
         \unit_memory/DRAM/n695 , \unit_memory/DRAM/n694 ,
         \unit_memory/DRAM/n693 , \unit_memory/DRAM/n692 ,
         \unit_memory/DRAM/n691 , \unit_memory/DRAM/n690 ,
         \unit_memory/DRAM/n689 , \unit_memory/DRAM/n688 ,
         \unit_memory/DRAM/n687 , \unit_memory/DRAM/n686 ,
         \unit_memory/DRAM/n685 , \unit_memory/DRAM/n684 ,
         \unit_memory/DRAM/n683 , \unit_memory/DRAM/n682 ,
         \unit_memory/DRAM/n681 , \unit_memory/DRAM/n680 ,
         \unit_memory/DRAM/n679 , \unit_memory/DRAM/n678 ,
         \unit_memory/DRAM/n677 , \unit_memory/DRAM/n676 ,
         \unit_memory/DRAM/n675 , \unit_memory/DRAM/n674 ,
         \unit_memory/DRAM/n673 , \unit_memory/DRAM/n672 ,
         \unit_memory/DRAM/n671 , \unit_memory/DRAM/n670 ,
         \unit_memory/DRAM/n669 , \unit_memory/DRAM/n668 ,
         \unit_memory/DRAM/n667 , \unit_memory/DRAM/n666 ,
         \unit_memory/DRAM/n665 , \unit_memory/DRAM/n664 ,
         \unit_memory/DRAM/n663 , \unit_memory/DRAM/n662 ,
         \unit_memory/DRAM/n661 , \unit_memory/DRAM/n660 ,
         \unit_memory/DRAM/n659 , \unit_memory/DRAM/n658 ,
         \unit_memory/DRAM/n657 , \unit_memory/DRAM/n656 ,
         \unit_memory/DRAM/n655 , \unit_memory/DRAM/n654 ,
         \unit_memory/DRAM/n653 , \unit_memory/DRAM/n652 ,
         \unit_memory/DRAM/n651 , \unit_memory/DRAM/n650 ,
         \unit_memory/DRAM/n649 , \unit_memory/DRAM/n648 ,
         \unit_memory/DRAM/n647 , \unit_memory/DRAM/n646 ,
         \unit_memory/DRAM/n645 , \unit_memory/DRAM/n644 ,
         \unit_memory/DRAM/n643 , \unit_memory/DRAM/n642 ,
         \unit_memory/DRAM/n641 , \unit_memory/DRAM/n640 ,
         \unit_memory/DRAM/n639 , \unit_memory/DRAM/n638 ,
         \unit_memory/DRAM/n637 , \unit_memory/DRAM/n636 ,
         \unit_memory/DRAM/n635 , \unit_memory/DRAM/n634 ,
         \unit_memory/DRAM/n633 , \unit_memory/DRAM/n632 ,
         \unit_memory/DRAM/n631 , \unit_memory/DRAM/n630 ,
         \unit_memory/DRAM/n629 , \unit_memory/DRAM/n628 ,
         \unit_memory/DRAM/n627 , \unit_memory/DRAM/n626 ,
         \unit_memory/DRAM/n625 , \unit_memory/DRAM/n624 ,
         \unit_memory/DRAM/n623 , \unit_memory/DRAM/n622 ,
         \unit_memory/DRAM/n621 , \unit_memory/DRAM/n620 ,
         \unit_memory/DRAM/n619 , \unit_memory/DRAM/n618 ,
         \unit_memory/DRAM/n617 , \unit_memory/DRAM/n616 ,
         \unit_memory/DRAM/n615 , \unit_memory/DRAM/n614 ,
         \unit_memory/DRAM/n613 , \unit_memory/DRAM/n612 ,
         \unit_memory/DRAM/n611 , \unit_memory/DRAM/n610 ,
         \unit_memory/DRAM/n609 , \unit_memory/DRAM/n608 ,
         \unit_memory/DRAM/n607 , \unit_memory/DRAM/n606 ,
         \unit_memory/DRAM/n605 , \unit_memory/DRAM/n604 ,
         \unit_memory/DRAM/n603 , \unit_memory/DRAM/n602 ,
         \unit_memory/DRAM/n601 , \unit_memory/DRAM/n600 ,
         \unit_memory/DRAM/n599 , \unit_memory/DRAM/n598 ,
         \unit_memory/DRAM/n597 , \unit_memory/DRAM/n596 ,
         \unit_memory/DRAM/n595 , \unit_memory/DRAM/n594 ,
         \unit_memory/DRAM/n593 , \unit_memory/DRAM/n592 ,
         \unit_memory/DRAM/n591 , \unit_memory/DRAM/n590 ,
         \unit_memory/DRAM/n589 , \unit_memory/DRAM/n588 ,
         \unit_memory/DRAM/n587 , \unit_memory/DRAM/n586 ,
         \unit_memory/DRAM/n585 , \unit_memory/DRAM/n584 ,
         \unit_memory/DRAM/n583 , \unit_memory/DRAM/n582 ,
         \unit_memory/DRAM/n581 , \unit_memory/DRAM/n580 ,
         \unit_memory/DRAM/n579 , \unit_memory/DRAM/n578 ,
         \unit_memory/DRAM/n577 , \unit_memory/DRAM/n576 ,
         \unit_memory/DRAM/n575 , \unit_memory/DRAM/n574 ,
         \unit_memory/DRAM/n573 , \unit_memory/DRAM/n572 ,
         \unit_memory/DRAM/n571 , \unit_memory/DRAM/n570 ,
         \unit_memory/DRAM/n569 , \unit_memory/DRAM/n568 ,
         \unit_memory/DRAM/n567 , \unit_memory/DRAM/n566 ,
         \unit_memory/DRAM/n565 , \unit_memory/DRAM/n564 ,
         \unit_memory/DRAM/n563 , \unit_memory/DRAM/n561 ,
         \unit_memory/DRAM/n552 , \unit_memory/DRAM/n551 ,
         \unit_memory/DRAM/n550 , \unit_memory/DRAM/n549 ,
         \unit_memory/DRAM/n548 , \unit_memory/DRAM/n547 ,
         \unit_memory/DRAM/n546 , \unit_memory/DRAM/n512 ,
         \unit_memory/DRAM/n511 , \unit_memory/DRAM/n510 ,
         \unit_memory/DRAM/n509 , \unit_memory/DRAM/n508 ,
         \unit_memory/DRAM/n507 , \unit_memory/DRAM/n506 ,
         \unit_memory/DRAM/n505 , \unit_memory/DRAM/n504 ,
         \unit_memory/DRAM/n503 , \unit_memory/DRAM/n502 ,
         \unit_memory/DRAM/n501 , \unit_memory/DRAM/n500 ,
         \unit_memory/DRAM/n499 , \unit_memory/DRAM/n498 ,
         \unit_memory/DRAM/n497 , \unit_memory/DRAM/n496 ,
         \unit_memory/DRAM/n495 , \unit_memory/DRAM/n494 ,
         \unit_memory/DRAM/n493 , \unit_memory/DRAM/n492 ,
         \unit_memory/DRAM/n491 , \unit_memory/DRAM/n490 ,
         \unit_memory/DRAM/n489 , \unit_memory/DRAM/n488 ,
         \unit_memory/DRAM/n487 , \unit_memory/DRAM/n486 ,
         \unit_memory/DRAM/n485 , \unit_memory/DRAM/n484 ,
         \unit_memory/DRAM/n483 , \unit_memory/DRAM/n482 ,
         \unit_memory/DRAM/n481 , \unit_memory/DRAM/n480 ,
         \unit_memory/DRAM/n479 , \unit_memory/DRAM/n478 ,
         \unit_memory/DRAM/n477 , \unit_memory/DRAM/n476 ,
         \unit_memory/DRAM/n475 , \unit_memory/DRAM/n474 ,
         \unit_memory/DRAM/n473 , \unit_memory/DRAM/n472 ,
         \unit_memory/DRAM/n471 , \unit_memory/DRAM/n470 ,
         \unit_memory/DRAM/n469 , \unit_memory/DRAM/n468 ,
         \unit_memory/DRAM/n467 , \unit_memory/DRAM/n466 ,
         \unit_memory/DRAM/n465 , \unit_memory/DRAM/n464 ,
         \unit_memory/DRAM/n463 , \unit_memory/DRAM/n462 ,
         \unit_memory/DRAM/n461 , \unit_memory/DRAM/n460 ,
         \unit_memory/DRAM/n459 , \unit_memory/DRAM/n458 ,
         \unit_memory/DRAM/n457 , \unit_memory/DRAM/n456 ,
         \unit_memory/DRAM/n455 , \unit_memory/DRAM/n454 ,
         \unit_memory/DRAM/n453 , \unit_memory/DRAM/n452 ,
         \unit_memory/DRAM/n451 , \unit_memory/DRAM/n450 ,
         \unit_memory/DRAM/n449 , \unit_memory/DRAM/n448 ,
         \unit_memory/DRAM/n447 , \unit_memory/DRAM/n446 ,
         \unit_memory/DRAM/n445 , \unit_memory/DRAM/n444 ,
         \unit_memory/DRAM/n443 , \unit_memory/DRAM/n442 ,
         \unit_memory/DRAM/n441 , \unit_memory/DRAM/n440 ,
         \unit_memory/DRAM/n439 , \unit_memory/DRAM/n438 ,
         \unit_memory/DRAM/n437 , \unit_memory/DRAM/n436 ,
         \unit_memory/DRAM/n435 , \unit_memory/DRAM/n434 ,
         \unit_memory/DRAM/n433 , \unit_memory/DRAM/n432 ,
         \unit_memory/DRAM/n431 , \unit_memory/DRAM/n430 ,
         \unit_memory/DRAM/n429 , \unit_memory/DRAM/n428 ,
         \unit_memory/DRAM/n427 , \unit_memory/DRAM/n426 ,
         \unit_memory/DRAM/n425 , \unit_memory/DRAM/n424 ,
         \unit_memory/DRAM/n423 , \unit_memory/DRAM/n422 ,
         \unit_memory/DRAM/n421 , \unit_memory/DRAM/n420 ,
         \unit_memory/DRAM/n419 , \unit_memory/DRAM/n418 ,
         \unit_memory/DRAM/n417 , \unit_memory/DRAM/n416 ,
         \unit_memory/DRAM/n415 , \unit_memory/DRAM/n414 ,
         \unit_memory/DRAM/n413 , \unit_memory/DRAM/n412 ,
         \unit_memory/DRAM/n411 , \unit_memory/DRAM/n410 ,
         \unit_memory/DRAM/n409 , \unit_memory/DRAM/n408 ,
         \unit_memory/DRAM/n407 , \unit_memory/DRAM/n406 ,
         \unit_memory/DRAM/n405 , \unit_memory/DRAM/n404 ,
         \unit_memory/DRAM/n403 , \unit_memory/DRAM/n402 ,
         \unit_memory/DRAM/n401 , \unit_memory/DRAM/n400 ,
         \unit_memory/DRAM/n399 , \unit_memory/DRAM/n398 ,
         \unit_memory/DRAM/n397 , \unit_memory/DRAM/n396 ,
         \unit_memory/DRAM/n395 , \unit_memory/DRAM/n394 ,
         \unit_memory/DRAM/n393 , \unit_memory/DRAM/n392 ,
         \unit_memory/DRAM/n391 , \unit_memory/DRAM/n390 ,
         \unit_memory/DRAM/n389 , \unit_memory/DRAM/n388 ,
         \unit_memory/DRAM/n387 , \unit_memory/DRAM/n386 ,
         \unit_memory/DRAM/n385 , \unit_memory/DRAM/n384 ,
         \unit_memory/DRAM/n383 , \unit_memory/DRAM/n382 ,
         \unit_memory/DRAM/n381 , \unit_memory/DRAM/n380 ,
         \unit_memory/DRAM/n379 , \unit_memory/DRAM/n378 ,
         \unit_memory/DRAM/n377 , \unit_memory/DRAM/n376 ,
         \unit_memory/DRAM/n375 , \unit_memory/DRAM/n374 ,
         \unit_memory/DRAM/n373 , \unit_memory/DRAM/n372 ,
         \unit_memory/DRAM/n371 , \unit_memory/DRAM/n370 ,
         \unit_memory/DRAM/n369 , \unit_memory/DRAM/n368 ,
         \unit_memory/DRAM/n367 , \unit_memory/DRAM/n366 ,
         \unit_memory/DRAM/n365 , \unit_memory/DRAM/n364 ,
         \unit_memory/DRAM/n363 , \unit_memory/DRAM/n362 ,
         \unit_memory/DRAM/n361 , \unit_memory/DRAM/n360 ,
         \unit_memory/DRAM/n359 , \unit_memory/DRAM/n358 ,
         \unit_memory/DRAM/n357 , \unit_memory/DRAM/n356 ,
         \unit_memory/DRAM/n355 , \unit_memory/DRAM/n354 ,
         \unit_memory/DRAM/n353 , \unit_memory/DRAM/n352 ,
         \unit_memory/DRAM/n351 , \unit_memory/DRAM/n350 ,
         \unit_memory/DRAM/n349 , \unit_memory/DRAM/n348 ,
         \unit_memory/DRAM/n347 , \unit_memory/DRAM/n346 ,
         \unit_memory/DRAM/n345 , \unit_memory/DRAM/n344 ,
         \unit_memory/DRAM/n343 , \unit_memory/DRAM/n342 ,
         \unit_memory/DRAM/n341 , \unit_memory/DRAM/n340 ,
         \unit_memory/DRAM/n339 , \unit_memory/DRAM/n338 ,
         \unit_memory/DRAM/n337 , \unit_memory/DRAM/n336 ,
         \unit_memory/DRAM/n335 , \unit_memory/DRAM/n334 ,
         \unit_memory/DRAM/n333 , \unit_memory/DRAM/n332 ,
         \unit_memory/DRAM/n331 , \unit_memory/DRAM/n330 ,
         \unit_memory/DRAM/n329 , \unit_memory/DRAM/n328 ,
         \unit_memory/DRAM/n327 , \unit_memory/DRAM/n326 ,
         \unit_memory/DRAM/n325 , \unit_memory/DRAM/n324 ,
         \unit_memory/DRAM/n323 , \unit_memory/DRAM/n322 ,
         \unit_memory/DRAM/n321 , \unit_memory/DRAM/n320 ,
         \unit_memory/DRAM/n319 , \unit_memory/DRAM/n318 ,
         \unit_memory/DRAM/n317 , \unit_memory/DRAM/n316 ,
         \unit_memory/DRAM/n315 , \unit_memory/DRAM/n314 ,
         \unit_memory/DRAM/n313 , \unit_memory/DRAM/n312 ,
         \unit_memory/DRAM/n311 , \unit_memory/DRAM/n310 ,
         \unit_memory/DRAM/n309 , \unit_memory/DRAM/n308 ,
         \unit_memory/DRAM/n307 , \unit_memory/DRAM/n306 ,
         \unit_memory/DRAM/n305 , \unit_memory/DRAM/n304 ,
         \unit_memory/DRAM/n303 , \unit_memory/DRAM/n302 ,
         \unit_memory/DRAM/n301 , \unit_memory/DRAM/n300 ,
         \unit_memory/DRAM/n299 , \unit_memory/DRAM/n298 ,
         \unit_memory/DRAM/n297 , \unit_memory/DRAM/n296 ,
         \unit_memory/DRAM/n295 , \unit_memory/DRAM/n294 ,
         \unit_memory/DRAM/n293 , \unit_memory/DRAM/n292 ,
         \unit_memory/DRAM/n291 , \unit_memory/DRAM/n290 ,
         \unit_memory/DRAM/n289 , \unit_memory/DRAM/n288 ,
         \unit_memory/DRAM/n287 , \unit_memory/DRAM/n286 ,
         \unit_memory/DRAM/n285 , \unit_memory/DRAM/n284 ,
         \unit_memory/DRAM/n283 , \unit_memory/DRAM/n282 ,
         \unit_memory/DRAM/n281 , \unit_memory/DRAM/n280 ,
         \unit_memory/DRAM/n279 , \unit_memory/DRAM/n278 ,
         \unit_memory/DRAM/n277 , \unit_memory/DRAM/n276 ,
         \unit_memory/DRAM/n275 , \unit_memory/DRAM/n274 ,
         \unit_memory/DRAM/n273 , \unit_memory/DRAM/n272 ,
         \unit_memory/DRAM/n271 , \unit_memory/DRAM/n270 ,
         \unit_memory/DRAM/n269 , \unit_memory/DRAM/n268 ,
         \unit_memory/DRAM/n267 , \unit_memory/DRAM/n266 ,
         \unit_memory/DRAM/n265 , \unit_memory/DRAM/n264 ,
         \unit_memory/DRAM/n263 , \unit_memory/DRAM/n262 ,
         \unit_memory/DRAM/n261 , \unit_memory/DRAM/n260 ,
         \unit_memory/DRAM/n259 , \unit_memory/DRAM/n258 ,
         \unit_memory/DRAM/n257 , \unit_memory/DRAM/n256 ,
         \unit_memory/DRAM/n255 , \unit_memory/DRAM/n254 ,
         \unit_memory/DRAM/n253 , \unit_memory/DRAM/n252 ,
         \unit_memory/DRAM/n251 , \unit_memory/DRAM/n250 ,
         \unit_memory/DRAM/n249 , \unit_memory/DRAM/n248 ,
         \unit_memory/DRAM/n247 , \unit_memory/DRAM/n246 ,
         \unit_memory/DRAM/n245 , \unit_memory/DRAM/n244 ,
         \unit_memory/DRAM/n243 , \unit_memory/DRAM/n242 ,
         \unit_memory/DRAM/n241 , \unit_memory/DRAM/n240 ,
         \unit_memory/DRAM/n239 , \unit_memory/DRAM/n238 ,
         \unit_memory/DRAM/n237 , \unit_memory/DRAM/n236 ,
         \unit_memory/DRAM/n235 , \unit_memory/DRAM/n234 ,
         \unit_memory/DRAM/n233 , \unit_memory/DRAM/n232 ,
         \unit_memory/DRAM/n231 , \unit_memory/DRAM/n230 ,
         \unit_memory/DRAM/n229 , \unit_memory/DRAM/n228 ,
         \unit_memory/DRAM/n227 , \unit_memory/DRAM/n226 ,
         \unit_memory/DRAM/n225 , \unit_memory/DRAM/n224 ,
         \unit_memory/DRAM/n223 , \unit_memory/DRAM/n222 ,
         \unit_memory/DRAM/n221 , \unit_memory/DRAM/n220 ,
         \unit_memory/DRAM/n219 , \unit_memory/DRAM/n218 ,
         \unit_memory/DRAM/n217 , \unit_memory/DRAM/n216 ,
         \unit_memory/DRAM/n215 , \unit_memory/DRAM/n214 ,
         \unit_memory/DRAM/n213 , \unit_memory/DRAM/n212 ,
         \unit_memory/DRAM/n211 , \unit_memory/DRAM/n210 ,
         \unit_memory/DRAM/n209 , \unit_memory/DRAM/n208 ,
         \unit_memory/DRAM/n207 , \unit_memory/DRAM/n206 ,
         \unit_memory/DRAM/n205 , \unit_memory/DRAM/n204 ,
         \unit_memory/DRAM/n203 , \unit_memory/DRAM/n202 ,
         \unit_memory/DRAM/n201 , \unit_memory/DRAM/n200 ,
         \unit_memory/DRAM/n199 , \unit_memory/DRAM/n198 ,
         \unit_memory/DRAM/n197 , \unit_memory/DRAM/n196 ,
         \unit_memory/DRAM/n195 , \unit_memory/DRAM/n194 ,
         \unit_memory/DRAM/n193 , \unit_memory/DRAM/n192 ,
         \unit_memory/DRAM/n191 , \unit_memory/DRAM/n190 ,
         \unit_memory/DRAM/n189 , \unit_memory/DRAM/n188 ,
         \unit_memory/DRAM/n187 , \unit_memory/DRAM/n186 ,
         \unit_memory/DRAM/n185 , \unit_memory/DRAM/n184 ,
         \unit_memory/DRAM/n183 , \unit_memory/DRAM/n182 ,
         \unit_memory/DRAM/n181 , \unit_memory/DRAM/n180 ,
         \unit_memory/DRAM/n179 , \unit_memory/DRAM/n178 ,
         \unit_memory/DRAM/n177 , \unit_memory/DRAM/n176 ,
         \unit_memory/DRAM/n175 , \unit_memory/DRAM/n174 ,
         \unit_memory/DRAM/n173 , \unit_memory/DRAM/n172 ,
         \unit_memory/DRAM/n171 , \unit_memory/DRAM/n170 ,
         \unit_memory/DRAM/n169 , \unit_memory/DRAM/n168 ,
         \unit_memory/DRAM/n167 , \unit_memory/DRAM/n166 ,
         \unit_memory/DRAM/n165 , \unit_memory/DRAM/n164 ,
         \unit_memory/DRAM/n163 , \unit_memory/DRAM/n162 ,
         \unit_memory/DRAM/n161 , \unit_memory/DRAM/n160 ,
         \unit_memory/DRAM/n159 , \unit_memory/DRAM/n158 ,
         \unit_memory/DRAM/n157 , \unit_memory/DRAM/n156 ,
         \unit_memory/DRAM/n155 , \unit_memory/DRAM/n154 ,
         \unit_memory/DRAM/n153 , \unit_memory/DRAM/n152 ,
         \unit_memory/DRAM/n151 , \unit_memory/DRAM/n150 ,
         \unit_memory/DRAM/n149 , \unit_memory/DRAM/n148 ,
         \unit_memory/DRAM/n147 , \unit_memory/DRAM/n146 ,
         \unit_memory/DRAM/n145 , \unit_memory/DRAM/n144 ,
         \unit_memory/DRAM/n143 , \unit_memory/DRAM/n142 ,
         \unit_memory/DRAM/n141 , \unit_memory/DRAM/n140 ,
         \unit_memory/DRAM/n139 , \unit_memory/DRAM/n138 ,
         \unit_memory/DRAM/n137 , \unit_memory/DRAM/n136 ,
         \unit_memory/DRAM/n135 , \unit_memory/DRAM/n134 ,
         \unit_memory/DRAM/n133 , \unit_memory/DRAM/n132 ,
         \unit_memory/DRAM/n131 , \unit_memory/DRAM/n130 ,
         \unit_memory/DRAM/n129 , \unit_memory/DRAM/n128 ,
         \unit_memory/DRAM/n127 , \unit_memory/DRAM/n126 ,
         \unit_memory/DRAM/n125 , \unit_memory/DRAM/n124 ,
         \unit_memory/DRAM/n123 , \unit_memory/DRAM/n122 ,
         \unit_memory/DRAM/n121 , \unit_memory/DRAM/n120 ,
         \unit_memory/DRAM/n119 , \unit_memory/DRAM/n118 ,
         \unit_memory/DRAM/n117 , \unit_memory/DRAM/n116 ,
         \unit_memory/DRAM/n115 , \unit_memory/DRAM/n114 ,
         \unit_memory/DRAM/n113 , \unit_memory/DRAM/n112 ,
         \unit_memory/DRAM/n111 , \unit_memory/DRAM/n110 ,
         \unit_memory/DRAM/n109 , \unit_memory/DRAM/n108 ,
         \unit_memory/DRAM/n107 , \unit_memory/DRAM/n106 ,
         \unit_memory/DRAM/n105 , \unit_memory/DRAM/n104 ,
         \unit_memory/DRAM/n103 , \unit_memory/DRAM/n102 ,
         \unit_memory/DRAM/n101 , \unit_memory/DRAM/n100 ,
         \unit_memory/DRAM/n99 , \unit_memory/DRAM/n98 ,
         \unit_memory/DRAM/n97 , \unit_memory/DRAM/n96 ,
         \unit_memory/DRAM/n95 , \unit_memory/DRAM/n94 ,
         \unit_memory/DRAM/n93 , \unit_memory/DRAM/n92 ,
         \unit_memory/DRAM/n91 , \unit_memory/DRAM/n90 ,
         \unit_memory/DRAM/n89 , \unit_memory/DRAM/n88 ,
         \unit_memory/DRAM/n87 , \unit_memory/DRAM/n86 ,
         \unit_memory/DRAM/n85 , \unit_memory/DRAM/n84 ,
         \unit_memory/DRAM/n83 , \unit_memory/DRAM/n82 ,
         \unit_memory/DRAM/n81 , \unit_memory/DRAM/n80 ,
         \unit_memory/DRAM/n79 , \unit_memory/DRAM/n78 ,
         \unit_memory/DRAM/n77 , \unit_memory/DRAM/n76 ,
         \unit_memory/DRAM/n75 , \unit_memory/DRAM/n74 ,
         \unit_memory/DRAM/n73 , \unit_memory/DRAM/n72 ,
         \unit_memory/DRAM/n71 , \unit_memory/DRAM/n70 ,
         \unit_memory/DRAM/n69 , \unit_memory/DRAM/n68 ,
         \unit_memory/DRAM/n67 , \unit_memory/DRAM/n66 ,
         \unit_memory/DRAM/n65 , \unit_memory/DRAM/n64 ,
         \unit_memory/DRAM/n63 , \unit_memory/DRAM/n62 ,
         \unit_memory/DRAM/n61 , \unit_memory/DRAM/n60 ,
         \unit_memory/DRAM/n59 , \unit_memory/DRAM/n58 ,
         \unit_memory/DRAM/n57 , \unit_memory/DRAM/n56 ,
         \unit_memory/DRAM/n55 , \unit_memory/DRAM/n54 ,
         \unit_memory/DRAM/n53 , \unit_memory/DRAM/n52 ,
         \unit_memory/DRAM/n51 , \unit_memory/DRAM/n50 ,
         \unit_memory/DRAM/n49 , \unit_memory/DRAM/n48 ,
         \unit_memory/DRAM/n47 , \unit_memory/DRAM/n46 ,
         \unit_memory/DRAM/n45 , \unit_memory/DRAM/n44 ,
         \unit_memory/DRAM/n43 , \unit_memory/DRAM/n42 ,
         \unit_memory/DRAM/n41 , \unit_memory/DRAM/n40 ,
         \unit_memory/DRAM/n39 , \unit_memory/DRAM/n38 ,
         \unit_memory/DRAM/n37 , \unit_memory/DRAM/n36 ,
         \unit_memory/DRAM/n35 , \unit_memory/DRAM/n34 ,
         \unit_memory/DRAM/n33 , \unit_memory/DRAM/n32 ,
         \unit_memory/DRAM/n31 , \unit_memory/DRAM/n30 ,
         \unit_memory/DRAM/n29 , \unit_memory/DRAM/n28 ,
         \unit_memory/DRAM/n27 , \unit_memory/DRAM/n26 ,
         \unit_memory/DRAM/n25 , \unit_memory/DRAM/n24 ,
         \unit_memory/DRAM/n23 , \unit_memory/DRAM/n22 ,
         \unit_memory/DRAM/n21 , \unit_memory/DRAM/n20 ,
         \unit_memory/DRAM/n19 , \unit_memory/DRAM/n18 ,
         \unit_memory/DRAM/n17 , \unit_memory/DRAM/n16 ,
         \unit_memory/DRAM/n15 , \unit_memory/DRAM/n14 ,
         \unit_memory/DRAM/n13 , \unit_memory/DRAM/n12 ,
         \unit_memory/DRAM/n11 , \unit_memory/DRAM/n10 , \unit_memory/DRAM/n9 ,
         \unit_memory/DRAM/n8 , \unit_memory/DRAM/n7 , \unit_memory/DRAM/n6 ,
         \unit_memory/DRAM/n5 , \unit_memory/DRAM/n4 , \unit_memory/DRAM/n3 ,
         \unit_memory/DRAM/n2 , \unit_memory/DRAM/n1 ,
         \unit_memory/DRAM/n2180 , \unit_memory/DRAM/n2179 ,
         \unit_memory/DRAM/n2178 , \unit_memory/DRAM/n2177 ,
         \unit_memory/DRAM/n2176 , \unit_memory/DRAM/n2175 ,
         \unit_memory/DRAM/n2174 , \unit_memory/DRAM/n2173 ,
         \unit_memory/DRAM/n2172 , \unit_memory/DRAM/n2171 ,
         \unit_memory/DRAM/n2170 , \unit_memory/DRAM/n2169 ,
         \unit_memory/DRAM/n2168 , \unit_memory/DRAM/n2167 ,
         \unit_memory/DRAM/n2166 , \unit_memory/DRAM/n2165 ,
         \unit_memory/DRAM/n2164 , \unit_memory/DRAM/n2163 ,
         \unit_memory/DRAM/n2162 , \unit_memory/DRAM/n2161 ,
         \unit_memory/DRAM/n2160 , \unit_memory/DRAM/n2159 ,
         \unit_memory/DRAM/n2158 , \unit_memory/DRAM/n2157 ,
         \unit_memory/DRAM/n2156 , \unit_memory/DRAM/n2155 ,
         \unit_memory/DRAM/n2154 , \unit_memory/DRAM/n2153 ,
         \unit_memory/DRAM/n2152 , \unit_memory/DRAM/n2151 ,
         \unit_memory/DRAM/n2150 , \unit_memory/DRAM/n2149 ,
         \unit_memory/DRAM/n2148 , \unit_memory/DRAM/n2147 ,
         \unit_memory/DRAM/n2146 , \unit_memory/DRAM/n2145 ,
         \unit_memory/DRAM/n2144 , \unit_memory/DRAM/n2143 ,
         \unit_memory/DRAM/n2142 , \unit_memory/DRAM/n2141 ,
         \unit_memory/DRAM/n2140 , \unit_memory/DRAM/n2139 ,
         \unit_memory/DRAM/n2138 , \unit_memory/DRAM/n2137 ,
         \unit_memory/DRAM/n2136 , \unit_memory/DRAM/n2135 ,
         \unit_memory/DRAM/n2134 , \unit_memory/DRAM/n2133 ,
         \unit_memory/DRAM/n2132 , \unit_memory/DRAM/n2131 ,
         \unit_memory/DRAM/n2130 , \unit_memory/DRAM/n2129 ,
         \unit_memory/DRAM/n2128 , \unit_memory/DRAM/n2127 ,
         \unit_memory/DRAM/n2126 , \unit_memory/DRAM/n2125 ,
         \unit_memory/DRAM/n2124 , \unit_memory/DRAM/n2123 ,
         \unit_memory/DRAM/n2122 , \unit_memory/DRAM/n2121 ,
         \unit_memory/DRAM/n2120 , \unit_memory/DRAM/n2119 ,
         \unit_memory/DRAM/n2118 , \unit_memory/DRAM/n2117 ,
         \unit_memory/DRAM/n2116 , \unit_memory/DRAM/n2115 ,
         \unit_memory/DRAM/n2114 , \unit_memory/DRAM/n2113 ,
         \unit_memory/DRAM/n2112 , \unit_memory/DRAM/n2111 ,
         \unit_memory/DRAM/n2110 , \unit_memory/DRAM/n2109 ,
         \unit_memory/DRAM/n2108 , \unit_memory/DRAM/n2107 ,
         \unit_memory/DRAM/n2106 , \unit_memory/DRAM/n2105 ,
         \unit_memory/DRAM/n2104 , \unit_memory/DRAM/n2103 ,
         \unit_memory/DRAM/n2102 , \unit_memory/DRAM/n2101 ,
         \unit_memory/DRAM/n2100 , \unit_memory/DRAM/n2099 ,
         \unit_memory/DRAM/n2098 , \unit_memory/DRAM/n2097 ,
         \unit_memory/DRAM/n2096 , \unit_memory/DRAM/n2095 ,
         \unit_memory/DRAM/n2094 , \unit_memory/DRAM/n2093 ,
         \unit_memory/DRAM/n2092 , \unit_memory/DRAM/n2091 ,
         \unit_memory/DRAM/n2090 , \unit_memory/DRAM/n2089 ,
         \unit_memory/DRAM/n2088 , \unit_memory/DRAM/n2087 ,
         \unit_memory/DRAM/n2086 , \unit_memory/DRAM/n2085 ,
         \unit_memory/DRAM/n2084 , \unit_memory/DRAM/n2083 ,
         \unit_memory/DRAM/n2082 , \unit_memory/DRAM/n2081 ,
         \unit_memory/DRAM/n2080 , \unit_memory/DRAM/n2079 ,
         \unit_memory/DRAM/n2078 , \unit_memory/DRAM/n2077 ,
         \unit_memory/DRAM/n2076 , \unit_memory/DRAM/n2075 ,
         \unit_memory/DRAM/n2074 , \unit_memory/DRAM/n2073 ,
         \unit_memory/DRAM/n2072 , \unit_memory/DRAM/n2071 ,
         \unit_memory/DRAM/n2070 , \unit_memory/DRAM/n2069 ,
         \unit_memory/DRAM/n2068 , \unit_memory/DRAM/n2067 ,
         \unit_memory/DRAM/n2066 , \unit_memory/DRAM/n2065 ,
         \unit_memory/DRAM/n2064 , \unit_memory/DRAM/n2063 ,
         \unit_memory/DRAM/n2062 , \unit_memory/DRAM/n2061 ,
         \unit_memory/DRAM/n2060 , \unit_memory/DRAM/n2059 ,
         \unit_memory/DRAM/n2058 , \unit_memory/DRAM/n2057 ,
         \unit_memory/DRAM/n2056 , \unit_memory/DRAM/n2055 ,
         \unit_memory/DRAM/n2054 , \unit_memory/DRAM/n2053 ,
         \unit_memory/DRAM/n2052 , \unit_memory/DRAM/n2051 ,
         \unit_memory/DRAM/n2050 , \unit_memory/DRAM/n2049 ,
         \unit_memory/DRAM/n2048 , \unit_memory/DRAM/n2047 ,
         \unit_memory/DRAM/n2046 , \unit_memory/DRAM/n2045 ,
         \unit_memory/DRAM/n2044 , \unit_memory/DRAM/n2043 ,
         \unit_memory/DRAM/n2042 , \unit_memory/DRAM/n2041 ,
         \unit_memory/DRAM/n2040 , \unit_memory/DRAM/n2039 ,
         \unit_memory/DRAM/n2038 , \unit_memory/DRAM/n2037 ,
         \unit_memory/DRAM/n2036 , \unit_memory/DRAM/n2035 ,
         \unit_memory/DRAM/n2034 , \unit_memory/DRAM/n2033 ,
         \unit_memory/DRAM/n2032 , \unit_memory/DRAM/n2031 ,
         \unit_memory/DRAM/n2030 , \unit_memory/DRAM/n2029 ,
         \unit_memory/DRAM/n2028 , \unit_memory/DRAM/n2027 ,
         \unit_memory/DRAM/n2026 , \unit_memory/DRAM/n2025 ,
         \unit_memory/DRAM/n2024 , \unit_memory/DRAM/n2023 ,
         \unit_memory/DRAM/n2022 , \unit_memory/DRAM/n2021 ,
         \unit_memory/DRAM/n2020 , \unit_memory/DRAM/n2019 ,
         \unit_memory/DRAM/n2018 , \unit_memory/DRAM/n2017 ,
         \unit_memory/DRAM/n2016 , \unit_memory/DRAM/n2015 ,
         \unit_memory/DRAM/n2014 , \unit_memory/DRAM/n2013 ,
         \unit_memory/DRAM/n2012 , \unit_memory/DRAM/n2011 ,
         \unit_memory/DRAM/n2010 , \unit_memory/DRAM/n2009 ,
         \unit_memory/DRAM/n2008 , \unit_memory/DRAM/n2007 ,
         \unit_memory/DRAM/n2006 , \unit_memory/DRAM/n2005 ,
         \unit_memory/DRAM/n2004 , \unit_memory/DRAM/n2003 ,
         \unit_memory/DRAM/n2002 , \unit_memory/DRAM/n2001 ,
         \unit_memory/DRAM/n2000 , \unit_memory/DRAM/n1999 ,
         \unit_memory/DRAM/n1998 , \unit_memory/DRAM/n1997 ,
         \unit_memory/DRAM/n1996 , \unit_memory/DRAM/n1995 ,
         \unit_memory/DRAM/n1994 , \unit_memory/DRAM/n1993 ,
         \unit_memory/DRAM/n1992 , \unit_memory/DRAM/n1991 ,
         \unit_memory/DRAM/n1990 , \unit_memory/DRAM/n1989 ,
         \unit_memory/DRAM/n1988 , \unit_memory/DRAM/n1987 ,
         \unit_memory/DRAM/n1986 , \unit_memory/DRAM/n1985 ,
         \unit_memory/DRAM/n1984 , \unit_memory/DRAM/n1983 ,
         \unit_memory/DRAM/n1982 , \unit_memory/DRAM/n1981 ,
         \unit_memory/DRAM/n1980 , \unit_memory/DRAM/n1979 ,
         \unit_memory/DRAM/n1978 , \unit_memory/DRAM/n1977 ,
         \unit_memory/DRAM/n1976 , \unit_memory/DRAM/n1975 ,
         \unit_memory/DRAM/n1974 , \unit_memory/DRAM/n1973 ,
         \unit_memory/DRAM/n1972 , \unit_memory/DRAM/n1971 ,
         \unit_memory/DRAM/n1970 , \unit_memory/DRAM/n1969 ,
         \unit_memory/DRAM/n1968 , \unit_memory/DRAM/n1967 ,
         \unit_memory/DRAM/n1966 , \unit_memory/DRAM/n1965 ,
         \unit_memory/DRAM/n1964 , \unit_memory/DRAM/n1963 ,
         \unit_memory/DRAM/n1962 , \unit_memory/DRAM/n1961 ,
         \unit_memory/DRAM/n1960 , \unit_memory/DRAM/n1959 ,
         \unit_memory/DRAM/n1958 , \unit_memory/DRAM/n1957 ,
         \unit_memory/DRAM/n1956 , \unit_memory/DRAM/n1955 ,
         \unit_memory/DRAM/n1954 , \unit_memory/DRAM/n1953 ,
         \unit_memory/DRAM/n1952 , \unit_memory/DRAM/n1951 ,
         \unit_memory/DRAM/n1950 , \unit_memory/DRAM/n1949 ,
         \unit_memory/DRAM/n1948 , \unit_memory/DRAM/n1947 ,
         \unit_memory/DRAM/n1946 , \unit_memory/DRAM/n1945 ,
         \unit_memory/DRAM/n1944 , \unit_memory/DRAM/n1943 ,
         \unit_memory/DRAM/n1942 , \unit_memory/DRAM/n1941 ,
         \unit_memory/DRAM/n1940 , \unit_memory/DRAM/n1939 ,
         \unit_memory/DRAM/n1938 , \unit_memory/DRAM/n1937 ,
         \unit_memory/DRAM/n1936 , \unit_memory/DRAM/n1935 ,
         \unit_memory/DRAM/n1934 , \unit_memory/DRAM/n1933 ,
         \unit_memory/DRAM/n1932 , \unit_memory/DRAM/n1931 ,
         \unit_memory/DRAM/n1930 , \unit_memory/DRAM/n1929 ,
         \unit_memory/DRAM/n1928 , \unit_memory/DRAM/n1927 ,
         \unit_memory/DRAM/n1926 , \unit_memory/DRAM/n1925 ,
         \unit_memory/DRAM/n1924 , \unit_memory/DRAM/n1923 ,
         \unit_memory/DRAM/n1922 , \unit_memory/DRAM/n1921 ,
         \unit_memory/DRAM/n1920 , \unit_memory/DRAM/n1919 ,
         \unit_memory/DRAM/n1918 , \unit_memory/DRAM/n1917 ,
         \unit_memory/DRAM/n1916 , \unit_memory/DRAM/n1915 ,
         \unit_memory/DRAM/n1914 , \unit_memory/DRAM/n1913 ,
         \unit_memory/DRAM/n1912 , \unit_memory/DRAM/n1911 ,
         \unit_memory/DRAM/n1910 , \unit_memory/DRAM/n1909 ,
         \unit_memory/DRAM/n1908 , \unit_memory/DRAM/n1907 ,
         \unit_memory/DRAM/n1906 , \unit_memory/DRAM/n1905 ,
         \unit_memory/DRAM/n1904 , \unit_memory/DRAM/n1903 ,
         \unit_memory/DRAM/n1902 , \unit_memory/DRAM/n1901 ,
         \unit_memory/DRAM/n1900 , \unit_memory/DRAM/n1899 ,
         \unit_memory/DRAM/n1898 , \unit_memory/DRAM/n1897 ,
         \unit_memory/DRAM/n1896 , \unit_memory/DRAM/n1895 ,
         \unit_memory/DRAM/n1894 , \unit_memory/DRAM/n1893 ,
         \unit_memory/DRAM/n1892 , \unit_memory/DRAM/n1891 ,
         \unit_memory/DRAM/n1890 , \unit_memory/DRAM/n1889 ,
         \unit_memory/DRAM/n1888 , \unit_memory/DRAM/n1887 ,
         \unit_memory/DRAM/n1886 , \unit_memory/DRAM/n1885 ,
         \unit_memory/DRAM/n1884 , \unit_memory/DRAM/n1883 ,
         \unit_memory/DRAM/n1882 , \unit_memory/DRAM/n1881 ,
         \unit_memory/DRAM/n1880 , \unit_memory/DRAM/n1879 ,
         \unit_memory/DRAM/n1878 , \unit_memory/DRAM/n1877 ,
         \unit_memory/DRAM/n1876 , \unit_memory/DRAM/n1875 ,
         \unit_memory/DRAM/n1874 , \unit_memory/DRAM/n1873 ,
         \unit_memory/DRAM/n1872 , \unit_memory/DRAM/n1871 ,
         \unit_memory/DRAM/n1870 , \unit_memory/DRAM/n1869 ,
         \unit_memory/DRAM/n1868 , \unit_memory/DRAM/n1867 ,
         \unit_memory/DRAM/n1866 , \unit_memory/DRAM/n1865 ,
         \unit_memory/DRAM/n1864 , \unit_memory/DRAM/n1863 ,
         \unit_memory/DRAM/n1862 , \unit_memory/DRAM/n1861 ,
         \unit_memory/DRAM/n1860 , \unit_memory/DRAM/n1859 ,
         \unit_memory/DRAM/n1858 , \unit_memory/DRAM/n1857 ,
         \unit_memory/DRAM/n1856 , \unit_memory/DRAM/n1855 ,
         \unit_memory/DRAM/n1854 , \unit_memory/DRAM/n1853 ,
         \unit_memory/DRAM/n1852 , \unit_memory/DRAM/n1851 ,
         \unit_memory/DRAM/n1850 , \unit_memory/DRAM/n1849 ,
         \unit_memory/DRAM/n1848 , \unit_memory/DRAM/n1847 ,
         \unit_memory/DRAM/n1846 , \unit_memory/DRAM/n1845 ,
         \unit_memory/DRAM/n1844 , \unit_memory/DRAM/n1843 ,
         \unit_memory/DRAM/n1842 , \unit_memory/DRAM/n1841 ,
         \unit_memory/DRAM/n1840 , \unit_memory/DRAM/n1839 ,
         \unit_memory/DRAM/n1838 , \unit_memory/DRAM/n1837 ,
         \unit_memory/DRAM/n1836 , \unit_memory/DRAM/n1835 ,
         \unit_memory/DRAM/n1834 , \unit_memory/DRAM/n1833 ,
         \unit_memory/DRAM/n1832 , \unit_memory/DRAM/n1831 ,
         \unit_memory/DRAM/n1830 , \unit_memory/DRAM/n1829 ,
         \unit_memory/DRAM/n1828 , \unit_memory/DRAM/n1827 ,
         \unit_memory/DRAM/n1826 , \unit_memory/DRAM/n1825 ,
         \unit_memory/DRAM/n1824 , \unit_memory/DRAM/n1823 ,
         \unit_memory/DRAM/n1822 , \unit_memory/DRAM/n1821 ,
         \unit_memory/DRAM/n1820 , \unit_memory/DRAM/n1819 ,
         \unit_memory/DRAM/n1818 , \unit_memory/DRAM/n1817 ,
         \unit_memory/DRAM/n1816 , \unit_memory/DRAM/n1815 ,
         \unit_memory/DRAM/n1814 , \unit_memory/DRAM/n1813 ,
         \unit_memory/DRAM/n1812 , \unit_memory/DRAM/n1811 ,
         \unit_memory/DRAM/n1810 , \unit_memory/DRAM/n1809 ,
         \unit_memory/DRAM/n1808 , \unit_memory/DRAM/n1807 ,
         \unit_memory/DRAM/n1806 , \unit_memory/DRAM/n1805 ,
         \unit_memory/DRAM/n1804 , \unit_memory/DRAM/n1803 ,
         \unit_memory/DRAM/n1802 , \unit_memory/DRAM/n1801 ,
         \unit_memory/DRAM/n1800 , \unit_memory/DRAM/n1799 ,
         \unit_memory/DRAM/n1798 , \unit_memory/DRAM/n1797 ,
         \unit_memory/DRAM/n1796 , \unit_memory/DRAM/n1795 ,
         \unit_memory/DRAM/n1794 , \unit_memory/DRAM/n1793 ,
         \unit_memory/DRAM/n1792 , \unit_memory/DRAM/n1791 ,
         \unit_memory/DRAM/n1790 , \unit_memory/DRAM/n1789 ,
         \unit_memory/DRAM/n1788 , \unit_memory/DRAM/n1787 ,
         \unit_memory/DRAM/n1786 , \unit_memory/DRAM/n1785 ,
         \unit_memory/DRAM/n1784 , \unit_memory/DRAM/n1783 ,
         \unit_memory/DRAM/n1782 , \unit_memory/DRAM/n1781 ,
         \unit_memory/DRAM/n1780 , \unit_memory/DRAM/n1779 ,
         \unit_memory/DRAM/n1778 , \unit_memory/DRAM/n1777 ,
         \unit_memory/DRAM/n1776 , \unit_memory/DRAM/n1775 ,
         \unit_memory/DRAM/n1774 , \unit_memory/DRAM/n1773 ,
         \unit_memory/DRAM/n1772 , \unit_memory/DRAM/n1771 ,
         \unit_memory/DRAM/n1770 , \unit_memory/DRAM/n1769 ,
         \unit_memory/DRAM/n1768 , \unit_memory/DRAM/n1767 ,
         \unit_memory/DRAM/n1766 , \unit_memory/DRAM/n1765 ,
         \unit_memory/DRAM/n1764 , \unit_memory/DRAM/n1763 ,
         \unit_memory/DRAM/n1762 , \unit_memory/DRAM/n1761 ,
         \unit_memory/DRAM/n1760 , \unit_memory/DRAM/n1759 ,
         \unit_memory/DRAM/n1758 , \unit_memory/DRAM/n1757 ,
         \unit_memory/DRAM/n1756 , \unit_memory/DRAM/n1755 ,
         \unit_memory/DRAM/n1754 , \unit_memory/DRAM/n1753 ,
         \unit_memory/DRAM/n1752 , \unit_memory/DRAM/n1751 ,
         \unit_memory/DRAM/n1750 , \unit_memory/DRAM/n1749 ,
         \unit_memory/DRAM/n1748 , \unit_memory/DRAM/n1747 ,
         \unit_memory/DRAM/n1746 , \unit_memory/DRAM/n1745 ,
         \unit_memory/DRAM/n1744 , \unit_memory/DRAM/n1743 ,
         \unit_memory/DRAM/n1742 , \unit_memory/DRAM/n1741 ,
         \unit_memory/DRAM/n1740 , \unit_memory/DRAM/n1739 ,
         \unit_memory/DRAM/n1738 , \unit_memory/DRAM/n1737 ,
         \unit_memory/DRAM/n1736 , \unit_memory/DRAM/n1735 ,
         \unit_memory/DRAM/n1734 , \unit_memory/DRAM/n1733 ,
         \unit_memory/DRAM/n1732 , \unit_memory/DRAM/n1731 ,
         \unit_memory/DRAM/n1730 , \unit_memory/DRAM/n1729 ,
         \unit_memory/DRAM/n1728 , \unit_memory/DRAM/n1727 ,
         \unit_memory/DRAM/n1726 , \unit_memory/DRAM/n1725 ,
         \unit_memory/DRAM/n1724 , \unit_memory/DRAM/n1723 ,
         \unit_memory/DRAM/n1722 , \unit_memory/DRAM/n1721 ,
         \unit_memory/DRAM/n1720 , \unit_memory/DRAM/n1719 ,
         \unit_memory/DRAM/n1718 , \unit_memory/DRAM/n1717 ,
         \unit_memory/DRAM/n1716 , \unit_memory/DRAM/n1715 ,
         \unit_memory/DRAM/n1714 , \unit_memory/DRAM/n1713 ,
         \unit_memory/DRAM/n1712 , \unit_memory/DRAM/n1711 ,
         \unit_memory/DRAM/n1710 , \unit_memory/DRAM/n1709 ,
         \unit_memory/DRAM/n1708 , \unit_memory/DRAM/n1707 ,
         \unit_memory/DRAM/n1706 , \unit_memory/DRAM/n1705 ,
         \unit_memory/DRAM/n1704 , \unit_memory/DRAM/n1703 ,
         \unit_memory/DRAM/n1702 , \unit_memory/DRAM/n1701 ,
         \unit_memory/DRAM/n1700 , \unit_memory/DRAM/n1699 ,
         \unit_memory/DRAM/n1698 , \unit_memory/DRAM/n1697 ,
         \unit_memory/DRAM/n1696 , \unit_memory/DRAM/n1695 ,
         \unit_memory/DRAM/n1694 , \unit_memory/DRAM/n1693 ,
         \unit_memory/DRAM/n1692 , \unit_memory/DRAM/n1691 ,
         \unit_memory/DRAM/n1690 , \unit_memory/DRAM/n1689 ,
         \unit_memory/DRAM/n1688 , \unit_memory/DRAM/n1687 ,
         \unit_memory/DRAM/n1686 , \unit_memory/DRAM/n1685 ,
         \unit_memory/DRAM/n1684 , \unit_memory/DRAM/n1683 ,
         \unit_memory/DRAM/n1682 , \unit_memory/DRAM/n1681 ,
         \unit_memory/DRAM/n1680 , \unit_memory/DRAM/n1679 ,
         \unit_memory/DRAM/n1678 , \unit_memory/DRAM/n1677 ,
         \unit_memory/DRAM/n1676 , \unit_memory/DRAM/n1675 ,
         \unit_memory/DRAM/n1674 , \unit_memory/DRAM/n1673 ,
         \unit_memory/DRAM/n1672 , \unit_memory/DRAM/n1671 ,
         \unit_memory/DRAM/n1670 , \unit_memory/DRAM/n1669 ,
         \unit_memory/DRAM/n1668 , \unit_memory/DRAM/n1667 ,
         \unit_memory/DRAM/n1666 , \unit_memory/DRAM/n1665 ,
         \unit_memory/DRAM/n1664 , \unit_memory/DRAM/n1663 ,
         \unit_memory/DRAM/n1662 , \unit_memory/DRAM/n1661 ,
         \unit_memory/DRAM/n1660 , \unit_memory/DRAM/n1659 ,
         \unit_memory/DRAM/n1658 , \unit_memory/DRAM/n1657 ,
         \unit_memory/DRAM/n1656 , \unit_memory/DRAM/n1655 ,
         \unit_memory/DRAM/n1654 , \unit_memory/DRAM/n1653 ,
         \unit_memory/DRAM/n1652 , \unit_memory/DRAM/n1651 ,
         \unit_memory/DRAM/n1650 , \unit_memory/DRAM/n1649 ,
         \unit_memory/DRAM/n1648 , \unit_memory/DRAM/n1647 ,
         \unit_memory/DRAM/n1646 , \unit_memory/DRAM/n1645 ,
         \unit_memory/DRAM/n1644 , \unit_memory/DRAM/n1643 ,
         \unit_memory/DRAM/n1642 , \unit_memory/DRAM/n1641 ,
         \unit_memory/DRAM/n1640 , \unit_memory/DRAM/n1639 ,
         \unit_memory/DRAM/n1638 , \unit_memory/DRAM/n1637 ,
         \unit_memory/DRAM/n1636 , \unit_memory/DRAM/n1635 ,
         \unit_memory/DRAM/n1634 , \unit_memory/DRAM/n1633 ,
         \unit_memory/DRAM/n1632 , \unit_memory/DRAM/n1631 ,
         \unit_memory/DRAM/n1630 , \unit_memory/DRAM/n1629 ,
         \unit_memory/DRAM/n1628 , \unit_memory/DRAM/n1627 ,
         \unit_memory/DRAM/n1626 , \unit_memory/DRAM/n1625 ,
         \unit_memory/DRAM/n1624 , \unit_memory/DRAM/n1623 ,
         \unit_memory/DRAM/n1622 , \unit_memory/DRAM/n1621 ,
         \unit_memory/DRAM/n1620 , \unit_memory/DRAM/n1619 ,
         \unit_memory/DRAM/n1618 , \unit_memory/DRAM/n1617 ,
         \unit_memory/DRAM/n1616 , \unit_memory/DRAM/n1615 ,
         \unit_memory/DRAM/n1614 , \unit_memory/DRAM/n1613 ,
         \unit_memory/DRAM/n1612 , \unit_memory/DRAM/n1611 ,
         \unit_memory/DRAM/n1610 , \unit_memory/DRAM/n1609 ,
         \unit_memory/DRAM/n1608 , \unit_memory/DRAM/n1607 ,
         \unit_memory/DRAM/n1606 , \unit_memory/DRAM/n1605 ,
         \unit_memory/DRAM/n1604 , \unit_memory/DRAM/n1603 ,
         \unit_memory/DRAM/n1602 , \unit_memory/DRAM/n1601 ,
         \unit_memory/DRAM/n1600 , \unit_memory/DRAM/n1599 ,
         \unit_memory/DRAM/n1598 , \unit_memory/DRAM/n1597 ,
         \unit_memory/DRAM/n1596 , \unit_memory/DRAM/n1595 ,
         \unit_memory/DRAM/n1594 , \unit_memory/DRAM/n1593 ,
         \unit_memory/DRAM/n1592 , \unit_memory/DRAM/n1591 ,
         \unit_memory/DRAM/n1590 , \unit_memory/DRAM/n1589 ,
         \unit_memory/DRAM/n1588 , \unit_memory/DRAM/n1587 ,
         \unit_memory/DRAM/n1586 , \unit_memory/DRAM/n1585 ,
         \unit_memory/DRAM/n1584 , \unit_memory/DRAM/n1583 ,
         \unit_memory/DRAM/n1582 , \unit_memory/DRAM/n1581 ,
         \unit_memory/DRAM/n1580 , \unit_memory/DRAM/n1579 ,
         \unit_memory/DRAM/n1578 , \unit_memory/DRAM/n1577 ,
         \unit_memory/DRAM/n1576 , \unit_memory/DRAM/n1575 ,
         \unit_memory/DRAM/n1574 , \unit_memory/DRAM/n1573 ,
         \unit_memory/DRAM/n1572 , \unit_memory/DRAM/n1571 ,
         \unit_memory/DRAM/n1570 , \unit_memory/DRAM/n1569 ,
         \unit_memory/DRAM/n1568 , \unit_memory/DRAM/n1567 ,
         \unit_memory/DRAM/n1566 , \unit_memory/DRAM/n1565 ,
         \unit_memory/DRAM/n1564 , \unit_memory/DRAM/n1563 ,
         \unit_memory/DRAM/n1562 , \unit_memory/DRAM/n1561 ,
         \unit_memory/DRAM/n1560 , \unit_memory/DRAM/n1559 ,
         \unit_memory/DRAM/n1558 , \unit_memory/DRAM/n1557 ,
         \unit_memory/DRAM/n1556 , \unit_memory/DRAM/n1555 ,
         \unit_memory/DRAM/n1554 , \unit_memory/DRAM/n1553 ,
         \unit_memory/DRAM/n1552 , \unit_memory/DRAM/n1551 ,
         \unit_memory/DRAM/n1550 , \unit_memory/DRAM/n1549 ,
         \unit_memory/DRAM/n1548 , \unit_memory/DRAM/n1547 ,
         \unit_memory/DRAM/n1546 , \unit_memory/DRAM/n1545 ,
         \unit_memory/DRAM/n1544 , \unit_memory/DRAM/n1543 ,
         \unit_memory/DRAM/n1542 , \unit_memory/DRAM/n1541 ,
         \unit_memory/DRAM/n1540 , \unit_memory/DRAM/n1539 ,
         \unit_memory/DRAM/n1538 , \unit_memory/DRAM/n1537 ,
         \unit_memory/DRAM/n1536 , \unit_memory/DRAM/n1535 ,
         \unit_memory/DRAM/n1534 , \unit_memory/DRAM/n1533 ,
         \unit_memory/DRAM/n1532 , \unit_memory/DRAM/n1531 ,
         \unit_memory/DRAM/n1530 , \unit_memory/DRAM/n1529 ,
         \unit_memory/DRAM/n1528 , \unit_memory/DRAM/n1527 ,
         \unit_memory/DRAM/n1526 , \unit_memory/DRAM/n1525 ,
         \unit_memory/DRAM/n1524 , \unit_memory/DRAM/n1523 ,
         \unit_memory/DRAM/n1522 , \unit_memory/DRAM/n1521 ,
         \unit_memory/DRAM/n1520 , \unit_memory/DRAM/n1519 ,
         \unit_memory/DRAM/n1518 , \unit_memory/DRAM/n1517 ,
         \unit_memory/DRAM/n1516 , \unit_memory/DRAM/n1515 ,
         \unit_memory/DRAM/n1514 , \unit_memory/DRAM/n1513 ,
         \unit_memory/DRAM/n1512 , \unit_memory/DRAM/n1511 ,
         \unit_memory/DRAM/n1510 , \unit_memory/DRAM/n1509 ,
         \unit_memory/DRAM/n1508 , \unit_memory/DRAM/n1507 ,
         \unit_memory/DRAM/n1506 , \unit_memory/DRAM/n1505 ,
         \unit_memory/DRAM/n1504 , \unit_memory/DRAM/n1503 ,
         \unit_memory/DRAM/n1502 , \unit_memory/DRAM/n1501 ,
         \unit_memory/DRAM/n1500 , \unit_memory/DRAM/n1499 ,
         \unit_memory/DRAM/n1498 , \unit_memory/DRAM/n1497 ,
         \unit_memory/DRAM/n1496 , \unit_memory/DRAM/n1495 ,
         \unit_memory/DRAM/n1494 , \unit_memory/DRAM/n1493 ,
         \unit_memory/DRAM/n1492 , \unit_memory/DRAM/n1491 ,
         \unit_memory/DRAM/n1490 , \unit_memory/DRAM/n1489 ,
         \unit_memory/DRAM/n1488 , \unit_memory/DRAM/n1487 ,
         \unit_memory/DRAM/n1486 , \unit_memory/DRAM/n1485 ,
         \unit_memory/DRAM/n1484 , \unit_memory/DRAM/n1483 ,
         \unit_memory/DRAM/n1482 , \unit_memory/DRAM/n1481 ,
         \unit_memory/DRAM/n1480 , \unit_memory/DRAM/n1479 ,
         \unit_memory/DRAM/n1478 , \unit_memory/DRAM/n1477 ,
         \unit_memory/DRAM/n1476 , \unit_memory/DRAM/n1475 ,
         \unit_memory/DRAM/n1474 , \unit_memory/DRAM/n1473 ,
         \unit_memory/DRAM/n1472 , \unit_memory/DRAM/n1471 ,
         \unit_memory/DRAM/n1470 , \unit_memory/DRAM/n1469 ,
         \unit_memory/DRAM/n1468 , \unit_memory/DRAM/n1467 ,
         \unit_memory/DRAM/n1466 , \unit_memory/DRAM/n1465 ,
         \unit_memory/DRAM/n1464 , \unit_memory/DRAM/n1463 ,
         \unit_memory/DRAM/n1462 , \unit_memory/DRAM/n1461 ,
         \unit_memory/DRAM/n1460 , \unit_memory/DRAM/n1459 ,
         \unit_memory/DRAM/n1458 , \unit_memory/DRAM/n1457 ,
         \unit_memory/DRAM/n1456 , \unit_memory/DRAM/n1455 ,
         \unit_memory/DRAM/n1454 , \unit_memory/DRAM/n1453 ,
         \unit_memory/DRAM/n1452 , \unit_memory/DRAM/n1451 ,
         \unit_memory/DRAM/n1450 , \unit_memory/DRAM/n1449 ,
         \unit_memory/DRAM/n1448 , \unit_memory/DRAM/n1447 ,
         \unit_memory/DRAM/n1446 , \unit_memory/DRAM/n1445 ,
         \unit_memory/DRAM/n1444 , \unit_memory/DRAM/n1443 ,
         \unit_memory/DRAM/n1442 , \unit_memory/DRAM/n1441 ,
         \unit_memory/DRAM/n1440 , \unit_memory/DRAM/n1439 ,
         \unit_memory/DRAM/n1438 , \unit_memory/DRAM/n1437 ,
         \unit_memory/DRAM/n1436 , \unit_memory/DRAM/n1435 ,
         \unit_memory/DRAM/n1434 , \unit_memory/DRAM/n1433 ,
         \unit_memory/DRAM/n1432 , \unit_memory/DRAM/n1431 ,
         \unit_memory/DRAM/n1430 , \unit_memory/DRAM/n1429 ,
         \unit_memory/DRAM/n1428 , \unit_memory/DRAM/n1427 ,
         \unit_memory/DRAM/n1426 , \unit_memory/DRAM/n1425 ,
         \unit_memory/DRAM/n1424 , \unit_memory/DRAM/n1423 ,
         \unit_memory/DRAM/n1422 , \unit_memory/DRAM/n1421 ,
         \unit_memory/DRAM/n1420 , \unit_memory/DRAM/n1419 ,
         \unit_memory/DRAM/n1418 , \unit_memory/DRAM/n1417 ,
         \unit_memory/DRAM/n1416 , \unit_memory/DRAM/n1415 ,
         \unit_memory/DRAM/n1414 , \unit_memory/DRAM/n1413 ,
         \unit_memory/DRAM/n1412 , \unit_memory/DRAM/n1411 ,
         \unit_memory/DRAM/n1410 , \unit_memory/DRAM/n1409 ,
         \unit_memory/DRAM/n1408 , \unit_memory/DRAM/n1407 ,
         \unit_memory/DRAM/n1406 , \unit_memory/DRAM/n1405 ,
         \unit_memory/DRAM/n1404 , \unit_memory/DRAM/n1403 ,
         \unit_memory/DRAM/n1402 , \unit_memory/DRAM/n1401 ,
         \unit_memory/DRAM/n1400 , \unit_memory/DRAM/n1399 ,
         \unit_memory/DRAM/n1398 , \unit_memory/DRAM/n1397 ,
         \unit_memory/DRAM/n1396 , \unit_memory/DRAM/n1395 ,
         \unit_memory/DRAM/n1394 , \unit_memory/DRAM/n1393 ,
         \unit_memory/DRAM/n1392 , \unit_memory/DRAM/n1391 ,
         \unit_memory/DRAM/n1390 , \unit_memory/DRAM/n1389 ,
         \unit_memory/DRAM/n1388 , \unit_memory/DRAM/n1387 ,
         \unit_memory/DRAM/n1386 , \unit_memory/DRAM/n1385 ,
         \unit_memory/DRAM/n1384 , \unit_memory/DRAM/n1383 ,
         \unit_memory/DRAM/n1382 , \unit_memory/DRAM/n1381 ,
         \unit_memory/DRAM/n1380 , \unit_memory/DRAM/n1379 ,
         \unit_memory/DRAM/n1378 , \unit_memory/DRAM/n1377 ,
         \unit_memory/DRAM/n1376 , \unit_memory/DRAM/n1375 ,
         \unit_memory/DRAM/n1374 , \unit_memory/DRAM/n1373 ,
         \unit_memory/DRAM/n1372 , \unit_memory/DRAM/n1371 ,
         \unit_memory/DRAM/n1370 , \unit_memory/DRAM/n1369 ,
         \unit_memory/DRAM/n1368 , \unit_memory/DRAM/n1367 ,
         \unit_memory/DRAM/n1366 , \unit_memory/DRAM/n1365 ,
         \unit_memory/DRAM/n1364 , \unit_memory/DRAM/n1363 ,
         \unit_memory/DRAM/n1362 , \unit_memory/DRAM/n1361 ,
         \unit_memory/DRAM/n1360 , \unit_memory/DRAM/n1359 ,
         \unit_memory/DRAM/n1358 , \unit_memory/DRAM/n1357 ,
         \unit_memory/DRAM/n1356 , \unit_memory/DRAM/n1355 ,
         \unit_memory/DRAM/n1354 , \unit_memory/DRAM/n1353 ,
         \unit_memory/DRAM/n1352 , \unit_memory/DRAM/n1351 ,
         \unit_memory/DRAM/n1350 , \unit_memory/DRAM/n1349 ,
         \unit_memory/DRAM/n1348 , \unit_memory/DRAM/n1347 ,
         \unit_memory/DRAM/n1346 , \unit_memory/DRAM/n1345 ,
         \unit_memory/DRAM/n1344 , \unit_memory/DRAM/n1343 ,
         \unit_memory/DRAM/n1342 , \unit_memory/DRAM/n1341 ,
         \unit_memory/DRAM/n1340 , \unit_memory/DRAM/n1339 ,
         \unit_memory/DRAM/n1338 , \unit_memory/DRAM/n1337 ,
         \unit_memory/DRAM/n1336 , \unit_memory/DRAM/n1335 ,
         \unit_memory/DRAM/n1334 , \unit_memory/DRAM/n1333 ,
         \unit_memory/DRAM/n1332 , \unit_memory/DRAM/n1331 ,
         \unit_memory/DRAM/n1330 , \unit_memory/DRAM/n1329 ,
         \unit_memory/DRAM/n1328 , \unit_memory/DRAM/n1327 ,
         \unit_memory/DRAM/n1326 , \unit_memory/DRAM/n1325 ,
         \unit_memory/DRAM/n1324 , \unit_memory/DRAM/n1323 ,
         \unit_memory/DRAM/n1322 , \unit_memory/DRAM/n1321 ,
         \unit_memory/DRAM/n1320 , \unit_memory/DRAM/n1319 ,
         \unit_memory/DRAM/n1318 , \unit_memory/DRAM/n1317 ,
         \unit_memory/DRAM/n1316 , \unit_memory/DRAM/n1315 ,
         \unit_memory/DRAM/n1314 , \unit_memory/DRAM/n1313 ,
         \unit_memory/DRAM/n1312 , \unit_memory/DRAM/n1311 ,
         \unit_memory/DRAM/n1310 , \unit_memory/DRAM/n1309 ,
         \unit_memory/DRAM/n1308 , \unit_memory/DRAM/n1307 ,
         \unit_memory/DRAM/n1306 , \unit_memory/DRAM/n1305 ,
         \unit_memory/DRAM/n1304 , \unit_memory/DRAM/n1303 ,
         \unit_memory/DRAM/n1302 , \unit_memory/DRAM/n1301 ,
         \unit_memory/DRAM/n1300 , \unit_memory/DRAM/n1299 ,
         \unit_memory/DRAM/n1298 , \unit_memory/DRAM/n1297 ,
         \unit_memory/DRAM/n1296 , \unit_memory/DRAM/n1295 ,
         \unit_memory/DRAM/n1294 , \unit_memory/DRAM/n1293 ,
         \unit_memory/DRAM/n1292 , \unit_memory/DRAM/n1291 ,
         \unit_memory/DRAM/n1290 , \unit_memory/DRAM/n1289 ,
         \unit_memory/DRAM/n1288 , \unit_memory/DRAM/n1287 ,
         \unit_memory/DRAM/n1286 , \unit_memory/DRAM/n1285 ,
         \unit_memory/DRAM/n1284 , \unit_memory/DRAM/n1283 ,
         \unit_memory/DRAM/n1282 , \unit_memory/DRAM/n1281 ,
         \unit_memory/DRAM/n1280 , \unit_memory/DRAM/n1279 ,
         \unit_memory/DRAM/n1278 , \unit_memory/DRAM/n1277 ,
         \unit_memory/DRAM/n1276 , \unit_memory/DRAM/n1275 ,
         \unit_memory/DRAM/n1274 , \unit_memory/DRAM/n1273 ,
         \unit_memory/DRAM/n1272 , \unit_memory/DRAM/n1271 ,
         \unit_memory/DRAM/n1270 , \unit_memory/DRAM/n1269 ,
         \unit_memory/DRAM/n1268 , \unit_memory/DRAM/n1267 ,
         \unit_memory/DRAM/n1266 , \unit_memory/DRAM/n1265 ,
         \unit_memory/DRAM/n1264 , \unit_memory/DRAM/n1263 ,
         \unit_memory/DRAM/n1262 , \unit_memory/DRAM/n1261 ,
         \unit_memory/DRAM/n1260 , \unit_memory/DRAM/n1259 ,
         \unit_memory/DRAM/n1258 , \unit_memory/DRAM/n1257 ,
         \unit_memory/DRAM/n1256 , \unit_memory/DRAM/n1255 ,
         \unit_memory/DRAM/n1254 , \unit_memory/DRAM/n1253 ,
         \unit_memory/DRAM/n1252 , \unit_memory/DRAM/n1251 ,
         \unit_memory/DRAM/n1250 , \unit_memory/DRAM/n1249 ,
         \unit_memory/DRAM/n1248 , \unit_memory/DRAM/n1247 ,
         \unit_memory/DRAM/n1246 , \unit_memory/DRAM/n1245 ,
         \unit_memory/DRAM/n1244 , \unit_memory/DRAM/n1243 ,
         \unit_memory/DRAM/n1242 , \unit_memory/DRAM/n1241 ,
         \unit_memory/DRAM/n1240 , \unit_memory/DRAM/n1239 ,
         \unit_memory/DRAM/n1238 , \unit_memory/DRAM/n1237 ,
         \unit_memory/DRAM/n1236 , \unit_memory/DRAM/n1235 ,
         \unit_memory/DRAM/n1234 , \unit_memory/DRAM/n1233 ,
         \unit_memory/DRAM/n1232 , \unit_memory/DRAM/n1231 ,
         \unit_memory/DRAM/n1230 , \unit_memory/DRAM/n1229 ,
         \unit_memory/DRAM/n1228 , \unit_memory/DRAM/n1227 ,
         \unit_memory/DRAM/n1226 , \unit_memory/DRAM/n1225 ,
         \unit_memory/DRAM/n1224 , \unit_memory/DRAM/n1223 ,
         \unit_memory/DRAM/n1222 , \unit_memory/DRAM/n1221 ,
         \unit_memory/DRAM/n1220 , \unit_memory/DRAM/n1219 ,
         \unit_memory/DRAM/n1218 , \unit_memory/DRAM/n1217 ,
         \unit_memory/DRAM/n1216 , \unit_memory/DRAM/n1215 ,
         \unit_memory/DRAM/n1214 , \unit_memory/DRAM/n1213 ,
         \unit_memory/DRAM/n1212 , \unit_memory/DRAM/n1211 ,
         \unit_memory/DRAM/n1210 , \unit_memory/DRAM/n1209 ,
         \unit_memory/DRAM/n1208 , \unit_memory/DRAM/n1207 ,
         \unit_memory/DRAM/n1206 , \unit_memory/DRAM/n1205 ,
         \unit_memory/DRAM/n1204 , \unit_memory/DRAM/n1203 ,
         \unit_memory/DRAM/n1202 , \unit_memory/DRAM/n1201 ,
         \unit_memory/DRAM/n1200 , \unit_memory/DRAM/n1199 ,
         \unit_memory/DRAM/n1198 , \unit_memory/DRAM/n1197 ,
         \unit_memory/DRAM/n1196 , \unit_memory/DRAM/n1195 ,
         \unit_memory/DRAM/n1194 , \unit_memory/DRAM/n1193 ,
         \unit_memory/DRAM/n1192 , \unit_memory/DRAM/n1191 ,
         \unit_memory/DRAM/n1190 , \unit_memory/DRAM/n1189 ,
         \unit_memory/DRAM/n1188 , \unit_memory/DRAM/n1187 ,
         \unit_memory/DRAM/n1186 , \unit_memory/DRAM/n1185 ,
         \unit_memory/DRAM/n1184 , \unit_memory/DRAM/n1183 ,
         \unit_memory/DRAM/n1182 , \unit_memory/DRAM/n1181 ,
         \unit_memory/DRAM/n1180 , \unit_memory/DRAM/n1179 ,
         \unit_memory/DRAM/n1178 , \unit_memory/DRAM/n1177 ,
         \unit_memory/DRAM/n1176 , \unit_memory/DRAM/n1175 ,
         \unit_memory/DRAM/n1174 , \unit_memory/DRAM/n1173 ,
         \unit_memory/DRAM/n1172 , \unit_memory/DRAM/n1171 ,
         \unit_memory/DRAM/n1170 , \unit_memory/DRAM/n1169 ,
         \unit_memory/DRAM/n1168 , \unit_memory/DRAM/n1167 ,
         \unit_memory/DRAM/n1166 , \unit_memory/DRAM/n1165 ,
         \unit_memory/DRAM/n1164 , \unit_memory/DRAM/n1163 ,
         \unit_memory/DRAM/n1162 , \unit_memory/DRAM/n1161 ,
         \unit_memory/DRAM/n1160 , \unit_memory/DRAM/n1159 ,
         \unit_memory/DRAM/n1158 , \unit_memory/DRAM/n1157 ,
         \unit_memory/DRAM/N597 , \unit_memory/DRAM/N596 ,
         \unit_memory/DRAM/N595 , \unit_memory/DRAM/N594 ,
         \unit_memory/DRAM/N593 , \unit_memory/DRAM/N592 ,
         \unit_memory/DRAM/N591 , \unit_memory/DRAM/N590 ,
         \unit_memory/DRAM/N589 , \unit_memory/DRAM/N588 ,
         \unit_memory/DRAM/N587 , \unit_memory/DRAM/N586 ,
         \unit_memory/DRAM/N585 , \unit_memory/DRAM/N584 ,
         \unit_memory/DRAM/N583 , \unit_memory/DRAM/N582 ,
         \unit_memory/DRAM/N573 , \unit_memory/DRAM/N572 ,
         \unit_memory/DRAM/N571 , \unit_memory/DRAM/N570 ,
         \unit_memory/DRAM/N569 , \unit_memory/DRAM/N568 ,
         \unit_memory/DRAM/N567 , \unit_memory/DRAM/N566 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_0/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_0/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_31/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_31/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_30/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_30/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_29/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_29/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_28/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_28/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_27/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_27/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_26/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_26/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_25/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_25/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_24/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_24/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_23/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_23/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_22/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_22/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_21/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_21/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_20/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_20/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_19/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_19/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_18/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_18/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_17/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_17/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_16/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_16/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_15/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_15/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_14/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_14/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_13/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_13/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_12/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_12/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_11/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_11/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_10/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_10/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_9/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_9/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_8/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_8/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_7/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_7/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_6/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_6/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_5/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_5/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_4/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_4/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_3/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_3/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_2/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_2/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_1/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_1/Y1 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_0/Y2 ,
         \unit_memory/MUX21_NPCWB/MUX21GENI_0/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_31/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_31/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_30/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_30/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_29/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_29/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_28/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_28/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_27/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_27/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_26/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_26/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_25/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_25/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_24/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_24/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_23/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_23/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_22/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_22/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_21/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_21/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_20/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_20/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_19/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_19/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_18/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_18/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_17/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_17/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_16/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_16/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_15/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_15/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_14/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_14/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_13/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_13/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_12/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_12/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_11/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_11/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_10/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_10/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_9/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_9/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_8/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_8/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_7/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_7/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_6/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_6/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_5/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_5/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_4/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_4/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_3/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_3/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_2/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_2/Y1 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_1/Y2 ,
         \unit_memory/MUX21_ALMEM/MUX21GENI_1/Y1 , net126982, net126984,
         net127003, net130312, net130310, net130308, net130306, net130304,
         net130302, net130328, net130326, net130324, net130903, net130914,
         net130925, net141182, net141181, net141231, net141230, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
  wire   [4:0] rd1_out;
  wire   [4:0] cw_dec;
  wire   [10:0] cw_ex;
  wire   [8:0] cw_mem;
  wire   [31:0] alu_out;
  wire   [31:0] IR_OUT;
  wire   [4:0] wr_address;
  wire   [31:0] wr_data;
  wire   [31:0] npc1_out;
  wire   [31:0] rega_out;
  wire   [31:0] regb_out;
  wire   [31:0] imm_out;
  wire   [31:0] aluout_regn;
  wire   [31:0] bout_regn;
  wire   [31:0] npc2_out;

  EXUNIT_N32 unit_execution ( .NPC1(npc1_out), .RD1(rd1_out), .A(rega_out), 
        .B(regb_out), .IMM(imm_out), .S1_A_NPC(net141231), .S2_IMM_B(1'b0), 
        .ALU_OPCODE(cw_ex[5:0]), .CLK(CLK), .RST(n1322), .JUMP_EN({1'b0, 
        cw_ex[6]}), .EN_REGN_ALU_OUT(cw_ex[8]), .JUMP(jump), .ALUOUT(alu_out), 
        .ALU_OUT_REGN(aluout_regn), .B_OUT_REGN(bout_regn), .NPC2(npc2_out), 
        .RD2_OUT_REGN(wr_address) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_3/n6 ), .CK(CLK), .Q(cw_mem[3]), 
        .QN(n33) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_4/n5 ), .CK(CLK), .Q(cw_mem[4]) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_5/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_5/n5 ), .CK(CLK), .QN(n109) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_6/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_6/n6 ), .CK(CLK), .Q(cw_mem[6]), 
        .QN(n34) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_7/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_7/n5 ), .CK(CLK), .QN(n108) );
  DFF_X1 \unit_control/uut_third_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_3/n5 ), .CK(CLK), .QN(
        \unit_control/n383 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_4/n5 ), .CK(CLK), .QN(
        \unit_control/n400 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_5/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_5/n5 ), .CK(CLK), .QN(
        \unit_control/n399 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_6/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_6/n5 ), .CK(CLK), .QN(
        \unit_control/n382 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_7/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_7/n5 ), .CK(CLK), .QN(
        \unit_control/n398 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_13/n5 ), .CK(CLK), .Q(cw_ex[4]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_14/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_14/n5 ), .CK(CLK), .Q(cw_ex[5]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_15/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_15/n5 ), .CK(CLK), .Q(cw_ex[6]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_17/n6 ), .CK(CLK), .Q(cw_ex[8]) );
  DFF_X1 \unit_control/uut_second_stage/ffi_23/Q_reg  ( .D(n99), .CK(CLK), .Q(
        cw_dec[3]) );
  DFF_X1 \unit_control/uut_second_stage/ffi_22/Q_reg  ( .D(n1352), .CK(CLK), 
        .Q(cw_dec[2]), .QN(n2) );
  DFF_X1 \unit_control/uut_second_stage/ffi_21/Q_reg  ( .D(\unit_control/n418 ), .CK(CLK), .Q(cw_dec[1]), .QN(\unit_decode/n2189 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_17/n5 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_17/n2 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_14/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_14/n5 ), .CK(CLK), .QN(
        \unit_control/n386 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_13/n5 ), .CK(CLK), .QN(
        \unit_control/n387 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_12/n5 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_12/n2 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_11/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_11/n5 ), .CK(CLK), .QN(
        \unit_control/n378 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_10/n5 ), .CK(CLK), .QN(
        \unit_control/n379 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_9/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_9/n5 ), .CK(CLK), .QN(
        \unit_control/n381 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_7/Q_reg  ( .D(n99), .CK(CLK), .QN(
        \unit_control/n389 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_6/Q_reg  ( .D(n99), .CK(CLK), .QN(
        \unit_control/n390 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_5/Q_reg  ( .D(n99), .CK(CLK), .QN(
        \unit_control/n391 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_4/n5 ), .CK(CLK), .QN(
        \unit_control/n392 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_3/Q_reg  ( .D(n49), .CK(CLK), .QN(
        \unit_control/n393 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_19/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_19/n6 ), .CK(CLK), .QN(net141230) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_13/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_13/n5 ), .CK(CLK), .QN(n112) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[16]  ( .D(
        \unit_fetch/n447 ), .CK(CLK), .Q(IR_OUT[16]), .QN(\unit_decode/n2100 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[21]  ( .D(
        \unit_fetch/n462 ), .CK(CLK), .Q(IR_OUT[21]), .QN(\unit_decode/n2095 )
         );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_1/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_1/n5 ), .CK(CLK), .Q(n36), .QN(
        \unit_fetch/n329 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_2/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_2/n5 ), .CK(CLK), .QN(
        \unit_decode/n2146 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_3/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_3/n5 ), .CK(CLK), .QN(
        \unit_decode/n2145 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_5/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_5/n5 ), .CK(CLK), .QN(
        \unit_decode/n2143 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_7/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_7/n5 ), .CK(CLK), .QN(
        \unit_decode/n2141 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_27/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_27/n5 ), .CK(CLK), .QN(
        \unit_decode/n2121 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_29/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_29/n5 ), .CK(CLK), .QN(
        \unit_decode/n2119 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_9/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_9/n5 ), .CK(CLK), .QN(
        \unit_decode/n2139 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_11/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_11/n5 ), .CK(CLK), .QN(
        \unit_decode/n2137 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_13/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_13/n5 ), .CK(CLK), .QN(
        \unit_decode/n2135 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_15/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_15/n5 ), .CK(CLK), .QN(
        \unit_decode/n2133 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_17/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_17/n5 ), .CK(CLK), .QN(
        \unit_decode/n2131 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_19/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_19/n5 ), .CK(CLK), .QN(
        \unit_decode/n2129 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_21/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_21/n5 ), .CK(CLK), .QN(
        \unit_decode/n2127 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_23/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_23/n5 ), .CK(CLK), .QN(
        \unit_decode/n2125 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_25/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_25/n5 ), .CK(CLK), .QN(
        \unit_decode/n2123 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[0]  ( .D(
        \unit_fetch/unit_instructionRegister/n98 ), .CK(CLK), .QN(
        \unit_decode/n2116 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[1]  ( .D(
        \unit_fetch/unit_instructionRegister/n97 ), .CK(CLK), .QN(
        \unit_decode/n2115 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[3]  ( .D(
        \unit_fetch/unit_instructionRegister/n95 ), .CK(CLK), .QN(
        \unit_decode/n2113 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[5]  ( .D(
        \unit_fetch/unit_instructionRegister/n93 ), .CK(CLK), .QN(
        \unit_decode/n2111 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[17]  ( .D(
        \unit_fetch/unit_instructionRegister/n81 ), .CK(CLK), .Q(IR_OUT[17]), 
        .QN(\unit_decode/n2099 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[4]  ( .D(
        \unit_fetch/unit_instructionRegister/n92 ), .CK(CLK), .QN(
        \unit_decode/n2112 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[12]  ( .D(
        \unit_fetch/unit_instructionRegister/n84 ), .CK(CLK), .Q(IR_OUT[12]), 
        .QN(\unit_decode/n2104 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[14]  ( .D(
        \unit_fetch/unit_instructionRegister/n84 ), .CK(CLK), .Q(IR_OUT[14]), 
        .QN(\unit_decode/n2102 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[30]  ( .D(
        \unit_fetch/unit_instructionRegister/n69 ), .CK(CLK), .QN(n63) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[6]  ( .D(
        \unit_fetch/unit_instructionRegister/n92 ), .CK(CLK), .QN(
        \unit_decode/n2110 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[20]  ( .D(n100), .CK(
        CLK), .Q(IR_OUT[20]), .QN(\unit_decode/n2096 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_31/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_31/n5 ), .CK(CLK), .QN(
        \unit_decode/n2117 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_30/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_30/n5 ), .CK(CLK), .QN(
        \unit_decode/n2118 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_28/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_28/n5 ), .CK(CLK), .QN(
        \unit_decode/n2120 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_26/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_26/n5 ), .CK(CLK), .QN(
        \unit_decode/n2122 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_24/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_24/n5 ), .CK(CLK), .QN(
        \unit_decode/n2124 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_22/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_22/n5 ), .CK(CLK), .QN(
        \unit_decode/n2126 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_20/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_20/n5 ), .CK(CLK), .QN(
        \unit_decode/n2128 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_18/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_18/n5 ), .CK(CLK), .QN(
        \unit_decode/n2130 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_16/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_16/n5 ), .CK(CLK), .QN(
        \unit_decode/n2132 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_14/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_14/n5 ), .CK(CLK), .QN(
        \unit_decode/n2134 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_12/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_12/n5 ), .CK(CLK), .QN(
        \unit_decode/n2136 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_10/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_10/n5 ), .CK(CLK), .QN(
        \unit_decode/n2138 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_8/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_8/n5 ), .CK(CLK), .QN(
        \unit_decode/n2140 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_6/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_6/n5 ), .CK(CLK), .QN(
        \unit_decode/n2142 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[24]  ( .D(
        \unit_fetch/unit_instructionRegister/n75 ), .CK(CLK), .Q(IR_OUT[24]), 
        .QN(\unit_decode/n2092 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[23]  ( .D(
        \unit_fetch/unit_instructionRegister/n67 ), .CK(CLK), .Q(IR_OUT[23]), 
        .QN(\unit_decode/n2093 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[19]  ( .D(
        \unit_fetch/unit_instructionRegister/n79 ), .CK(CLK), .Q(IR_OUT[19]), 
        .QN(\unit_decode/n2097 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[18]  ( .D(
        \unit_fetch/unit_instructionRegister/n80 ), .CK(CLK), .Q(IR_OUT[18]), 
        .QN(\unit_decode/n2098 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[15]  ( .D(
        \unit_fetch/unit_instructionRegister/n83 ), .CK(CLK), .Q(IR_OUT[15]), 
        .QN(\unit_decode/n2101 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[13]  ( .D(
        \unit_fetch/unit_instructionRegister/n85 ), .CK(CLK), .Q(IR_OUT[13]), 
        .QN(\unit_decode/n2103 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[11]  ( .D(
        \unit_fetch/unit_instructionRegister/n87 ), .CK(CLK), .Q(IR_OUT[11]), 
        .QN(\unit_decode/n2105 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[10]  ( .D(
        \unit_fetch/unit_instructionRegister/n88 ), .CK(CLK), .QN(
        \unit_decode/n2106 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[9]  ( .D(
        \unit_fetch/unit_instructionRegister/n89 ), .CK(CLK), .QN(
        \unit_decode/n2107 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[8]  ( .D(
        \unit_fetch/unit_instructionRegister/n90 ), .CK(CLK), .QN(
        \unit_decode/n2108 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[7]  ( .D(
        \unit_fetch/unit_instructionRegister/n91 ), .CK(CLK), .QN(
        \unit_decode/n2109 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[2]  ( .D(
        \unit_fetch/unit_instructionRegister/n96 ), .CK(CLK), .QN(
        \unit_decode/n2114 ) );
  NAND3_X1 \unit_decode/U3638  ( .A1(wr_address[1]), .A2(wr_address[0]), .A3(
        wr_address[2]), .ZN(\unit_decode/n2243 ) );
  NAND3_X1 \unit_decode/U3637  ( .A1(wr_address[3]), .A2(\unit_decode/n2244 ), 
        .A3(wr_address[4]), .ZN(\unit_decode/n2264 ) );
  NAND3_X1 \unit_decode/U3636  ( .A1(wr_address[1]), .A2(\unit_decode/n2185 ), 
        .A3(wr_address[2]), .ZN(\unit_decode/n2241 ) );
  NAND3_X1 \unit_decode/U3635  ( .A1(wr_address[0]), .A2(\unit_decode/n2184 ), 
        .A3(wr_address[2]), .ZN(\unit_decode/n2239 ) );
  NAND3_X1 \unit_decode/U3634  ( .A1(\unit_decode/n2185 ), .A2(
        \unit_decode/n2184 ), .A3(wr_address[2]), .ZN(\unit_decode/n2237 ) );
  NAND3_X1 \unit_decode/U3633  ( .A1(wr_address[0]), .A2(\unit_decode/n2183 ), 
        .A3(wr_address[1]), .ZN(\unit_decode/n2235 ) );
  NAND3_X1 \unit_decode/U3632  ( .A1(\unit_decode/n2185 ), .A2(
        \unit_decode/n2183 ), .A3(wr_address[1]), .ZN(\unit_decode/n2233 ) );
  NAND3_X1 \unit_decode/U3631  ( .A1(\unit_decode/n2184 ), .A2(
        \unit_decode/n2183 ), .A3(wr_address[0]), .ZN(\unit_decode/n2231 ) );
  NAND3_X1 \unit_decode/U3630  ( .A1(\unit_decode/n2184 ), .A2(
        \unit_decode/n2183 ), .A3(\unit_decode/n2185 ), .ZN(
        \unit_decode/n2229 ) );
  NAND3_X1 \unit_decode/U3629  ( .A1(\unit_decode/n2244 ), .A2(
        \unit_decode/n2182 ), .A3(wr_address[4]), .ZN(\unit_decode/n2255 ) );
  NAND3_X1 \unit_decode/U3628  ( .A1(\unit_decode/n2244 ), .A2(
        \unit_decode/n2165 ), .A3(wr_address[3]), .ZN(\unit_decode/n2246 ) );
  NAND3_X1 \unit_decode/U3627  ( .A1(\unit_decode/n2182 ), .A2(
        \unit_decode/n2165 ), .A3(\unit_decode/n2244 ), .ZN(
        \unit_decode/n2228 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][23]  ( .D(
        \unit_decode/RegisterFile/n1675 ), .CK(CLK), .QN(\unit_decode/n2084 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][23]  ( .D(
        \unit_decode/RegisterFile/n1643 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n9 ), .QN(\unit_decode/n2060 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][0]  ( .D(
        \unit_decode/RegisterFile/n1588 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n64 ), .QN(\unit_decode/n2059 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][1]  ( .D(
        \unit_decode/RegisterFile/n1589 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n63 ), .QN(\unit_decode/n2058 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][2]  ( .D(
        \unit_decode/RegisterFile/n1590 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n62 ), .QN(\unit_decode/n2057 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][3]  ( .D(
        \unit_decode/RegisterFile/n1591 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n61 ), .QN(\unit_decode/n2056 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][4]  ( .D(
        \unit_decode/RegisterFile/n1592 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n60 ), .QN(\unit_decode/n2055 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][5]  ( .D(
        \unit_decode/RegisterFile/n1593 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n59 ), .QN(\unit_decode/n2054 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][6]  ( .D(
        \unit_decode/RegisterFile/n1594 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n58 ), .QN(\unit_decode/n2053 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][7]  ( .D(
        \unit_decode/RegisterFile/n1595 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n57 ), .QN(\unit_decode/n2052 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][8]  ( .D(
        \unit_decode/RegisterFile/n1596 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n56 ), .QN(\unit_decode/n2051 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][9]  ( .D(
        \unit_decode/RegisterFile/n1597 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n55 ), .QN(\unit_decode/n2050 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][10]  ( .D(
        \unit_decode/RegisterFile/n1598 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n54 ), .QN(\unit_decode/n2049 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][11]  ( .D(
        \unit_decode/RegisterFile/n1599 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n53 ), .QN(\unit_decode/n2048 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][12]  ( .D(
        \unit_decode/RegisterFile/n1600 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n52 ), .QN(\unit_decode/n2047 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][13]  ( .D(
        \unit_decode/RegisterFile/n1601 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n51 ), .QN(\unit_decode/n2046 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][14]  ( .D(
        \unit_decode/RegisterFile/n1602 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n50 ), .QN(\unit_decode/n2045 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][15]  ( .D(
        \unit_decode/RegisterFile/n1603 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n49 ), .QN(\unit_decode/n2044 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][16]  ( .D(
        \unit_decode/RegisterFile/n1604 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n48 ), .QN(\unit_decode/n2043 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][17]  ( .D(
        \unit_decode/RegisterFile/n1605 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n47 ), .QN(\unit_decode/n2042 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][18]  ( .D(
        \unit_decode/RegisterFile/n1606 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n46 ), .QN(\unit_decode/n2041 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][19]  ( .D(
        \unit_decode/RegisterFile/n1607 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n45 ), .QN(\unit_decode/n2040 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][20]  ( .D(
        \unit_decode/RegisterFile/n1608 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n44 ), .QN(\unit_decode/n2039 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][21]  ( .D(
        \unit_decode/RegisterFile/n1609 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n43 ), .QN(\unit_decode/n2038 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][22]  ( .D(
        \unit_decode/RegisterFile/n1610 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n42 ), .QN(\unit_decode/n2037 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][23]  ( .D(
        \unit_decode/RegisterFile/n1611 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n41 ), .QN(\unit_decode/n2036 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][0]  ( .D(
        \unit_decode/RegisterFile/n1556 ), .CK(CLK), .QN(\unit_decode/n2035 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][1]  ( .D(
        \unit_decode/RegisterFile/n1557 ), .CK(CLK), .QN(\unit_decode/n2034 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][2]  ( .D(
        \unit_decode/RegisterFile/n1558 ), .CK(CLK), .QN(\unit_decode/n2033 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][3]  ( .D(
        \unit_decode/RegisterFile/n1559 ), .CK(CLK), .QN(\unit_decode/n2032 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][4]  ( .D(
        \unit_decode/RegisterFile/n1560 ), .CK(CLK), .QN(\unit_decode/n2031 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][5]  ( .D(
        \unit_decode/RegisterFile/n1561 ), .CK(CLK), .QN(\unit_decode/n2030 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][6]  ( .D(
        \unit_decode/RegisterFile/n1562 ), .CK(CLK), .QN(\unit_decode/n2029 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][7]  ( .D(
        \unit_decode/RegisterFile/n1563 ), .CK(CLK), .QN(\unit_decode/n2028 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][8]  ( .D(
        \unit_decode/RegisterFile/n1564 ), .CK(CLK), .QN(\unit_decode/n2027 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][9]  ( .D(
        \unit_decode/RegisterFile/n1565 ), .CK(CLK), .QN(\unit_decode/n2026 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][10]  ( .D(
        \unit_decode/RegisterFile/n1566 ), .CK(CLK), .QN(\unit_decode/n2025 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][11]  ( .D(
        \unit_decode/RegisterFile/n1567 ), .CK(CLK), .QN(\unit_decode/n2024 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][12]  ( .D(
        \unit_decode/RegisterFile/n1568 ), .CK(CLK), .QN(\unit_decode/n2023 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][13]  ( .D(
        \unit_decode/RegisterFile/n1569 ), .CK(CLK), .QN(\unit_decode/n2022 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][14]  ( .D(
        \unit_decode/RegisterFile/n1570 ), .CK(CLK), .QN(\unit_decode/n2021 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][15]  ( .D(
        \unit_decode/RegisterFile/n1571 ), .CK(CLK), .QN(\unit_decode/n2020 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][16]  ( .D(
        \unit_decode/RegisterFile/n1572 ), .CK(CLK), .QN(\unit_decode/n2019 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][17]  ( .D(
        \unit_decode/RegisterFile/n1573 ), .CK(CLK), .QN(\unit_decode/n2018 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][18]  ( .D(
        \unit_decode/RegisterFile/n1574 ), .CK(CLK), .QN(\unit_decode/n2017 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][19]  ( .D(
        \unit_decode/RegisterFile/n1575 ), .CK(CLK), .QN(\unit_decode/n2016 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][20]  ( .D(
        \unit_decode/RegisterFile/n1576 ), .CK(CLK), .QN(\unit_decode/n2015 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][21]  ( .D(
        \unit_decode/RegisterFile/n1577 ), .CK(CLK), .QN(\unit_decode/n2014 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][22]  ( .D(
        \unit_decode/RegisterFile/n1578 ), .CK(CLK), .QN(\unit_decode/n2013 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][23]  ( .D(
        \unit_decode/RegisterFile/n1579 ), .CK(CLK), .QN(\unit_decode/n2012 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][0]  ( .D(
        \unit_decode/RegisterFile/n1140 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n512 ), .QN(\unit_decode/n1963 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][1]  ( .D(
        \unit_decode/RegisterFile/n1141 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n511 ), .QN(\unit_decode/n1962 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][2]  ( .D(
        \unit_decode/RegisterFile/n1142 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n510 ), .QN(\unit_decode/n1961 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][3]  ( .D(
        \unit_decode/RegisterFile/n1143 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n509 ), .QN(\unit_decode/n1960 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][4]  ( .D(
        \unit_decode/RegisterFile/n1144 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n508 ), .QN(\unit_decode/n1959 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][5]  ( .D(
        \unit_decode/RegisterFile/n1145 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n507 ), .QN(\unit_decode/n1958 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][6]  ( .D(
        \unit_decode/RegisterFile/n1146 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n506 ), .QN(\unit_decode/n1957 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][7]  ( .D(
        \unit_decode/RegisterFile/n1147 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n505 ), .QN(\unit_decode/n1956 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][24]  ( .D(
        \unit_decode/RegisterFile/n2156 ), .CK(CLK), .Q(\unit_decode/n4112 ), 
        .QN(\unit_decode/n1955 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][25]  ( .D(
        \unit_decode/RegisterFile/n2157 ), .CK(CLK), .Q(\unit_decode/n4108 ), 
        .QN(\unit_decode/n1954 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][26]  ( .D(
        \unit_decode/RegisterFile/n2158 ), .CK(CLK), .Q(\unit_decode/n4104 ), 
        .QN(\unit_decode/n1953 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][27]  ( .D(
        \unit_decode/RegisterFile/n2159 ), .CK(CLK), .Q(\unit_decode/n4100 ), 
        .QN(\unit_decode/n1952 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][28]  ( .D(
        \unit_decode/RegisterFile/n2160 ), .CK(CLK), .Q(\unit_decode/n4096 ), 
        .QN(\unit_decode/n1951 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][29]  ( .D(
        \unit_decode/RegisterFile/n2161 ), .CK(CLK), .Q(\unit_decode/n4092 ), 
        .QN(\unit_decode/n1950 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][30]  ( .D(
        \unit_decode/RegisterFile/n2162 ), .CK(CLK), .Q(\unit_decode/n4016 ), 
        .QN(\unit_decode/n1949 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][31]  ( .D(
        \unit_decode/RegisterFile/n2163 ), .CK(CLK), .Q(\unit_decode/n4012 ), 
        .QN(\unit_decode/n1948 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][24]  ( .D(
        \unit_decode/RegisterFile/n2124 ), .CK(CLK), .Q(\unit_decode/n3862 ), 
        .QN(\unit_decode/n1947 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][25]  ( .D(
        \unit_decode/RegisterFile/n2125 ), .CK(CLK), .Q(\unit_decode/n3856 ), 
        .QN(\unit_decode/n1946 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][26]  ( .D(
        \unit_decode/RegisterFile/n2126 ), .CK(CLK), .Q(\unit_decode/n3850 ), 
        .QN(\unit_decode/n1945 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][27]  ( .D(
        \unit_decode/RegisterFile/n2127 ), .CK(CLK), .Q(\unit_decode/n3844 ), 
        .QN(\unit_decode/n1944 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][28]  ( .D(
        \unit_decode/RegisterFile/n2128 ), .CK(CLK), .Q(\unit_decode/n3838 ), 
        .QN(\unit_decode/n1943 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][29]  ( .D(
        \unit_decode/RegisterFile/n2129 ), .CK(CLK), .Q(\unit_decode/n3832 ), 
        .QN(\unit_decode/n1942 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][30]  ( .D(
        \unit_decode/RegisterFile/n2130 ), .CK(CLK), .Q(\unit_decode/n3646 ), 
        .QN(\unit_decode/n1941 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][31]  ( .D(
        \unit_decode/RegisterFile/n2131 ), .CK(CLK), .Q(\unit_decode/n3640 ), 
        .QN(\unit_decode/n1940 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][24]  ( .D(
        \unit_decode/RegisterFile/n2092 ), .CK(CLK), .QN(\unit_decode/n1939 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][25]  ( .D(
        \unit_decode/RegisterFile/n2093 ), .CK(CLK), .QN(\unit_decode/n1938 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][26]  ( .D(
        \unit_decode/RegisterFile/n2094 ), .CK(CLK), .QN(\unit_decode/n1937 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][27]  ( .D(
        \unit_decode/RegisterFile/n2095 ), .CK(CLK), .QN(\unit_decode/n1936 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][28]  ( .D(
        \unit_decode/RegisterFile/n2096 ), .CK(CLK), .QN(\unit_decode/n1935 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][29]  ( .D(
        \unit_decode/RegisterFile/n2097 ), .CK(CLK), .QN(\unit_decode/n1934 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][30]  ( .D(
        \unit_decode/RegisterFile/n2098 ), .CK(CLK), .QN(\unit_decode/n1933 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][31]  ( .D(
        \unit_decode/RegisterFile/n2099 ), .CK(CLK), .QN(\unit_decode/n1932 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][24]  ( .D(
        \unit_decode/RegisterFile/n2060 ), .CK(CLK), .QN(\unit_decode/n1931 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][25]  ( .D(
        \unit_decode/RegisterFile/n2061 ), .CK(CLK), .QN(\unit_decode/n1930 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][26]  ( .D(
        \unit_decode/RegisterFile/n2062 ), .CK(CLK), .QN(\unit_decode/n1929 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][27]  ( .D(
        \unit_decode/RegisterFile/n2063 ), .CK(CLK), .QN(\unit_decode/n1928 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][28]  ( .D(
        \unit_decode/RegisterFile/n2064 ), .CK(CLK), .QN(\unit_decode/n1927 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][29]  ( .D(
        \unit_decode/RegisterFile/n2065 ), .CK(CLK), .QN(\unit_decode/n1926 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][30]  ( .D(
        \unit_decode/RegisterFile/n2066 ), .CK(CLK), .QN(\unit_decode/n1925 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][31]  ( .D(
        \unit_decode/RegisterFile/n2067 ), .CK(CLK), .QN(\unit_decode/n1924 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][24]  ( .D(
        \unit_decode/RegisterFile/n2028 ), .CK(CLK), .Q(\unit_decode/n4114 ), 
        .QN(\unit_decode/n1923 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][25]  ( .D(
        \unit_decode/RegisterFile/n2029 ), .CK(CLK), .Q(\unit_decode/n4110 ), 
        .QN(\unit_decode/n1922 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][26]  ( .D(
        \unit_decode/RegisterFile/n2030 ), .CK(CLK), .Q(\unit_decode/n4106 ), 
        .QN(\unit_decode/n1921 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][27]  ( .D(
        \unit_decode/RegisterFile/n2031 ), .CK(CLK), .Q(\unit_decode/n4102 ), 
        .QN(\unit_decode/n1920 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][28]  ( .D(
        \unit_decode/RegisterFile/n2032 ), .CK(CLK), .Q(\unit_decode/n4098 ), 
        .QN(\unit_decode/n1919 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][29]  ( .D(
        \unit_decode/RegisterFile/n2033 ), .CK(CLK), .Q(\unit_decode/n4094 ), 
        .QN(\unit_decode/n1918 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][30]  ( .D(
        \unit_decode/RegisterFile/n2034 ), .CK(CLK), .Q(\unit_decode/n4018 ), 
        .QN(\unit_decode/n1917 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][31]  ( .D(
        \unit_decode/RegisterFile/n2035 ), .CK(CLK), .Q(\unit_decode/n4014 ), 
        .QN(\unit_decode/n1916 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][24]  ( .D(
        \unit_decode/RegisterFile/n1996 ), .CK(CLK), .Q(\unit_decode/n3682 ), 
        .QN(\unit_decode/n1915 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][25]  ( .D(
        \unit_decode/RegisterFile/n1997 ), .CK(CLK), .Q(\unit_decode/n3676 ), 
        .QN(\unit_decode/n1914 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][26]  ( .D(
        \unit_decode/RegisterFile/n1998 ), .CK(CLK), .Q(\unit_decode/n3670 ), 
        .QN(\unit_decode/n1913 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][27]  ( .D(
        \unit_decode/RegisterFile/n1999 ), .CK(CLK), .Q(\unit_decode/n3664 ), 
        .QN(\unit_decode/n1912 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][28]  ( .D(
        \unit_decode/RegisterFile/n2000 ), .CK(CLK), .Q(\unit_decode/n3658 ), 
        .QN(\unit_decode/n1911 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][29]  ( .D(
        \unit_decode/RegisterFile/n2001 ), .CK(CLK), .Q(\unit_decode/n3652 ), 
        .QN(\unit_decode/n1910 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][30]  ( .D(
        \unit_decode/RegisterFile/n2002 ), .CK(CLK), .Q(\unit_decode/n3634 ), 
        .QN(\unit_decode/n1909 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][31]  ( .D(
        \unit_decode/RegisterFile/n2003 ), .CK(CLK), .Q(\unit_decode/n3628 ), 
        .QN(\unit_decode/n1908 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][24]  ( .D(
        \unit_decode/RegisterFile/n1964 ), .CK(CLK), .QN(\unit_decode/n1907 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][25]  ( .D(
        \unit_decode/RegisterFile/n1965 ), .CK(CLK), .QN(\unit_decode/n1906 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][26]  ( .D(
        \unit_decode/RegisterFile/n1966 ), .CK(CLK), .QN(\unit_decode/n1905 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][27]  ( .D(
        \unit_decode/RegisterFile/n1967 ), .CK(CLK), .QN(\unit_decode/n1904 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][28]  ( .D(
        \unit_decode/RegisterFile/n1968 ), .CK(CLK), .QN(\unit_decode/n1903 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][29]  ( .D(
        \unit_decode/RegisterFile/n1969 ), .CK(CLK), .QN(\unit_decode/n1902 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][30]  ( .D(
        \unit_decode/RegisterFile/n1970 ), .CK(CLK), .QN(\unit_decode/n1901 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][31]  ( .D(
        \unit_decode/RegisterFile/n1971 ), .CK(CLK), .QN(\unit_decode/n1900 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][24]  ( .D(
        \unit_decode/RegisterFile/n1932 ), .CK(CLK), .QN(\unit_decode/n1899 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][25]  ( .D(
        \unit_decode/RegisterFile/n1933 ), .CK(CLK), .QN(\unit_decode/n1898 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][26]  ( .D(
        \unit_decode/RegisterFile/n1934 ), .CK(CLK), .QN(\unit_decode/n1897 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][27]  ( .D(
        \unit_decode/RegisterFile/n1935 ), .CK(CLK), .QN(\unit_decode/n1896 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][28]  ( .D(
        \unit_decode/RegisterFile/n1936 ), .CK(CLK), .QN(\unit_decode/n1895 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][29]  ( .D(
        \unit_decode/RegisterFile/n1937 ), .CK(CLK), .QN(\unit_decode/n1894 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][30]  ( .D(
        \unit_decode/RegisterFile/n1938 ), .CK(CLK), .QN(\unit_decode/n1893 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][31]  ( .D(
        \unit_decode/RegisterFile/n1939 ), .CK(CLK), .QN(\unit_decode/n1892 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][24]  ( .D(
        \unit_decode/RegisterFile/n1260 ), .CK(CLK), .QN(\unit_decode/n1875 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][25]  ( .D(
        \unit_decode/RegisterFile/n1261 ), .CK(CLK), .QN(\unit_decode/n1874 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][26]  ( .D(
        \unit_decode/RegisterFile/n1262 ), .CK(CLK), .QN(\unit_decode/n1873 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][27]  ( .D(
        \unit_decode/RegisterFile/n1263 ), .CK(CLK), .QN(\unit_decode/n1872 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][28]  ( .D(
        \unit_decode/RegisterFile/n1264 ), .CK(CLK), .QN(\unit_decode/n1871 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][24]  ( .D(
        \unit_decode/RegisterFile/n1228 ), .CK(CLK), .QN(\unit_decode/n1870 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][25]  ( .D(
        \unit_decode/RegisterFile/n1229 ), .CK(CLK), .QN(\unit_decode/n1869 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][26]  ( .D(
        \unit_decode/RegisterFile/n1230 ), .CK(CLK), .QN(\unit_decode/n1868 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][27]  ( .D(
        \unit_decode/RegisterFile/n1231 ), .CK(CLK), .QN(\unit_decode/n1867 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][28]  ( .D(
        \unit_decode/RegisterFile/n1232 ), .CK(CLK), .QN(\unit_decode/n1866 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][29]  ( .D(
        \unit_decode/RegisterFile/n1233 ), .CK(CLK), .QN(\unit_decode/n1865 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][30]  ( .D(
        \unit_decode/RegisterFile/n1234 ), .CK(CLK), .QN(\unit_decode/n1864 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][31]  ( .D(
        \unit_decode/RegisterFile/n1235 ), .CK(CLK), .QN(\unit_decode/n1863 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][24]  ( .D(
        \unit_decode/RegisterFile/n1196 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n456 ), .QN(\unit_decode/n1862 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][25]  ( .D(
        \unit_decode/RegisterFile/n1197 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n455 ), .QN(\unit_decode/n1861 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][26]  ( .D(
        \unit_decode/RegisterFile/n1198 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n454 ), .QN(\unit_decode/n1860 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][27]  ( .D(
        \unit_decode/RegisterFile/n1199 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n453 ), .QN(\unit_decode/n1859 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][28]  ( .D(
        \unit_decode/RegisterFile/n1200 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n452 ), .QN(\unit_decode/n1858 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][29]  ( .D(
        \unit_decode/RegisterFile/n1201 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n451 ), .QN(\unit_decode/n1857 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][30]  ( .D(
        \unit_decode/RegisterFile/n1202 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n450 ), .QN(\unit_decode/n1856 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][31]  ( .D(
        \unit_decode/RegisterFile/n1203 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n449 ), .QN(\unit_decode/n1855 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][24]  ( .D(
        \unit_decode/RegisterFile/n1900 ), .CK(CLK), .Q(\unit_decode/n4111 ), 
        .QN(\unit_decode/n1854 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][25]  ( .D(
        \unit_decode/RegisterFile/n1901 ), .CK(CLK), .Q(\unit_decode/n4107 ), 
        .QN(\unit_decode/n1853 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][26]  ( .D(
        \unit_decode/RegisterFile/n1902 ), .CK(CLK), .Q(\unit_decode/n4103 ), 
        .QN(\unit_decode/n1852 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][27]  ( .D(
        \unit_decode/RegisterFile/n1903 ), .CK(CLK), .Q(\unit_decode/n4099 ), 
        .QN(\unit_decode/n1851 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][28]  ( .D(
        \unit_decode/RegisterFile/n1904 ), .CK(CLK), .Q(\unit_decode/n4095 ), 
        .QN(\unit_decode/n1850 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][29]  ( .D(
        \unit_decode/RegisterFile/n1905 ), .CK(CLK), .Q(\unit_decode/n4091 ), 
        .QN(\unit_decode/n1849 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][30]  ( .D(
        \unit_decode/RegisterFile/n1906 ), .CK(CLK), .Q(\unit_decode/n4015 ), 
        .QN(\unit_decode/n1848 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][31]  ( .D(
        \unit_decode/RegisterFile/n1907 ), .CK(CLK), .Q(\unit_decode/n4011 ), 
        .QN(\unit_decode/n1847 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][24]  ( .D(
        \unit_decode/RegisterFile/n1868 ), .CK(CLK), .Q(\unit_decode/n3861 ), 
        .QN(\unit_decode/n1846 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][25]  ( .D(
        \unit_decode/RegisterFile/n1869 ), .CK(CLK), .Q(\unit_decode/n3855 ), 
        .QN(\unit_decode/n1845 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][26]  ( .D(
        \unit_decode/RegisterFile/n1870 ), .CK(CLK), .Q(\unit_decode/n3849 ), 
        .QN(\unit_decode/n1844 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][27]  ( .D(
        \unit_decode/RegisterFile/n1871 ), .CK(CLK), .Q(\unit_decode/n3843 ), 
        .QN(\unit_decode/n1843 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][28]  ( .D(
        \unit_decode/RegisterFile/n1872 ), .CK(CLK), .Q(\unit_decode/n3837 ), 
        .QN(\unit_decode/n1842 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][29]  ( .D(
        \unit_decode/RegisterFile/n1873 ), .CK(CLK), .Q(\unit_decode/n3831 ), 
        .QN(\unit_decode/n1841 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][30]  ( .D(
        \unit_decode/RegisterFile/n1874 ), .CK(CLK), .Q(\unit_decode/n3645 ), 
        .QN(\unit_decode/n1840 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][31]  ( .D(
        \unit_decode/RegisterFile/n1875 ), .CK(CLK), .Q(\unit_decode/n3639 ), 
        .QN(\unit_decode/n1839 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][24]  ( .D(
        \unit_decode/RegisterFile/n1836 ), .CK(CLK), .QN(\unit_decode/n1838 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][25]  ( .D(
        \unit_decode/RegisterFile/n1837 ), .CK(CLK), .QN(\unit_decode/n1837 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][26]  ( .D(
        \unit_decode/RegisterFile/n1838 ), .CK(CLK), .QN(\unit_decode/n1836 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][27]  ( .D(
        \unit_decode/RegisterFile/n1839 ), .CK(CLK), .QN(\unit_decode/n1835 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][28]  ( .D(
        \unit_decode/RegisterFile/n1840 ), .CK(CLK), .QN(\unit_decode/n1834 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][29]  ( .D(
        \unit_decode/RegisterFile/n1841 ), .CK(CLK), .QN(\unit_decode/n1833 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][30]  ( .D(
        \unit_decode/RegisterFile/n1842 ), .CK(CLK), .QN(\unit_decode/n1832 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][31]  ( .D(
        \unit_decode/RegisterFile/n1843 ), .CK(CLK), .QN(\unit_decode/n1831 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][24]  ( .D(
        \unit_decode/RegisterFile/n1804 ), .CK(CLK), .QN(\unit_decode/n1830 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][25]  ( .D(
        \unit_decode/RegisterFile/n1805 ), .CK(CLK), .QN(\unit_decode/n1829 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][26]  ( .D(
        \unit_decode/RegisterFile/n1806 ), .CK(CLK), .QN(\unit_decode/n1828 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][27]  ( .D(
        \unit_decode/RegisterFile/n1807 ), .CK(CLK), .QN(\unit_decode/n1827 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][28]  ( .D(
        \unit_decode/RegisterFile/n1808 ), .CK(CLK), .QN(\unit_decode/n1826 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][29]  ( .D(
        \unit_decode/RegisterFile/n1809 ), .CK(CLK), .QN(\unit_decode/n1825 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][30]  ( .D(
        \unit_decode/RegisterFile/n1810 ), .CK(CLK), .QN(\unit_decode/n1824 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][31]  ( .D(
        \unit_decode/RegisterFile/n1811 ), .CK(CLK), .QN(\unit_decode/n1823 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][24]  ( .D(
        \unit_decode/RegisterFile/n1772 ), .CK(CLK), .Q(\unit_decode/n4113 ), 
        .QN(\unit_decode/n1822 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][25]  ( .D(
        \unit_decode/RegisterFile/n1773 ), .CK(CLK), .Q(\unit_decode/n4109 ), 
        .QN(\unit_decode/n1821 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][26]  ( .D(
        \unit_decode/RegisterFile/n1774 ), .CK(CLK), .Q(\unit_decode/n4105 ), 
        .QN(\unit_decode/n1820 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][27]  ( .D(
        \unit_decode/RegisterFile/n1775 ), .CK(CLK), .Q(\unit_decode/n4101 ), 
        .QN(\unit_decode/n1819 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][28]  ( .D(
        \unit_decode/RegisterFile/n1776 ), .CK(CLK), .Q(\unit_decode/n4097 ), 
        .QN(\unit_decode/n1818 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][29]  ( .D(
        \unit_decode/RegisterFile/n1777 ), .CK(CLK), .Q(\unit_decode/n4093 ), 
        .QN(\unit_decode/n1817 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][30]  ( .D(
        \unit_decode/RegisterFile/n1778 ), .CK(CLK), .Q(\unit_decode/n4017 ), 
        .QN(\unit_decode/n1816 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][31]  ( .D(
        \unit_decode/RegisterFile/n1779 ), .CK(CLK), .Q(\unit_decode/n4013 ), 
        .QN(\unit_decode/n1815 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][24]  ( .D(
        \unit_decode/RegisterFile/n1740 ), .CK(CLK), .Q(\unit_decode/n3681 ), 
        .QN(\unit_decode/n1814 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][25]  ( .D(
        \unit_decode/RegisterFile/n1741 ), .CK(CLK), .Q(\unit_decode/n3675 ), 
        .QN(\unit_decode/n1813 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][26]  ( .D(
        \unit_decode/RegisterFile/n1742 ), .CK(CLK), .Q(\unit_decode/n3669 ), 
        .QN(\unit_decode/n1812 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][27]  ( .D(
        \unit_decode/RegisterFile/n1743 ), .CK(CLK), .Q(\unit_decode/n3663 ), 
        .QN(\unit_decode/n1811 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][28]  ( .D(
        \unit_decode/RegisterFile/n1744 ), .CK(CLK), .Q(\unit_decode/n3657 ), 
        .QN(\unit_decode/n1810 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][29]  ( .D(
        \unit_decode/RegisterFile/n1745 ), .CK(CLK), .Q(\unit_decode/n3651 ), 
        .QN(\unit_decode/n1809 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][30]  ( .D(
        \unit_decode/RegisterFile/n1746 ), .CK(CLK), .Q(\unit_decode/n3633 ), 
        .QN(\unit_decode/n1808 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][31]  ( .D(
        \unit_decode/RegisterFile/n1747 ), .CK(CLK), .Q(\unit_decode/n3627 ), 
        .QN(\unit_decode/n1807 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][24]  ( .D(
        \unit_decode/RegisterFile/n1708 ), .CK(CLK), .QN(\unit_decode/n1806 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][25]  ( .D(
        \unit_decode/RegisterFile/n1709 ), .CK(CLK), .QN(\unit_decode/n1805 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][26]  ( .D(
        \unit_decode/RegisterFile/n1710 ), .CK(CLK), .QN(\unit_decode/n1804 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][27]  ( .D(
        \unit_decode/RegisterFile/n1711 ), .CK(CLK), .QN(\unit_decode/n1803 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][28]  ( .D(
        \unit_decode/RegisterFile/n1712 ), .CK(CLK), .QN(\unit_decode/n1802 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][29]  ( .D(
        \unit_decode/RegisterFile/n1713 ), .CK(CLK), .QN(\unit_decode/n1801 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][30]  ( .D(
        \unit_decode/RegisterFile/n1714 ), .CK(CLK), .QN(\unit_decode/n1800 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][31]  ( .D(
        \unit_decode/RegisterFile/n1715 ), .CK(CLK), .QN(\unit_decode/n1799 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][24]  ( .D(
        \unit_decode/RegisterFile/n1676 ), .CK(CLK), .QN(\unit_decode/n1798 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][25]  ( .D(
        \unit_decode/RegisterFile/n1677 ), .CK(CLK), .QN(\unit_decode/n1797 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][26]  ( .D(
        \unit_decode/RegisterFile/n1678 ), .CK(CLK), .QN(\unit_decode/n1796 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][27]  ( .D(
        \unit_decode/RegisterFile/n1679 ), .CK(CLK), .QN(\unit_decode/n1795 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][28]  ( .D(
        \unit_decode/RegisterFile/n1680 ), .CK(CLK), .QN(\unit_decode/n1794 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][29]  ( .D(
        \unit_decode/RegisterFile/n1681 ), .CK(CLK), .QN(\unit_decode/n1793 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][30]  ( .D(
        \unit_decode/RegisterFile/n1682 ), .CK(CLK), .QN(\unit_decode/n1792 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][31]  ( .D(
        \unit_decode/RegisterFile/n1683 ), .CK(CLK), .QN(\unit_decode/n1791 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][24]  ( .D(
        \unit_decode/RegisterFile/n1644 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n8 ), .QN(\unit_decode/n1790 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][25]  ( .D(
        \unit_decode/RegisterFile/n1645 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n7 ), .QN(\unit_decode/n1789 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][26]  ( .D(
        \unit_decode/RegisterFile/n1646 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n6 ), .QN(\unit_decode/n1788 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][27]  ( .D(
        \unit_decode/RegisterFile/n1647 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n5 ), .QN(\unit_decode/n1787 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][28]  ( .D(
        \unit_decode/RegisterFile/n1648 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n4 ), .QN(\unit_decode/n1786 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][24]  ( .D(
        \unit_decode/RegisterFile/n1612 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n40 ), .QN(\unit_decode/n1782 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][25]  ( .D(
        \unit_decode/RegisterFile/n1613 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n39 ), .QN(\unit_decode/n1781 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][26]  ( .D(
        \unit_decode/RegisterFile/n1614 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n38 ), .QN(\unit_decode/n1780 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][27]  ( .D(
        \unit_decode/RegisterFile/n1615 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n37 ), .QN(\unit_decode/n1779 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][28]  ( .D(
        \unit_decode/RegisterFile/n1616 ), .CK(CLK), .Q(
        \unit_decode/RegisterFile/n36 ), .QN(\unit_decode/n1778 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][24]  ( .D(
        \unit_decode/RegisterFile/n1580 ), .CK(CLK), .QN(\unit_decode/n1774 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][25]  ( .D(
        \unit_decode/RegisterFile/n1581 ), .CK(CLK), .QN(\unit_decode/n1773 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][26]  ( .D(
        \unit_decode/RegisterFile/n1582 ), .CK(CLK), .QN(\unit_decode/n1772 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][27]  ( .D(
        \unit_decode/RegisterFile/n1583 ), .CK(CLK), .QN(\unit_decode/n1771 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][28]  ( .D(
        \unit_decode/RegisterFile/n1584 ), .CK(CLK), .QN(\unit_decode/n1770 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][29]  ( .D(
        \unit_decode/RegisterFile/n1585 ), .CK(CLK), .QN(\unit_decode/n1769 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][30]  ( .D(
        \unit_decode/RegisterFile/n1586 ), .CK(CLK), .QN(\unit_decode/n1768 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[18][31]  ( .D(
        \unit_decode/RegisterFile/n1587 ), .CK(CLK), .QN(\unit_decode/n1767 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][29]  ( .D(
        \unit_decode/RegisterFile/n1553 ), .CK(CLK), .QN(\unit_decode/n1766 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][30]  ( .D(
        \unit_decode/RegisterFile/n1554 ), .CK(CLK), .QN(\unit_decode/n1765 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][31]  ( .D(
        \unit_decode/RegisterFile/n1555 ), .CK(CLK), .QN(\unit_decode/n1764 )
         );
  DFF_X1 \unit_decode/NPC1reg/ffi_17/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_17/n5 ), .CK(CLK), .Q(npc1_out[17]), .QN(
        \unit_decode/n3573 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_16/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_16/n5 ), .CK(CLK), .Q(npc1_out[16]), .QN(
        \unit_decode/n3574 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_15/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_15/n5 ), .CK(CLK), .Q(npc1_out[15]), .QN(
        \unit_decode/n3575 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_14/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_14/n5 ), .CK(CLK), .Q(npc1_out[14]), .QN(
        \unit_decode/n3576 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_13/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_13/n5 ), .CK(CLK), .Q(npc1_out[13]), .QN(
        \unit_decode/n3577 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_12/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_12/n5 ), .CK(CLK), .Q(npc1_out[12]), .QN(
        \unit_decode/n3578 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_11/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_11/n5 ), .CK(CLK), .Q(npc1_out[11]), .QN(
        \unit_decode/n3579 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_10/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_10/n5 ), .CK(CLK), .Q(npc1_out[10]), .QN(
        \unit_decode/n3580 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_9/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_9/n5 ), .CK(CLK), .Q(npc1_out[9]), .QN(\unit_decode/n3581 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_8/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_8/n5 ), .CK(CLK), .Q(npc1_out[8]), .QN(\unit_decode/n3582 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_7/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_7/n5 ), .CK(CLK), .Q(npc1_out[7]), .QN(\unit_decode/n3583 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_6/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_6/n5 ), .CK(CLK), .Q(npc1_out[6]), .QN(\unit_decode/n3584 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_5/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_5/n5 ), .CK(CLK), .Q(npc1_out[5]), .QN(\unit_decode/n3585 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_4/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_4/n5 ), .CK(CLK), .Q(npc1_out[4]), .QN(\unit_decode/n3586 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_3/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_3/n5 ), .CK(CLK), .Q(npc1_out[3]), .QN(\unit_decode/n217 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_1/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_1/n5 ), .CK(CLK), .Q(npc1_out[1]), .QN(\unit_decode/n205 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_0/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_0/n5 ), .CK(CLK), .Q(npc1_out[0]), .QN(\unit_decode/n201 ) );
  DFF_X1 \unit_decode/Areg/ffi_13/Q_reg  ( .D(\unit_decode/Areg/ffi_13/n5 ), 
        .CK(CLK), .Q(rega_out[13]), .QN(\unit_decode/n3528 ) );
  DFF_X1 \unit_decode/Areg/ffi_12/Q_reg  ( .D(\unit_decode/Areg/ffi_12/n5 ), 
        .CK(CLK), .Q(rega_out[12]), .QN(\unit_decode/n3529 ) );
  DFF_X1 \unit_decode/Areg/ffi_9/Q_reg  ( .D(\unit_decode/Areg/ffi_9/n5 ), 
        .CK(CLK), .Q(rega_out[9]), .QN(\unit_decode/n3532 ) );
  DFF_X1 \unit_decode/Areg/ffi_8/Q_reg  ( .D(\unit_decode/Areg/ffi_8/n5 ), 
        .CK(CLK), .Q(rega_out[8]), .QN(\unit_decode/n3533 ) );
  DFF_X1 \unit_decode/Areg/ffi_7/Q_reg  ( .D(\unit_decode/Areg/ffi_7/n5 ), 
        .CK(CLK), .Q(rega_out[7]), .QN(\unit_decode/n3534 ) );
  DFF_X1 \unit_decode/Areg/ffi_5/Q_reg  ( .D(\unit_decode/Areg/ffi_5/n5 ), 
        .CK(CLK), .Q(rega_out[5]), .QN(\unit_decode/n3536 ) );
  DFF_X1 \unit_decode/Areg/ffi_4/Q_reg  ( .D(\unit_decode/Areg/ffi_4/n5 ), 
        .CK(CLK), .Q(rega_out[4]), .QN(\unit_decode/n3537 ) );
  DFF_X1 \unit_decode/Areg/ffi_3/Q_reg  ( .D(\unit_decode/Areg/ffi_3/n5 ), 
        .CK(CLK), .Q(rega_out[3]), .QN(\unit_decode/n215 ) );
  DFF_X1 \unit_decode/Areg/ffi_1/Q_reg  ( .D(\unit_decode/Areg/ffi_1/n5 ), 
        .CK(CLK), .Q(rega_out[1]), .QN(\unit_decode/n203 ) );
  DFF_X1 \unit_decode/Areg/ffi_0/Q_reg  ( .D(\unit_decode/Areg/ffi_0/n5 ), 
        .CK(CLK), .Q(rega_out[0]), .QN(\unit_decode/n199 ) );
  DFF_X1 \unit_decode/Breg/ffi_30/Q_reg  ( .D(\unit_decode/Breg/ffi_30/n5 ), 
        .CK(CLK), .Q(regb_out[30]), .QN(\unit_decode/n3539 ) );
  DFF_X1 \unit_decode/Breg/ffi_29/Q_reg  ( .D(\unit_decode/Breg/ffi_29/n5 ), 
        .CK(CLK), .Q(regb_out[29]), .QN(\unit_decode/n3540 ) );
  DFF_X1 \unit_decode/Breg/ffi_28/Q_reg  ( .D(\unit_decode/Breg/ffi_28/n5 ), 
        .CK(CLK), .Q(regb_out[28]), .QN(\unit_decode/n3541 ) );
  DFF_X1 \unit_decode/Breg/ffi_27/Q_reg  ( .D(\unit_decode/Breg/ffi_27/n5 ), 
        .CK(CLK), .Q(regb_out[27]), .QN(\unit_decode/n3542 ) );
  DFF_X1 \unit_decode/Breg/ffi_26/Q_reg  ( .D(\unit_decode/Breg/ffi_26/n5 ), 
        .CK(CLK), .Q(regb_out[26]), .QN(\unit_decode/n3543 ) );
  DFF_X1 \unit_decode/Breg/ffi_25/Q_reg  ( .D(\unit_decode/Breg/ffi_25/n5 ), 
        .CK(CLK), .Q(regb_out[25]), .QN(\unit_decode/n3544 ) );
  DFF_X1 \unit_decode/Breg/ffi_24/Q_reg  ( .D(\unit_decode/Breg/ffi_24/n5 ), 
        .CK(CLK), .Q(regb_out[24]), .QN(\unit_decode/n3545 ) );
  DFF_X1 \unit_decode/Breg/ffi_23/Q_reg  ( .D(\unit_decode/Breg/ffi_23/n5 ), 
        .CK(CLK), .Q(regb_out[23]), .QN(\unit_decode/n3546 ) );
  DFF_X1 \unit_decode/Breg/ffi_22/Q_reg  ( .D(\unit_decode/Breg/ffi_22/n5 ), 
        .CK(CLK), .Q(regb_out[22]), .QN(\unit_decode/n3547 ) );
  DFF_X1 \unit_decode/Breg/ffi_21/Q_reg  ( .D(\unit_decode/Breg/ffi_21/n5 ), 
        .CK(CLK), .Q(regb_out[21]), .QN(\unit_decode/n3548 ) );
  DFF_X1 \unit_decode/Breg/ffi_20/Q_reg  ( .D(\unit_decode/Breg/ffi_20/n5 ), 
        .CK(CLK), .Q(regb_out[20]), .QN(\unit_decode/n3549 ) );
  DFF_X1 \unit_decode/Breg/ffi_3/Q_reg  ( .D(\unit_decode/Breg/ffi_3/n5 ), 
        .CK(CLK), .Q(regb_out[3]), .QN(\unit_decode/n235 ) );
  DFF_X1 \unit_decode/Breg/ffi_2/Q_reg  ( .D(\unit_decode/Breg/ffi_2/n5 ), 
        .CK(CLK), .Q(regb_out[2]), .QN(\unit_decode/n227 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_31/Q_reg  ( .D(\unit_decode/IMMreg/ffi_31/n5 ), .CK(CLK), .Q(imm_out[31]), .QN(\unit_decode/n3625 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_30/Q_reg  ( .D(\unit_decode/IMMreg/ffi_30/n5 ), .CK(CLK), .Q(imm_out[30]), .QN(\unit_decode/n3600 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_29/Q_reg  ( .D(\unit_decode/IMMreg/ffi_29/n5 ), .CK(CLK), .Q(imm_out[29]), .QN(\unit_decode/n3601 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_28/Q_reg  ( .D(\unit_decode/IMMreg/ffi_28/n5 ), .CK(CLK), .Q(imm_out[28]), .QN(\unit_decode/n3559 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_27/Q_reg  ( .D(\unit_decode/IMMreg/ffi_27/n5 ), .CK(CLK), .Q(imm_out[27]), .QN(\unit_decode/n3602 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_26/Q_reg  ( .D(\unit_decode/IMMreg/ffi_26/n5 ), .CK(CLK), .Q(imm_out[26]), .QN(\unit_decode/n3603 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_25/Q_reg  ( .D(\unit_decode/IMMreg/ffi_25/n5 ), .CK(CLK), .Q(imm_out[25]), .QN(\unit_decode/n3604 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_24/Q_reg  ( .D(\unit_decode/IMMreg/ffi_24/n5 ), .CK(CLK), .Q(imm_out[24]), .QN(\unit_decode/n3605 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_23/Q_reg  ( .D(\unit_decode/IMMreg/ffi_23/n5 ), .CK(CLK), .Q(imm_out[23]), .QN(\unit_decode/n3606 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_22/Q_reg  ( .D(\unit_decode/IMMreg/ffi_22/n5 ), .CK(CLK), .Q(imm_out[22]), .QN(\unit_decode/n3607 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_21/Q_reg  ( .D(\unit_decode/IMMreg/ffi_21/n5 ), .CK(CLK), .Q(imm_out[21]), .QN(\unit_decode/n3608 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_20/Q_reg  ( .D(\unit_decode/IMMreg/ffi_20/n5 ), .CK(CLK), .Q(imm_out[20]), .QN(\unit_decode/n3609 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_19/Q_reg  ( .D(\unit_decode/IMMreg/ffi_19/n5 ), .CK(CLK), .Q(imm_out[19]), .QN(\unit_decode/n3610 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_18/Q_reg  ( .D(\unit_decode/IMMreg/ffi_18/n5 ), .CK(CLK), .Q(imm_out[18]), .QN(\unit_decode/n3611 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_17/Q_reg  ( .D(\unit_decode/IMMreg/ffi_17/n5 ), .CK(CLK), .Q(imm_out[17]), .QN(\unit_decode/n3612 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_16/Q_reg  ( .D(\unit_decode/IMMreg/ffi_16/n5 ), .CK(CLK), .Q(imm_out[16]), .QN(\unit_decode/n3613 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_13/Q_reg  ( .D(\unit_decode/IMMreg/ffi_13/n5 ), .CK(CLK), .Q(imm_out[13]), .QN(\unit_decode/n3616 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_12/Q_reg  ( .D(\unit_decode/IMMreg/ffi_12/n5 ), .CK(CLK), .Q(imm_out[12]), .QN(\unit_decode/n3617 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_10/Q_reg  ( .D(\unit_decode/IMMreg/ffi_10/n5 ), .CK(CLK), .Q(imm_out[10]), .QN(\unit_decode/n3619 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_9/Q_reg  ( .D(\unit_decode/IMMreg/ffi_9/n5 ), 
        .CK(CLK), .Q(imm_out[9]), .QN(\unit_decode/n3620 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_8/Q_reg  ( .D(\unit_decode/IMMreg/ffi_8/n5 ), 
        .CK(CLK), .Q(imm_out[8]), .QN(\unit_decode/n3621 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_5/Q_reg  ( .D(\unit_decode/IMMreg/ffi_5/n5 ), 
        .CK(CLK), .Q(imm_out[5]), .QN(\unit_decode/n213 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_4/Q_reg  ( .D(\unit_decode/IMMreg/ffi_4/n5 ), 
        .CK(CLK), .Q(imm_out[4]), .QN(\unit_decode/n211 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_3/Q_reg  ( .D(\unit_decode/IMMreg/ffi_3/n5 ), 
        .CK(CLK), .Q(imm_out[3]), .QN(\unit_decode/n231 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_1/Q_reg  ( .D(\unit_decode/IMMreg/ffi_1/n5 ), 
        .CK(CLK), .Q(imm_out[1]), .QN(\unit_decode/n229 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][23]  ( .D(
        \unit_decode/RegisterFile/n2155 ), .CK(CLK), .Q(\unit_decode/n4116 ), 
        .QN(\unit_decode/n1747 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][22]  ( .D(
        \unit_decode/RegisterFile/n2154 ), .CK(CLK), .Q(\unit_decode/n4120 ), 
        .QN(\unit_decode/n1746 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][21]  ( .D(
        \unit_decode/RegisterFile/n2153 ), .CK(CLK), .Q(\unit_decode/n4124 ), 
        .QN(\unit_decode/n1745 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][20]  ( .D(
        \unit_decode/RegisterFile/n2152 ), .CK(CLK), .Q(\unit_decode/n4128 ), 
        .QN(\unit_decode/n1744 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][19]  ( .D(
        \unit_decode/RegisterFile/n2151 ), .CK(CLK), .Q(\unit_decode/n4132 ), 
        .QN(\unit_decode/n1743 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][18]  ( .D(
        \unit_decode/RegisterFile/n2150 ), .CK(CLK), .Q(\unit_decode/n4136 ), 
        .QN(\unit_decode/n1742 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][17]  ( .D(
        \unit_decode/RegisterFile/n2149 ), .CK(CLK), .Q(\unit_decode/n4020 ), 
        .QN(\unit_decode/n1741 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][16]  ( .D(
        \unit_decode/RegisterFile/n2148 ), .CK(CLK), .Q(\unit_decode/n4024 ), 
        .QN(\unit_decode/n1740 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][15]  ( .D(
        \unit_decode/RegisterFile/n2147 ), .CK(CLK), .Q(\unit_decode/n4028 ), 
        .QN(\unit_decode/n1739 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][14]  ( .D(
        \unit_decode/RegisterFile/n2146 ), .CK(CLK), .Q(\unit_decode/n4032 ), 
        .QN(\unit_decode/n1738 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][13]  ( .D(
        \unit_decode/RegisterFile/n2145 ), .CK(CLK), .Q(\unit_decode/n4036 ), 
        .QN(\unit_decode/n1737 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][12]  ( .D(
        \unit_decode/RegisterFile/n2144 ), .CK(CLK), .Q(\unit_decode/n4040 ), 
        .QN(\unit_decode/n1736 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][11]  ( .D(
        \unit_decode/RegisterFile/n2143 ), .CK(CLK), .Q(\unit_decode/n4044 ), 
        .QN(\unit_decode/n1735 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][10]  ( .D(
        \unit_decode/RegisterFile/n2142 ), .CK(CLK), .Q(\unit_decode/n4048 ), 
        .QN(\unit_decode/n1734 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][9]  ( .D(
        \unit_decode/RegisterFile/n2141 ), .CK(CLK), .Q(\unit_decode/n4052 ), 
        .QN(\unit_decode/n1733 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][8]  ( .D(
        \unit_decode/RegisterFile/n2140 ), .CK(CLK), .Q(\unit_decode/n4056 ), 
        .QN(\unit_decode/n1732 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][7]  ( .D(
        \unit_decode/RegisterFile/n2139 ), .CK(CLK), .Q(\unit_decode/n4060 ), 
        .QN(\unit_decode/n1731 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][6]  ( .D(
        \unit_decode/RegisterFile/n2138 ), .CK(CLK), .Q(\unit_decode/n4064 ), 
        .QN(\unit_decode/n1730 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][5]  ( .D(
        \unit_decode/RegisterFile/n2137 ), .CK(CLK), .Q(\unit_decode/n4068 ), 
        .QN(\unit_decode/n1729 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][4]  ( .D(
        \unit_decode/RegisterFile/n2136 ), .CK(CLK), .Q(\unit_decode/n4072 ), 
        .QN(\unit_decode/n1728 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][3]  ( .D(
        \unit_decode/RegisterFile/n2135 ), .CK(CLK), .Q(\unit_decode/n4076 ), 
        .QN(\unit_decode/n1727 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][2]  ( .D(
        \unit_decode/RegisterFile/n2134 ), .CK(CLK), .Q(\unit_decode/n4080 ), 
        .QN(\unit_decode/n1726 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][1]  ( .D(
        \unit_decode/RegisterFile/n2133 ), .CK(CLK), .Q(\unit_decode/n4084 ), 
        .QN(\unit_decode/n1725 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[0][0]  ( .D(
        \unit_decode/RegisterFile/n2132 ), .CK(CLK), .Q(\unit_decode/n4088 ), 
        .QN(\unit_decode/n1724 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][23]  ( .D(
        \unit_decode/RegisterFile/n2123 ), .CK(CLK), .Q(\unit_decode/n3868 ), 
        .QN(\unit_decode/n1723 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][22]  ( .D(
        \unit_decode/RegisterFile/n2122 ), .CK(CLK), .Q(\unit_decode/n3874 ), 
        .QN(\unit_decode/n1722 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][21]  ( .D(
        \unit_decode/RegisterFile/n2121 ), .CK(CLK), .Q(\unit_decode/n3880 ), 
        .QN(\unit_decode/n1721 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][20]  ( .D(
        \unit_decode/RegisterFile/n2120 ), .CK(CLK), .Q(\unit_decode/n3886 ), 
        .QN(\unit_decode/n1720 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][19]  ( .D(
        \unit_decode/RegisterFile/n2119 ), .CK(CLK), .Q(\unit_decode/n3892 ), 
        .QN(\unit_decode/n1719 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][18]  ( .D(
        \unit_decode/RegisterFile/n2118 ), .CK(CLK), .Q(\unit_decode/n3898 ), 
        .QN(\unit_decode/n1718 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][17]  ( .D(
        \unit_decode/RegisterFile/n2117 ), .CK(CLK), .Q(\unit_decode/n3904 ), 
        .QN(\unit_decode/n1717 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][16]  ( .D(
        \unit_decode/RegisterFile/n2116 ), .CK(CLK), .Q(\unit_decode/n3910 ), 
        .QN(\unit_decode/n1716 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][15]  ( .D(
        \unit_decode/RegisterFile/n2115 ), .CK(CLK), .Q(\unit_decode/n3916 ), 
        .QN(\unit_decode/n1715 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][14]  ( .D(
        \unit_decode/RegisterFile/n2114 ), .CK(CLK), .Q(\unit_decode/n3922 ), 
        .QN(\unit_decode/n1714 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][13]  ( .D(
        \unit_decode/RegisterFile/n2113 ), .CK(CLK), .Q(\unit_decode/n3928 ), 
        .QN(\unit_decode/n1713 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][12]  ( .D(
        \unit_decode/RegisterFile/n2112 ), .CK(CLK), .Q(\unit_decode/n3934 ), 
        .QN(\unit_decode/n1712 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][11]  ( .D(
        \unit_decode/RegisterFile/n2111 ), .CK(CLK), .Q(\unit_decode/n3940 ), 
        .QN(\unit_decode/n1711 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][10]  ( .D(
        \unit_decode/RegisterFile/n2110 ), .CK(CLK), .Q(\unit_decode/n3946 ), 
        .QN(\unit_decode/n1710 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][9]  ( .D(
        \unit_decode/RegisterFile/n2109 ), .CK(CLK), .Q(\unit_decode/n3952 ), 
        .QN(\unit_decode/n1709 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][8]  ( .D(
        \unit_decode/RegisterFile/n2108 ), .CK(CLK), .Q(\unit_decode/n3958 ), 
        .QN(\unit_decode/n1708 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][7]  ( .D(
        \unit_decode/RegisterFile/n2107 ), .CK(CLK), .Q(\unit_decode/n3964 ), 
        .QN(\unit_decode/n1707 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][6]  ( .D(
        \unit_decode/RegisterFile/n2106 ), .CK(CLK), .Q(\unit_decode/n3970 ), 
        .QN(\unit_decode/n1706 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][5]  ( .D(
        \unit_decode/RegisterFile/n2105 ), .CK(CLK), .Q(\unit_decode/n3976 ), 
        .QN(\unit_decode/n1705 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][4]  ( .D(
        \unit_decode/RegisterFile/n2104 ), .CK(CLK), .Q(\unit_decode/n3982 ), 
        .QN(\unit_decode/n1704 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][3]  ( .D(
        \unit_decode/RegisterFile/n2103 ), .CK(CLK), .Q(\unit_decode/n3988 ), 
        .QN(\unit_decode/n1703 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][2]  ( .D(
        \unit_decode/RegisterFile/n2102 ), .CK(CLK), .Q(\unit_decode/n3994 ), 
        .QN(\unit_decode/n1702 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][1]  ( .D(
        \unit_decode/RegisterFile/n2101 ), .CK(CLK), .Q(\unit_decode/n4000 ), 
        .QN(\unit_decode/n1701 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[1][0]  ( .D(
        \unit_decode/RegisterFile/n2100 ), .CK(CLK), .Q(\unit_decode/n4006 ), 
        .QN(\unit_decode/n1700 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][23]  ( .D(
        \unit_decode/RegisterFile/n2091 ), .CK(CLK), .QN(\unit_decode/n1699 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][22]  ( .D(
        \unit_decode/RegisterFile/n2090 ), .CK(CLK), .QN(\unit_decode/n1698 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][21]  ( .D(
        \unit_decode/RegisterFile/n2089 ), .CK(CLK), .QN(\unit_decode/n1697 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][20]  ( .D(
        \unit_decode/RegisterFile/n2088 ), .CK(CLK), .QN(\unit_decode/n1696 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][19]  ( .D(
        \unit_decode/RegisterFile/n2087 ), .CK(CLK), .QN(\unit_decode/n1695 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][18]  ( .D(
        \unit_decode/RegisterFile/n2086 ), .CK(CLK), .QN(\unit_decode/n1694 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][17]  ( .D(
        \unit_decode/RegisterFile/n2085 ), .CK(CLK), .QN(\unit_decode/n1693 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][16]  ( .D(
        \unit_decode/RegisterFile/n2084 ), .CK(CLK), .QN(\unit_decode/n1692 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][15]  ( .D(
        \unit_decode/RegisterFile/n2083 ), .CK(CLK), .QN(\unit_decode/n1691 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][14]  ( .D(
        \unit_decode/RegisterFile/n2082 ), .CK(CLK), .QN(\unit_decode/n1690 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][13]  ( .D(
        \unit_decode/RegisterFile/n2081 ), .CK(CLK), .QN(\unit_decode/n1689 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][12]  ( .D(
        \unit_decode/RegisterFile/n2080 ), .CK(CLK), .QN(\unit_decode/n1688 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][11]  ( .D(
        \unit_decode/RegisterFile/n2079 ), .CK(CLK), .QN(\unit_decode/n1687 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][10]  ( .D(
        \unit_decode/RegisterFile/n2078 ), .CK(CLK), .QN(\unit_decode/n1686 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][9]  ( .D(
        \unit_decode/RegisterFile/n2077 ), .CK(CLK), .QN(\unit_decode/n1685 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][8]  ( .D(
        \unit_decode/RegisterFile/n2076 ), .CK(CLK), .QN(\unit_decode/n1684 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][7]  ( .D(
        \unit_decode/RegisterFile/n2075 ), .CK(CLK), .QN(\unit_decode/n1683 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][6]  ( .D(
        \unit_decode/RegisterFile/n2074 ), .CK(CLK), .QN(\unit_decode/n1682 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][5]  ( .D(
        \unit_decode/RegisterFile/n2073 ), .CK(CLK), .QN(\unit_decode/n1681 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][4]  ( .D(
        \unit_decode/RegisterFile/n2072 ), .CK(CLK), .QN(\unit_decode/n1680 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][3]  ( .D(
        \unit_decode/RegisterFile/n2071 ), .CK(CLK), .QN(\unit_decode/n1679 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][2]  ( .D(
        \unit_decode/RegisterFile/n2070 ), .CK(CLK), .QN(\unit_decode/n1678 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][1]  ( .D(
        \unit_decode/RegisterFile/n2069 ), .CK(CLK), .QN(\unit_decode/n1677 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[2][0]  ( .D(
        \unit_decode/RegisterFile/n2068 ), .CK(CLK), .QN(\unit_decode/n1676 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][23]  ( .D(
        \unit_decode/RegisterFile/n2059 ), .CK(CLK), .QN(\unit_decode/n1675 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][22]  ( .D(
        \unit_decode/RegisterFile/n2058 ), .CK(CLK), .QN(\unit_decode/n1674 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][21]  ( .D(
        \unit_decode/RegisterFile/n2057 ), .CK(CLK), .QN(\unit_decode/n1673 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][20]  ( .D(
        \unit_decode/RegisterFile/n2056 ), .CK(CLK), .QN(\unit_decode/n1672 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][19]  ( .D(
        \unit_decode/RegisterFile/n2055 ), .CK(CLK), .QN(\unit_decode/n1671 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][18]  ( .D(
        \unit_decode/RegisterFile/n2054 ), .CK(CLK), .QN(\unit_decode/n1670 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][17]  ( .D(
        \unit_decode/RegisterFile/n2053 ), .CK(CLK), .QN(\unit_decode/n1669 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][16]  ( .D(
        \unit_decode/RegisterFile/n2052 ), .CK(CLK), .QN(\unit_decode/n1668 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][15]  ( .D(
        \unit_decode/RegisterFile/n2051 ), .CK(CLK), .QN(\unit_decode/n1667 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][14]  ( .D(
        \unit_decode/RegisterFile/n2050 ), .CK(CLK), .QN(\unit_decode/n1666 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][13]  ( .D(
        \unit_decode/RegisterFile/n2049 ), .CK(CLK), .QN(\unit_decode/n1665 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][12]  ( .D(
        \unit_decode/RegisterFile/n2048 ), .CK(CLK), .QN(\unit_decode/n1664 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][11]  ( .D(
        \unit_decode/RegisterFile/n2047 ), .CK(CLK), .QN(\unit_decode/n1663 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][10]  ( .D(
        \unit_decode/RegisterFile/n2046 ), .CK(CLK), .QN(\unit_decode/n1662 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][9]  ( .D(
        \unit_decode/RegisterFile/n2045 ), .CK(CLK), .QN(\unit_decode/n1661 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][8]  ( .D(
        \unit_decode/RegisterFile/n2044 ), .CK(CLK), .QN(\unit_decode/n1660 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][7]  ( .D(
        \unit_decode/RegisterFile/n2043 ), .CK(CLK), .QN(\unit_decode/n1659 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][6]  ( .D(
        \unit_decode/RegisterFile/n2042 ), .CK(CLK), .QN(\unit_decode/n1658 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][5]  ( .D(
        \unit_decode/RegisterFile/n2041 ), .CK(CLK), .QN(\unit_decode/n1657 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][4]  ( .D(
        \unit_decode/RegisterFile/n2040 ), .CK(CLK), .QN(\unit_decode/n1656 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][3]  ( .D(
        \unit_decode/RegisterFile/n2039 ), .CK(CLK), .QN(\unit_decode/n1655 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][2]  ( .D(
        \unit_decode/RegisterFile/n2038 ), .CK(CLK), .QN(\unit_decode/n1654 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][1]  ( .D(
        \unit_decode/RegisterFile/n2037 ), .CK(CLK), .QN(\unit_decode/n1653 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[3][0]  ( .D(
        \unit_decode/RegisterFile/n2036 ), .CK(CLK), .QN(\unit_decode/n1652 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][23]  ( .D(
        \unit_decode/RegisterFile/n2027 ), .CK(CLK), .Q(\unit_decode/n4118 ), 
        .QN(\unit_decode/n1651 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][22]  ( .D(
        \unit_decode/RegisterFile/n2026 ), .CK(CLK), .Q(\unit_decode/n4122 ), 
        .QN(\unit_decode/n1650 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][21]  ( .D(
        \unit_decode/RegisterFile/n2025 ), .CK(CLK), .Q(\unit_decode/n4126 ), 
        .QN(\unit_decode/n1649 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][20]  ( .D(
        \unit_decode/RegisterFile/n2024 ), .CK(CLK), .Q(\unit_decode/n4130 ), 
        .QN(\unit_decode/n1648 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][19]  ( .D(
        \unit_decode/RegisterFile/n2023 ), .CK(CLK), .Q(\unit_decode/n4134 ), 
        .QN(\unit_decode/n1647 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][18]  ( .D(
        \unit_decode/RegisterFile/n2022 ), .CK(CLK), .Q(\unit_decode/n4138 ), 
        .QN(\unit_decode/n1646 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][17]  ( .D(
        \unit_decode/RegisterFile/n2021 ), .CK(CLK), .Q(\unit_decode/n4022 ), 
        .QN(\unit_decode/n1645 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][16]  ( .D(
        \unit_decode/RegisterFile/n2020 ), .CK(CLK), .Q(\unit_decode/n4026 ), 
        .QN(\unit_decode/n1644 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][15]  ( .D(
        \unit_decode/RegisterFile/n2019 ), .CK(CLK), .Q(\unit_decode/n4030 ), 
        .QN(\unit_decode/n1643 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][14]  ( .D(
        \unit_decode/RegisterFile/n2018 ), .CK(CLK), .Q(\unit_decode/n4034 ), 
        .QN(\unit_decode/n1642 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][13]  ( .D(
        \unit_decode/RegisterFile/n2017 ), .CK(CLK), .Q(\unit_decode/n4038 ), 
        .QN(\unit_decode/n1641 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][12]  ( .D(
        \unit_decode/RegisterFile/n2016 ), .CK(CLK), .Q(\unit_decode/n4042 ), 
        .QN(\unit_decode/n1640 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][11]  ( .D(
        \unit_decode/RegisterFile/n2015 ), .CK(CLK), .Q(\unit_decode/n4046 ), 
        .QN(\unit_decode/n1639 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][10]  ( .D(
        \unit_decode/RegisterFile/n2014 ), .CK(CLK), .Q(\unit_decode/n4050 ), 
        .QN(\unit_decode/n1638 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][9]  ( .D(
        \unit_decode/RegisterFile/n2013 ), .CK(CLK), .Q(\unit_decode/n4054 ), 
        .QN(\unit_decode/n1637 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][8]  ( .D(
        \unit_decode/RegisterFile/n2012 ), .CK(CLK), .Q(\unit_decode/n4058 ), 
        .QN(\unit_decode/n1636 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][7]  ( .D(
        \unit_decode/RegisterFile/n2011 ), .CK(CLK), .Q(\unit_decode/n4062 ), 
        .QN(\unit_decode/n1635 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][6]  ( .D(
        \unit_decode/RegisterFile/n2010 ), .CK(CLK), .Q(\unit_decode/n4066 ), 
        .QN(\unit_decode/n1634 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][5]  ( .D(
        \unit_decode/RegisterFile/n2009 ), .CK(CLK), .Q(\unit_decode/n4070 ), 
        .QN(\unit_decode/n1633 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][4]  ( .D(
        \unit_decode/RegisterFile/n2008 ), .CK(CLK), .Q(\unit_decode/n4074 ), 
        .QN(\unit_decode/n1632 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][3]  ( .D(
        \unit_decode/RegisterFile/n2007 ), .CK(CLK), .Q(\unit_decode/n4078 ), 
        .QN(\unit_decode/n1631 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][2]  ( .D(
        \unit_decode/RegisterFile/n2006 ), .CK(CLK), .Q(\unit_decode/n4082 ), 
        .QN(\unit_decode/n1630 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][1]  ( .D(
        \unit_decode/RegisterFile/n2005 ), .CK(CLK), .Q(\unit_decode/n4086 ), 
        .QN(\unit_decode/n1629 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[4][0]  ( .D(
        \unit_decode/RegisterFile/n2004 ), .CK(CLK), .Q(\unit_decode/n4090 ), 
        .QN(\unit_decode/n1628 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][23]  ( .D(
        \unit_decode/RegisterFile/n1995 ), .CK(CLK), .Q(\unit_decode/n3688 ), 
        .QN(\unit_decode/n1627 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][22]  ( .D(
        \unit_decode/RegisterFile/n1994 ), .CK(CLK), .Q(\unit_decode/n3694 ), 
        .QN(\unit_decode/n1626 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][21]  ( .D(
        \unit_decode/RegisterFile/n1993 ), .CK(CLK), .Q(\unit_decode/n3700 ), 
        .QN(\unit_decode/n1625 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][20]  ( .D(
        \unit_decode/RegisterFile/n1992 ), .CK(CLK), .Q(\unit_decode/n3706 ), 
        .QN(\unit_decode/n1624 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][19]  ( .D(
        \unit_decode/RegisterFile/n1991 ), .CK(CLK), .Q(\unit_decode/n3712 ), 
        .QN(\unit_decode/n1623 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][18]  ( .D(
        \unit_decode/RegisterFile/n1990 ), .CK(CLK), .Q(\unit_decode/n3718 ), 
        .QN(\unit_decode/n1622 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][17]  ( .D(
        \unit_decode/RegisterFile/n1989 ), .CK(CLK), .Q(\unit_decode/n3724 ), 
        .QN(\unit_decode/n1621 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][16]  ( .D(
        \unit_decode/RegisterFile/n1988 ), .CK(CLK), .Q(\unit_decode/n3730 ), 
        .QN(\unit_decode/n1620 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][15]  ( .D(
        \unit_decode/RegisterFile/n1987 ), .CK(CLK), .Q(\unit_decode/n3736 ), 
        .QN(\unit_decode/n1619 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][14]  ( .D(
        \unit_decode/RegisterFile/n1986 ), .CK(CLK), .Q(\unit_decode/n3742 ), 
        .QN(\unit_decode/n1618 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][13]  ( .D(
        \unit_decode/RegisterFile/n1985 ), .CK(CLK), .Q(\unit_decode/n3748 ), 
        .QN(\unit_decode/n1617 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][12]  ( .D(
        \unit_decode/RegisterFile/n1984 ), .CK(CLK), .Q(\unit_decode/n3754 ), 
        .QN(\unit_decode/n1616 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][11]  ( .D(
        \unit_decode/RegisterFile/n1983 ), .CK(CLK), .Q(\unit_decode/n3760 ), 
        .QN(\unit_decode/n1615 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][10]  ( .D(
        \unit_decode/RegisterFile/n1982 ), .CK(CLK), .Q(\unit_decode/n3766 ), 
        .QN(\unit_decode/n1614 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][9]  ( .D(
        \unit_decode/RegisterFile/n1981 ), .CK(CLK), .Q(\unit_decode/n3772 ), 
        .QN(\unit_decode/n1613 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][8]  ( .D(
        \unit_decode/RegisterFile/n1980 ), .CK(CLK), .Q(\unit_decode/n3778 ), 
        .QN(\unit_decode/n1612 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][7]  ( .D(
        \unit_decode/RegisterFile/n1979 ), .CK(CLK), .Q(\unit_decode/n3784 ), 
        .QN(\unit_decode/n1611 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][6]  ( .D(
        \unit_decode/RegisterFile/n1978 ), .CK(CLK), .Q(\unit_decode/n3790 ), 
        .QN(\unit_decode/n1610 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][5]  ( .D(
        \unit_decode/RegisterFile/n1977 ), .CK(CLK), .Q(\unit_decode/n3796 ), 
        .QN(\unit_decode/n1609 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][4]  ( .D(
        \unit_decode/RegisterFile/n1976 ), .CK(CLK), .Q(\unit_decode/n3802 ), 
        .QN(\unit_decode/n1608 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][3]  ( .D(
        \unit_decode/RegisterFile/n1975 ), .CK(CLK), .Q(\unit_decode/n3808 ), 
        .QN(\unit_decode/n1607 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][2]  ( .D(
        \unit_decode/RegisterFile/n1974 ), .CK(CLK), .Q(\unit_decode/n3814 ), 
        .QN(\unit_decode/n1606 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][1]  ( .D(
        \unit_decode/RegisterFile/n1973 ), .CK(CLK), .Q(\unit_decode/n3820 ), 
        .QN(\unit_decode/n1605 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[5][0]  ( .D(
        \unit_decode/RegisterFile/n1972 ), .CK(CLK), .Q(\unit_decode/n3826 ), 
        .QN(\unit_decode/n1604 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][23]  ( .D(
        \unit_decode/RegisterFile/n1963 ), .CK(CLK), .QN(\unit_decode/n1603 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][22]  ( .D(
        \unit_decode/RegisterFile/n1962 ), .CK(CLK), .QN(\unit_decode/n1602 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][21]  ( .D(
        \unit_decode/RegisterFile/n1961 ), .CK(CLK), .QN(\unit_decode/n1601 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][20]  ( .D(
        \unit_decode/RegisterFile/n1960 ), .CK(CLK), .QN(\unit_decode/n1600 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][19]  ( .D(
        \unit_decode/RegisterFile/n1959 ), .CK(CLK), .QN(\unit_decode/n1599 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][18]  ( .D(
        \unit_decode/RegisterFile/n1958 ), .CK(CLK), .QN(\unit_decode/n1598 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][17]  ( .D(
        \unit_decode/RegisterFile/n1957 ), .CK(CLK), .QN(\unit_decode/n1597 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][16]  ( .D(
        \unit_decode/RegisterFile/n1956 ), .CK(CLK), .QN(\unit_decode/n1596 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][15]  ( .D(
        \unit_decode/RegisterFile/n1955 ), .CK(CLK), .QN(\unit_decode/n1595 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][14]  ( .D(
        \unit_decode/RegisterFile/n1954 ), .CK(CLK), .QN(\unit_decode/n1594 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][13]  ( .D(
        \unit_decode/RegisterFile/n1953 ), .CK(CLK), .QN(\unit_decode/n1593 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][12]  ( .D(
        \unit_decode/RegisterFile/n1952 ), .CK(CLK), .QN(\unit_decode/n1592 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][11]  ( .D(
        \unit_decode/RegisterFile/n1951 ), .CK(CLK), .QN(\unit_decode/n1591 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][10]  ( .D(
        \unit_decode/RegisterFile/n1950 ), .CK(CLK), .QN(\unit_decode/n1590 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][9]  ( .D(
        \unit_decode/RegisterFile/n1949 ), .CK(CLK), .QN(\unit_decode/n1589 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][8]  ( .D(
        \unit_decode/RegisterFile/n1948 ), .CK(CLK), .QN(\unit_decode/n1588 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][7]  ( .D(
        \unit_decode/RegisterFile/n1947 ), .CK(CLK), .QN(\unit_decode/n1587 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][6]  ( .D(
        \unit_decode/RegisterFile/n1946 ), .CK(CLK), .QN(\unit_decode/n1586 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][5]  ( .D(
        \unit_decode/RegisterFile/n1945 ), .CK(CLK), .QN(\unit_decode/n1585 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][4]  ( .D(
        \unit_decode/RegisterFile/n1944 ), .CK(CLK), .QN(\unit_decode/n1584 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][3]  ( .D(
        \unit_decode/RegisterFile/n1943 ), .CK(CLK), .QN(\unit_decode/n1583 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][2]  ( .D(
        \unit_decode/RegisterFile/n1942 ), .CK(CLK), .QN(\unit_decode/n1582 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][1]  ( .D(
        \unit_decode/RegisterFile/n1941 ), .CK(CLK), .QN(\unit_decode/n1581 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[6][0]  ( .D(
        \unit_decode/RegisterFile/n1940 ), .CK(CLK), .QN(\unit_decode/n1580 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][23]  ( .D(
        \unit_decode/RegisterFile/n1931 ), .CK(CLK), .QN(\unit_decode/n1579 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][22]  ( .D(
        \unit_decode/RegisterFile/n1930 ), .CK(CLK), .QN(\unit_decode/n1578 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][21]  ( .D(
        \unit_decode/RegisterFile/n1929 ), .CK(CLK), .QN(\unit_decode/n1577 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][20]  ( .D(
        \unit_decode/RegisterFile/n1928 ), .CK(CLK), .QN(\unit_decode/n1576 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][19]  ( .D(
        \unit_decode/RegisterFile/n1927 ), .CK(CLK), .QN(\unit_decode/n1575 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][18]  ( .D(
        \unit_decode/RegisterFile/n1926 ), .CK(CLK), .QN(\unit_decode/n1574 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][17]  ( .D(
        \unit_decode/RegisterFile/n1925 ), .CK(CLK), .QN(\unit_decode/n1573 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][16]  ( .D(
        \unit_decode/RegisterFile/n1924 ), .CK(CLK), .QN(\unit_decode/n1572 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][15]  ( .D(
        \unit_decode/RegisterFile/n1923 ), .CK(CLK), .QN(\unit_decode/n1571 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][14]  ( .D(
        \unit_decode/RegisterFile/n1922 ), .CK(CLK), .QN(\unit_decode/n1570 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][13]  ( .D(
        \unit_decode/RegisterFile/n1921 ), .CK(CLK), .QN(\unit_decode/n1569 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][12]  ( .D(
        \unit_decode/RegisterFile/n1920 ), .CK(CLK), .QN(\unit_decode/n1568 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][11]  ( .D(
        \unit_decode/RegisterFile/n1919 ), .CK(CLK), .QN(\unit_decode/n1567 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][10]  ( .D(
        \unit_decode/RegisterFile/n1918 ), .CK(CLK), .QN(\unit_decode/n1566 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][9]  ( .D(
        \unit_decode/RegisterFile/n1917 ), .CK(CLK), .QN(\unit_decode/n1565 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][8]  ( .D(
        \unit_decode/RegisterFile/n1916 ), .CK(CLK), .QN(\unit_decode/n1564 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][7]  ( .D(
        \unit_decode/RegisterFile/n1915 ), .CK(CLK), .QN(\unit_decode/n1563 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][6]  ( .D(
        \unit_decode/RegisterFile/n1914 ), .CK(CLK), .QN(\unit_decode/n1562 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][5]  ( .D(
        \unit_decode/RegisterFile/n1913 ), .CK(CLK), .QN(\unit_decode/n1561 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][4]  ( .D(
        \unit_decode/RegisterFile/n1912 ), .CK(CLK), .QN(\unit_decode/n1560 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][3]  ( .D(
        \unit_decode/RegisterFile/n1911 ), .CK(CLK), .QN(\unit_decode/n1559 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][2]  ( .D(
        \unit_decode/RegisterFile/n1910 ), .CK(CLK), .QN(\unit_decode/n1558 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][1]  ( .D(
        \unit_decode/RegisterFile/n1909 ), .CK(CLK), .QN(\unit_decode/n1557 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[7][0]  ( .D(
        \unit_decode/RegisterFile/n1908 ), .CK(CLK), .QN(\unit_decode/n1556 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][23]  ( .D(
        \unit_decode/RegisterFile/n1899 ), .CK(CLK), .Q(\unit_decode/n4115 ), 
        .QN(\unit_decode/n1555 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][22]  ( .D(
        \unit_decode/RegisterFile/n1898 ), .CK(CLK), .Q(\unit_decode/n4119 ), 
        .QN(\unit_decode/n1554 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][21]  ( .D(
        \unit_decode/RegisterFile/n1897 ), .CK(CLK), .Q(\unit_decode/n4123 ), 
        .QN(\unit_decode/n1553 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][20]  ( .D(
        \unit_decode/RegisterFile/n1896 ), .CK(CLK), .Q(\unit_decode/n4127 ), 
        .QN(\unit_decode/n1552 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][19]  ( .D(
        \unit_decode/RegisterFile/n1895 ), .CK(CLK), .Q(\unit_decode/n4131 ), 
        .QN(\unit_decode/n1551 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][18]  ( .D(
        \unit_decode/RegisterFile/n1894 ), .CK(CLK), .Q(\unit_decode/n4135 ), 
        .QN(\unit_decode/n1550 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][17]  ( .D(
        \unit_decode/RegisterFile/n1893 ), .CK(CLK), .Q(\unit_decode/n4019 ), 
        .QN(\unit_decode/n1549 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][16]  ( .D(
        \unit_decode/RegisterFile/n1892 ), .CK(CLK), .Q(\unit_decode/n4023 ), 
        .QN(\unit_decode/n1548 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][15]  ( .D(
        \unit_decode/RegisterFile/n1891 ), .CK(CLK), .Q(\unit_decode/n4027 ), 
        .QN(\unit_decode/n1547 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][14]  ( .D(
        \unit_decode/RegisterFile/n1890 ), .CK(CLK), .Q(\unit_decode/n4031 ), 
        .QN(\unit_decode/n1546 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][13]  ( .D(
        \unit_decode/RegisterFile/n1889 ), .CK(CLK), .Q(\unit_decode/n4035 ), 
        .QN(\unit_decode/n1545 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][12]  ( .D(
        \unit_decode/RegisterFile/n1888 ), .CK(CLK), .Q(\unit_decode/n4039 ), 
        .QN(\unit_decode/n1544 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][11]  ( .D(
        \unit_decode/RegisterFile/n1887 ), .CK(CLK), .Q(\unit_decode/n4043 ), 
        .QN(\unit_decode/n1543 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][10]  ( .D(
        \unit_decode/RegisterFile/n1886 ), .CK(CLK), .Q(\unit_decode/n4047 ), 
        .QN(\unit_decode/n1542 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][9]  ( .D(
        \unit_decode/RegisterFile/n1885 ), .CK(CLK), .Q(\unit_decode/n4051 ), 
        .QN(\unit_decode/n1541 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][8]  ( .D(
        \unit_decode/RegisterFile/n1884 ), .CK(CLK), .Q(\unit_decode/n4055 ), 
        .QN(\unit_decode/n1540 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][7]  ( .D(
        \unit_decode/RegisterFile/n1883 ), .CK(CLK), .Q(\unit_decode/n4059 ), 
        .QN(\unit_decode/n1539 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][6]  ( .D(
        \unit_decode/RegisterFile/n1882 ), .CK(CLK), .Q(\unit_decode/n4063 ), 
        .QN(\unit_decode/n1538 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][5]  ( .D(
        \unit_decode/RegisterFile/n1881 ), .CK(CLK), .Q(\unit_decode/n4067 ), 
        .QN(\unit_decode/n1537 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][4]  ( .D(
        \unit_decode/RegisterFile/n1880 ), .CK(CLK), .Q(\unit_decode/n4071 ), 
        .QN(\unit_decode/n1536 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][3]  ( .D(
        \unit_decode/RegisterFile/n1879 ), .CK(CLK), .Q(\unit_decode/n4075 ), 
        .QN(\unit_decode/n1535 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][2]  ( .D(
        \unit_decode/RegisterFile/n1878 ), .CK(CLK), .Q(\unit_decode/n4079 ), 
        .QN(\unit_decode/n1534 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][1]  ( .D(
        \unit_decode/RegisterFile/n1877 ), .CK(CLK), .Q(\unit_decode/n4083 ), 
        .QN(\unit_decode/n1533 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[8][0]  ( .D(
        \unit_decode/RegisterFile/n1876 ), .CK(CLK), .Q(\unit_decode/n4087 ), 
        .QN(\unit_decode/n1532 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][23]  ( .D(
        \unit_decode/RegisterFile/n1867 ), .CK(CLK), .Q(\unit_decode/n3867 ), 
        .QN(\unit_decode/n1531 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][22]  ( .D(
        \unit_decode/RegisterFile/n1866 ), .CK(CLK), .Q(\unit_decode/n3873 ), 
        .QN(\unit_decode/n1530 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][21]  ( .D(
        \unit_decode/RegisterFile/n1865 ), .CK(CLK), .Q(\unit_decode/n3879 ), 
        .QN(\unit_decode/n1529 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][20]  ( .D(
        \unit_decode/RegisterFile/n1864 ), .CK(CLK), .Q(\unit_decode/n3885 ), 
        .QN(\unit_decode/n1528 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][19]  ( .D(
        \unit_decode/RegisterFile/n1863 ), .CK(CLK), .Q(\unit_decode/n3891 ), 
        .QN(\unit_decode/n1527 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][18]  ( .D(
        \unit_decode/RegisterFile/n1862 ), .CK(CLK), .Q(\unit_decode/n3897 ), 
        .QN(\unit_decode/n1526 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][17]  ( .D(
        \unit_decode/RegisterFile/n1861 ), .CK(CLK), .Q(\unit_decode/n3903 ), 
        .QN(\unit_decode/n1525 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][16]  ( .D(
        \unit_decode/RegisterFile/n1860 ), .CK(CLK), .Q(\unit_decode/n3909 ), 
        .QN(\unit_decode/n1524 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][15]  ( .D(
        \unit_decode/RegisterFile/n1859 ), .CK(CLK), .Q(\unit_decode/n3915 ), 
        .QN(\unit_decode/n1523 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][14]  ( .D(
        \unit_decode/RegisterFile/n1858 ), .CK(CLK), .Q(\unit_decode/n3921 ), 
        .QN(\unit_decode/n1522 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][13]  ( .D(
        \unit_decode/RegisterFile/n1857 ), .CK(CLK), .Q(\unit_decode/n3927 ), 
        .QN(\unit_decode/n1521 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][12]  ( .D(
        \unit_decode/RegisterFile/n1856 ), .CK(CLK), .Q(\unit_decode/n3933 ), 
        .QN(\unit_decode/n1520 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][11]  ( .D(
        \unit_decode/RegisterFile/n1855 ), .CK(CLK), .Q(\unit_decode/n3939 ), 
        .QN(\unit_decode/n1519 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][10]  ( .D(
        \unit_decode/RegisterFile/n1854 ), .CK(CLK), .Q(\unit_decode/n3945 ), 
        .QN(\unit_decode/n1518 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][9]  ( .D(
        \unit_decode/RegisterFile/n1853 ), .CK(CLK), .Q(\unit_decode/n3951 ), 
        .QN(\unit_decode/n1517 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][8]  ( .D(
        \unit_decode/RegisterFile/n1852 ), .CK(CLK), .Q(\unit_decode/n3957 ), 
        .QN(\unit_decode/n1516 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][7]  ( .D(
        \unit_decode/RegisterFile/n1851 ), .CK(CLK), .Q(\unit_decode/n3963 ), 
        .QN(\unit_decode/n1515 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][6]  ( .D(
        \unit_decode/RegisterFile/n1850 ), .CK(CLK), .Q(\unit_decode/n3969 ), 
        .QN(\unit_decode/n1514 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][5]  ( .D(
        \unit_decode/RegisterFile/n1849 ), .CK(CLK), .Q(\unit_decode/n3975 ), 
        .QN(\unit_decode/n1513 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][4]  ( .D(
        \unit_decode/RegisterFile/n1848 ), .CK(CLK), .Q(\unit_decode/n3981 ), 
        .QN(\unit_decode/n1512 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][3]  ( .D(
        \unit_decode/RegisterFile/n1847 ), .CK(CLK), .Q(\unit_decode/n3987 ), 
        .QN(\unit_decode/n1511 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][2]  ( .D(
        \unit_decode/RegisterFile/n1846 ), .CK(CLK), .Q(\unit_decode/n3993 ), 
        .QN(\unit_decode/n1510 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][1]  ( .D(
        \unit_decode/RegisterFile/n1845 ), .CK(CLK), .Q(\unit_decode/n3999 ), 
        .QN(\unit_decode/n1509 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[9][0]  ( .D(
        \unit_decode/RegisterFile/n1844 ), .CK(CLK), .Q(\unit_decode/n4005 ), 
        .QN(\unit_decode/n1508 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][23]  ( .D(
        \unit_decode/RegisterFile/n1835 ), .CK(CLK), .QN(\unit_decode/n1507 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][22]  ( .D(
        \unit_decode/RegisterFile/n1834 ), .CK(CLK), .QN(\unit_decode/n1506 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][21]  ( .D(
        \unit_decode/RegisterFile/n1833 ), .CK(CLK), .QN(\unit_decode/n1505 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][20]  ( .D(
        \unit_decode/RegisterFile/n1832 ), .CK(CLK), .QN(\unit_decode/n1504 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][19]  ( .D(
        \unit_decode/RegisterFile/n1831 ), .CK(CLK), .QN(\unit_decode/n1503 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][18]  ( .D(
        \unit_decode/RegisterFile/n1830 ), .CK(CLK), .QN(\unit_decode/n1502 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][17]  ( .D(
        \unit_decode/RegisterFile/n1829 ), .CK(CLK), .QN(\unit_decode/n1501 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][16]  ( .D(
        \unit_decode/RegisterFile/n1828 ), .CK(CLK), .QN(\unit_decode/n1500 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][15]  ( .D(
        \unit_decode/RegisterFile/n1827 ), .CK(CLK), .QN(\unit_decode/n1499 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][14]  ( .D(
        \unit_decode/RegisterFile/n1826 ), .CK(CLK), .QN(\unit_decode/n1498 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][13]  ( .D(
        \unit_decode/RegisterFile/n1825 ), .CK(CLK), .QN(\unit_decode/n1497 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][12]  ( .D(
        \unit_decode/RegisterFile/n1824 ), .CK(CLK), .QN(\unit_decode/n1496 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][11]  ( .D(
        \unit_decode/RegisterFile/n1823 ), .CK(CLK), .QN(\unit_decode/n1495 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][10]  ( .D(
        \unit_decode/RegisterFile/n1822 ), .CK(CLK), .QN(\unit_decode/n1494 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][9]  ( .D(
        \unit_decode/RegisterFile/n1821 ), .CK(CLK), .QN(\unit_decode/n1493 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][8]  ( .D(
        \unit_decode/RegisterFile/n1820 ), .CK(CLK), .QN(\unit_decode/n1492 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][7]  ( .D(
        \unit_decode/RegisterFile/n1819 ), .CK(CLK), .QN(\unit_decode/n1491 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][6]  ( .D(
        \unit_decode/RegisterFile/n1818 ), .CK(CLK), .QN(\unit_decode/n1490 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][5]  ( .D(
        \unit_decode/RegisterFile/n1817 ), .CK(CLK), .QN(\unit_decode/n1489 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][4]  ( .D(
        \unit_decode/RegisterFile/n1816 ), .CK(CLK), .QN(\unit_decode/n1488 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][3]  ( .D(
        \unit_decode/RegisterFile/n1815 ), .CK(CLK), .QN(\unit_decode/n1487 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][2]  ( .D(
        \unit_decode/RegisterFile/n1814 ), .CK(CLK), .QN(\unit_decode/n1486 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][1]  ( .D(
        \unit_decode/RegisterFile/n1813 ), .CK(CLK), .QN(\unit_decode/n1485 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[10][0]  ( .D(
        \unit_decode/RegisterFile/n1812 ), .CK(CLK), .QN(\unit_decode/n1484 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][23]  ( .D(
        \unit_decode/RegisterFile/n1803 ), .CK(CLK), .QN(\unit_decode/n1483 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][22]  ( .D(
        \unit_decode/RegisterFile/n1802 ), .CK(CLK), .QN(\unit_decode/n1482 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][21]  ( .D(
        \unit_decode/RegisterFile/n1801 ), .CK(CLK), .QN(\unit_decode/n1481 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][20]  ( .D(
        \unit_decode/RegisterFile/n1800 ), .CK(CLK), .QN(\unit_decode/n1480 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][19]  ( .D(
        \unit_decode/RegisterFile/n1799 ), .CK(CLK), .QN(\unit_decode/n1479 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][18]  ( .D(
        \unit_decode/RegisterFile/n1798 ), .CK(CLK), .QN(\unit_decode/n1478 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][17]  ( .D(
        \unit_decode/RegisterFile/n1797 ), .CK(CLK), .QN(\unit_decode/n1477 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][16]  ( .D(
        \unit_decode/RegisterFile/n1796 ), .CK(CLK), .QN(\unit_decode/n1476 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][15]  ( .D(
        \unit_decode/RegisterFile/n1795 ), .CK(CLK), .QN(\unit_decode/n1475 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][14]  ( .D(
        \unit_decode/RegisterFile/n1794 ), .CK(CLK), .QN(\unit_decode/n1474 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][13]  ( .D(
        \unit_decode/RegisterFile/n1793 ), .CK(CLK), .QN(\unit_decode/n1473 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][12]  ( .D(
        \unit_decode/RegisterFile/n1792 ), .CK(CLK), .QN(\unit_decode/n1472 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][11]  ( .D(
        \unit_decode/RegisterFile/n1791 ), .CK(CLK), .QN(\unit_decode/n1471 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][10]  ( .D(
        \unit_decode/RegisterFile/n1790 ), .CK(CLK), .QN(\unit_decode/n1470 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][9]  ( .D(
        \unit_decode/RegisterFile/n1789 ), .CK(CLK), .QN(\unit_decode/n1469 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][8]  ( .D(
        \unit_decode/RegisterFile/n1788 ), .CK(CLK), .QN(\unit_decode/n1468 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][7]  ( .D(
        \unit_decode/RegisterFile/n1787 ), .CK(CLK), .QN(\unit_decode/n1467 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][6]  ( .D(
        \unit_decode/RegisterFile/n1786 ), .CK(CLK), .QN(\unit_decode/n1466 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][5]  ( .D(
        \unit_decode/RegisterFile/n1785 ), .CK(CLK), .QN(\unit_decode/n1465 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][4]  ( .D(
        \unit_decode/RegisterFile/n1784 ), .CK(CLK), .QN(\unit_decode/n1464 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][3]  ( .D(
        \unit_decode/RegisterFile/n1783 ), .CK(CLK), .QN(\unit_decode/n1463 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][2]  ( .D(
        \unit_decode/RegisterFile/n1782 ), .CK(CLK), .QN(\unit_decode/n1462 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][1]  ( .D(
        \unit_decode/RegisterFile/n1781 ), .CK(CLK), .QN(\unit_decode/n1461 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[11][0]  ( .D(
        \unit_decode/RegisterFile/n1780 ), .CK(CLK), .QN(\unit_decode/n1460 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][23]  ( .D(
        \unit_decode/RegisterFile/n1771 ), .CK(CLK), .Q(\unit_decode/n4117 ), 
        .QN(\unit_decode/n1459 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][22]  ( .D(
        \unit_decode/RegisterFile/n1770 ), .CK(CLK), .Q(\unit_decode/n4121 ), 
        .QN(\unit_decode/n1458 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][21]  ( .D(
        \unit_decode/RegisterFile/n1769 ), .CK(CLK), .Q(\unit_decode/n4125 ), 
        .QN(\unit_decode/n1457 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][20]  ( .D(
        \unit_decode/RegisterFile/n1768 ), .CK(CLK), .Q(\unit_decode/n4129 ), 
        .QN(\unit_decode/n1456 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][19]  ( .D(
        \unit_decode/RegisterFile/n1767 ), .CK(CLK), .Q(\unit_decode/n4133 ), 
        .QN(\unit_decode/n1455 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][18]  ( .D(
        \unit_decode/RegisterFile/n1766 ), .CK(CLK), .Q(\unit_decode/n4137 ), 
        .QN(\unit_decode/n1454 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][17]  ( .D(
        \unit_decode/RegisterFile/n1765 ), .CK(CLK), .Q(\unit_decode/n4021 ), 
        .QN(\unit_decode/n1453 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][16]  ( .D(
        \unit_decode/RegisterFile/n1764 ), .CK(CLK), .Q(\unit_decode/n4025 ), 
        .QN(\unit_decode/n1452 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][15]  ( .D(
        \unit_decode/RegisterFile/n1763 ), .CK(CLK), .Q(\unit_decode/n4029 ), 
        .QN(\unit_decode/n1451 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][14]  ( .D(
        \unit_decode/RegisterFile/n1762 ), .CK(CLK), .Q(\unit_decode/n4033 ), 
        .QN(\unit_decode/n1450 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][13]  ( .D(
        \unit_decode/RegisterFile/n1761 ), .CK(CLK), .Q(\unit_decode/n4037 ), 
        .QN(\unit_decode/n1449 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][12]  ( .D(
        \unit_decode/RegisterFile/n1760 ), .CK(CLK), .Q(\unit_decode/n4041 ), 
        .QN(\unit_decode/n1448 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][11]  ( .D(
        \unit_decode/RegisterFile/n1759 ), .CK(CLK), .Q(\unit_decode/n4045 ), 
        .QN(\unit_decode/n1447 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][10]  ( .D(
        \unit_decode/RegisterFile/n1758 ), .CK(CLK), .Q(\unit_decode/n4049 ), 
        .QN(\unit_decode/n1446 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][9]  ( .D(
        \unit_decode/RegisterFile/n1757 ), .CK(CLK), .Q(\unit_decode/n4053 ), 
        .QN(\unit_decode/n1445 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][8]  ( .D(
        \unit_decode/RegisterFile/n1756 ), .CK(CLK), .Q(\unit_decode/n4057 ), 
        .QN(\unit_decode/n1444 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][7]  ( .D(
        \unit_decode/RegisterFile/n1755 ), .CK(CLK), .Q(\unit_decode/n4061 ), 
        .QN(\unit_decode/n1443 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][6]  ( .D(
        \unit_decode/RegisterFile/n1754 ), .CK(CLK), .Q(\unit_decode/n4065 ), 
        .QN(\unit_decode/n1442 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][5]  ( .D(
        \unit_decode/RegisterFile/n1753 ), .CK(CLK), .Q(\unit_decode/n4069 ), 
        .QN(\unit_decode/n1441 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][4]  ( .D(
        \unit_decode/RegisterFile/n1752 ), .CK(CLK), .Q(\unit_decode/n4073 ), 
        .QN(\unit_decode/n1440 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][3]  ( .D(
        \unit_decode/RegisterFile/n1751 ), .CK(CLK), .Q(\unit_decode/n4077 ), 
        .QN(\unit_decode/n1439 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][2]  ( .D(
        \unit_decode/RegisterFile/n1750 ), .CK(CLK), .Q(\unit_decode/n4081 ), 
        .QN(\unit_decode/n1438 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][1]  ( .D(
        \unit_decode/RegisterFile/n1749 ), .CK(CLK), .Q(\unit_decode/n4085 ), 
        .QN(\unit_decode/n1437 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[12][0]  ( .D(
        \unit_decode/RegisterFile/n1748 ), .CK(CLK), .Q(\unit_decode/n4089 ), 
        .QN(\unit_decode/n1436 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][23]  ( .D(
        \unit_decode/RegisterFile/n1739 ), .CK(CLK), .Q(\unit_decode/n3687 ), 
        .QN(\unit_decode/n1435 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][22]  ( .D(
        \unit_decode/RegisterFile/n1738 ), .CK(CLK), .Q(\unit_decode/n3693 ), 
        .QN(\unit_decode/n1434 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][21]  ( .D(
        \unit_decode/RegisterFile/n1737 ), .CK(CLK), .Q(\unit_decode/n3699 ), 
        .QN(\unit_decode/n1433 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][20]  ( .D(
        \unit_decode/RegisterFile/n1736 ), .CK(CLK), .Q(\unit_decode/n3705 ), 
        .QN(\unit_decode/n1432 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][19]  ( .D(
        \unit_decode/RegisterFile/n1735 ), .CK(CLK), .Q(\unit_decode/n3711 ), 
        .QN(\unit_decode/n1431 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][18]  ( .D(
        \unit_decode/RegisterFile/n1734 ), .CK(CLK), .Q(\unit_decode/n3717 ), 
        .QN(\unit_decode/n1430 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][17]  ( .D(
        \unit_decode/RegisterFile/n1733 ), .CK(CLK), .Q(\unit_decode/n3723 ), 
        .QN(\unit_decode/n1429 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][16]  ( .D(
        \unit_decode/RegisterFile/n1732 ), .CK(CLK), .Q(\unit_decode/n3729 ), 
        .QN(\unit_decode/n1428 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][15]  ( .D(
        \unit_decode/RegisterFile/n1731 ), .CK(CLK), .Q(\unit_decode/n3735 ), 
        .QN(\unit_decode/n1427 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][14]  ( .D(
        \unit_decode/RegisterFile/n1730 ), .CK(CLK), .Q(\unit_decode/n3741 ), 
        .QN(\unit_decode/n1426 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][13]  ( .D(
        \unit_decode/RegisterFile/n1729 ), .CK(CLK), .Q(\unit_decode/n3747 ), 
        .QN(\unit_decode/n1425 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][12]  ( .D(
        \unit_decode/RegisterFile/n1728 ), .CK(CLK), .Q(\unit_decode/n3753 ), 
        .QN(\unit_decode/n1424 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][11]  ( .D(
        \unit_decode/RegisterFile/n1727 ), .CK(CLK), .Q(\unit_decode/n3759 ), 
        .QN(\unit_decode/n1423 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][10]  ( .D(
        \unit_decode/RegisterFile/n1726 ), .CK(CLK), .Q(\unit_decode/n3765 ), 
        .QN(\unit_decode/n1422 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][9]  ( .D(
        \unit_decode/RegisterFile/n1725 ), .CK(CLK), .Q(\unit_decode/n3771 ), 
        .QN(\unit_decode/n1421 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][8]  ( .D(
        \unit_decode/RegisterFile/n1724 ), .CK(CLK), .Q(\unit_decode/n3777 ), 
        .QN(\unit_decode/n1420 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][7]  ( .D(
        \unit_decode/RegisterFile/n1723 ), .CK(CLK), .Q(\unit_decode/n3783 ), 
        .QN(\unit_decode/n1419 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][6]  ( .D(
        \unit_decode/RegisterFile/n1722 ), .CK(CLK), .Q(\unit_decode/n3789 ), 
        .QN(\unit_decode/n1418 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][5]  ( .D(
        \unit_decode/RegisterFile/n1721 ), .CK(CLK), .Q(\unit_decode/n3795 ), 
        .QN(\unit_decode/n1417 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][4]  ( .D(
        \unit_decode/RegisterFile/n1720 ), .CK(CLK), .Q(\unit_decode/n3801 ), 
        .QN(\unit_decode/n1416 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][3]  ( .D(
        \unit_decode/RegisterFile/n1719 ), .CK(CLK), .Q(\unit_decode/n3807 ), 
        .QN(\unit_decode/n1415 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][2]  ( .D(
        \unit_decode/RegisterFile/n1718 ), .CK(CLK), .Q(\unit_decode/n3813 ), 
        .QN(\unit_decode/n1414 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][1]  ( .D(
        \unit_decode/RegisterFile/n1717 ), .CK(CLK), .Q(\unit_decode/n3819 ), 
        .QN(\unit_decode/n1413 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[13][0]  ( .D(
        \unit_decode/RegisterFile/n1716 ), .CK(CLK), .Q(\unit_decode/n3825 ), 
        .QN(\unit_decode/n1412 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][23]  ( .D(
        \unit_decode/RegisterFile/n1707 ), .CK(CLK), .QN(\unit_decode/n1411 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][22]  ( .D(
        \unit_decode/RegisterFile/n1706 ), .CK(CLK), .QN(\unit_decode/n1410 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][21]  ( .D(
        \unit_decode/RegisterFile/n1705 ), .CK(CLK), .QN(\unit_decode/n1409 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][20]  ( .D(
        \unit_decode/RegisterFile/n1704 ), .CK(CLK), .QN(\unit_decode/n1408 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][19]  ( .D(
        \unit_decode/RegisterFile/n1703 ), .CK(CLK), .QN(\unit_decode/n1407 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][18]  ( .D(
        \unit_decode/RegisterFile/n1702 ), .CK(CLK), .QN(\unit_decode/n1406 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][17]  ( .D(
        \unit_decode/RegisterFile/n1701 ), .CK(CLK), .QN(\unit_decode/n1405 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][16]  ( .D(
        \unit_decode/RegisterFile/n1700 ), .CK(CLK), .QN(\unit_decode/n1404 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][15]  ( .D(
        \unit_decode/RegisterFile/n1699 ), .CK(CLK), .QN(\unit_decode/n1403 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][14]  ( .D(
        \unit_decode/RegisterFile/n1698 ), .CK(CLK), .QN(\unit_decode/n1402 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][13]  ( .D(
        \unit_decode/RegisterFile/n1697 ), .CK(CLK), .QN(\unit_decode/n1401 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][12]  ( .D(
        \unit_decode/RegisterFile/n1696 ), .CK(CLK), .QN(\unit_decode/n1400 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][11]  ( .D(
        \unit_decode/RegisterFile/n1695 ), .CK(CLK), .QN(\unit_decode/n1399 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][10]  ( .D(
        \unit_decode/RegisterFile/n1694 ), .CK(CLK), .QN(\unit_decode/n1398 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][9]  ( .D(
        \unit_decode/RegisterFile/n1693 ), .CK(CLK), .QN(\unit_decode/n1397 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][8]  ( .D(
        \unit_decode/RegisterFile/n1692 ), .CK(CLK), .QN(\unit_decode/n1396 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][7]  ( .D(
        \unit_decode/RegisterFile/n1691 ), .CK(CLK), .QN(\unit_decode/n1395 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][6]  ( .D(
        \unit_decode/RegisterFile/n1690 ), .CK(CLK), .QN(\unit_decode/n1394 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][5]  ( .D(
        \unit_decode/RegisterFile/n1689 ), .CK(CLK), .QN(\unit_decode/n1393 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][4]  ( .D(
        \unit_decode/RegisterFile/n1688 ), .CK(CLK), .QN(\unit_decode/n1392 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][3]  ( .D(
        \unit_decode/RegisterFile/n1687 ), .CK(CLK), .QN(\unit_decode/n1391 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][2]  ( .D(
        \unit_decode/RegisterFile/n1686 ), .CK(CLK), .QN(\unit_decode/n1390 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][1]  ( .D(
        \unit_decode/RegisterFile/n1685 ), .CK(CLK), .QN(\unit_decode/n1389 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[14][0]  ( .D(
        \unit_decode/RegisterFile/n1684 ), .CK(CLK), .QN(\unit_decode/n1388 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][22]  ( .D(
        \unit_decode/RegisterFile/n1674 ), .CK(CLK), .QN(\unit_decode/n1387 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][21]  ( .D(
        \unit_decode/RegisterFile/n1673 ), .CK(CLK), .QN(\unit_decode/n1386 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][20]  ( .D(
        \unit_decode/RegisterFile/n1672 ), .CK(CLK), .QN(\unit_decode/n1385 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][19]  ( .D(
        \unit_decode/RegisterFile/n1671 ), .CK(CLK), .QN(\unit_decode/n1384 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][18]  ( .D(
        \unit_decode/RegisterFile/n1670 ), .CK(CLK), .QN(\unit_decode/n1383 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][17]  ( .D(
        \unit_decode/RegisterFile/n1669 ), .CK(CLK), .QN(\unit_decode/n1382 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][16]  ( .D(
        \unit_decode/RegisterFile/n1668 ), .CK(CLK), .QN(\unit_decode/n1381 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][15]  ( .D(
        \unit_decode/RegisterFile/n1667 ), .CK(CLK), .QN(\unit_decode/n1380 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][14]  ( .D(
        \unit_decode/RegisterFile/n1666 ), .CK(CLK), .QN(\unit_decode/n1379 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][13]  ( .D(
        \unit_decode/RegisterFile/n1665 ), .CK(CLK), .QN(\unit_decode/n1378 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][12]  ( .D(
        \unit_decode/RegisterFile/n1664 ), .CK(CLK), .QN(\unit_decode/n1377 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][11]  ( .D(
        \unit_decode/RegisterFile/n1663 ), .CK(CLK), .QN(\unit_decode/n1376 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][10]  ( .D(
        \unit_decode/RegisterFile/n1662 ), .CK(CLK), .QN(\unit_decode/n1375 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][9]  ( .D(
        \unit_decode/RegisterFile/n1661 ), .CK(CLK), .QN(\unit_decode/n1374 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][8]  ( .D(
        \unit_decode/RegisterFile/n1660 ), .CK(CLK), .QN(\unit_decode/n1373 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][7]  ( .D(
        \unit_decode/RegisterFile/n1659 ), .CK(CLK), .QN(\unit_decode/n1372 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][6]  ( .D(
        \unit_decode/RegisterFile/n1658 ), .CK(CLK), .QN(\unit_decode/n1371 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][5]  ( .D(
        \unit_decode/RegisterFile/n1657 ), .CK(CLK), .QN(\unit_decode/n1370 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][4]  ( .D(
        \unit_decode/RegisterFile/n1656 ), .CK(CLK), .QN(\unit_decode/n1369 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][3]  ( .D(
        \unit_decode/RegisterFile/n1655 ), .CK(CLK), .QN(\unit_decode/n1368 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][2]  ( .D(
        \unit_decode/RegisterFile/n1654 ), .CK(CLK), .QN(\unit_decode/n1367 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][1]  ( .D(
        \unit_decode/RegisterFile/n1653 ), .CK(CLK), .QN(\unit_decode/n1366 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[15][0]  ( .D(
        \unit_decode/RegisterFile/n1652 ), .CK(CLK), .QN(\unit_decode/n1365 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][23]  ( .D(
        \unit_decode/RegisterFile/n1387 ), .CK(CLK), .Q(\unit_decode/n187 ), 
        .QN(\unit_decode/n1364 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][22]  ( .D(
        \unit_decode/RegisterFile/n1386 ), .CK(CLK), .Q(\unit_decode/n188 ), 
        .QN(\unit_decode/n1363 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][21]  ( .D(
        \unit_decode/RegisterFile/n1385 ), .CK(CLK), .Q(\unit_decode/n189 ), 
        .QN(\unit_decode/n1362 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][20]  ( .D(
        \unit_decode/RegisterFile/n1384 ), .CK(CLK), .Q(\unit_decode/n190 ), 
        .QN(\unit_decode/n1361 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][19]  ( .D(
        \unit_decode/RegisterFile/n1383 ), .CK(CLK), .Q(\unit_decode/n191 ), 
        .QN(\unit_decode/n1360 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][18]  ( .D(
        \unit_decode/RegisterFile/n1382 ), .CK(CLK), .Q(\unit_decode/n192 ), 
        .QN(\unit_decode/n1359 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][17]  ( .D(
        \unit_decode/RegisterFile/n1381 ), .CK(CLK), .Q(\unit_decode/n169 ), 
        .QN(\unit_decode/n1358 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][16]  ( .D(
        \unit_decode/RegisterFile/n1380 ), .CK(CLK), .Q(\unit_decode/n170 ), 
        .QN(\unit_decode/n1357 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][15]  ( .D(
        \unit_decode/RegisterFile/n1379 ), .CK(CLK), .Q(\unit_decode/n171 ), 
        .QN(\unit_decode/n1356 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][14]  ( .D(
        \unit_decode/RegisterFile/n1378 ), .CK(CLK), .Q(\unit_decode/n172 ), 
        .QN(\unit_decode/n1355 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][13]  ( .D(
        \unit_decode/RegisterFile/n1377 ), .CK(CLK), .Q(\unit_decode/n173 ), 
        .QN(\unit_decode/n1354 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][12]  ( .D(
        \unit_decode/RegisterFile/n1376 ), .CK(CLK), .Q(\unit_decode/n174 ), 
        .QN(\unit_decode/n1353 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][11]  ( .D(
        \unit_decode/RegisterFile/n1375 ), .CK(CLK), .Q(\unit_decode/n175 ), 
        .QN(\unit_decode/n1352 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][10]  ( .D(
        \unit_decode/RegisterFile/n1374 ), .CK(CLK), .Q(\unit_decode/n176 ), 
        .QN(\unit_decode/n1351 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][9]  ( .D(
        \unit_decode/RegisterFile/n1373 ), .CK(CLK), .Q(\unit_decode/n177 ), 
        .QN(\unit_decode/n1350 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][8]  ( .D(
        \unit_decode/RegisterFile/n1372 ), .CK(CLK), .Q(\unit_decode/n178 ), 
        .QN(\unit_decode/n1349 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][7]  ( .D(
        \unit_decode/RegisterFile/n1371 ), .CK(CLK), .Q(\unit_decode/n179 ), 
        .QN(\unit_decode/n1348 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][6]  ( .D(
        \unit_decode/RegisterFile/n1370 ), .CK(CLK), .Q(\unit_decode/n180 ), 
        .QN(\unit_decode/n1347 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][5]  ( .D(
        \unit_decode/RegisterFile/n1369 ), .CK(CLK), .Q(\unit_decode/n181 ), 
        .QN(\unit_decode/n1346 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][4]  ( .D(
        \unit_decode/RegisterFile/n1368 ), .CK(CLK), .Q(\unit_decode/n182 ), 
        .QN(\unit_decode/n1345 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][3]  ( .D(
        \unit_decode/RegisterFile/n1367 ), .CK(CLK), .Q(\unit_decode/n183 ), 
        .QN(\unit_decode/n1344 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][2]  ( .D(
        \unit_decode/RegisterFile/n1366 ), .CK(CLK), .Q(\unit_decode/n184 ), 
        .QN(\unit_decode/n1343 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][1]  ( .D(
        \unit_decode/RegisterFile/n1365 ), .CK(CLK), .Q(\unit_decode/n185 ), 
        .QN(\unit_decode/n1342 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][0]  ( .D(
        \unit_decode/RegisterFile/n1364 ), .CK(CLK), .Q(\unit_decode/n186 ), 
        .QN(\unit_decode/n1341 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][23]  ( .D(
        \unit_decode/RegisterFile/n1355 ), .CK(CLK), .Q(\unit_decode/n97 ), 
        .QN(\unit_decode/n1340 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][22]  ( .D(
        \unit_decode/RegisterFile/n1354 ), .CK(CLK), .Q(\unit_decode/n100 ), 
        .QN(\unit_decode/n1339 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][21]  ( .D(
        \unit_decode/RegisterFile/n1353 ), .CK(CLK), .Q(\unit_decode/n103 ), 
        .QN(\unit_decode/n1338 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][20]  ( .D(
        \unit_decode/RegisterFile/n1352 ), .CK(CLK), .Q(\unit_decode/n106 ), 
        .QN(\unit_decode/n1337 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][19]  ( .D(
        \unit_decode/RegisterFile/n1351 ), .CK(CLK), .Q(\unit_decode/n109 ), 
        .QN(\unit_decode/n1336 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][18]  ( .D(
        \unit_decode/RegisterFile/n1350 ), .CK(CLK), .Q(\unit_decode/n112 ), 
        .QN(\unit_decode/n1335 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][17]  ( .D(
        \unit_decode/RegisterFile/n1349 ), .CK(CLK), .Q(\unit_decode/n115 ), 
        .QN(\unit_decode/n1334 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][16]  ( .D(
        \unit_decode/RegisterFile/n1348 ), .CK(CLK), .Q(\unit_decode/n118 ), 
        .QN(\unit_decode/n1333 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][15]  ( .D(
        \unit_decode/RegisterFile/n1347 ), .CK(CLK), .Q(\unit_decode/n121 ), 
        .QN(\unit_decode/n1332 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][14]  ( .D(
        \unit_decode/RegisterFile/n1346 ), .CK(CLK), .Q(\unit_decode/n124 ), 
        .QN(\unit_decode/n1331 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][13]  ( .D(
        \unit_decode/RegisterFile/n1345 ), .CK(CLK), .Q(\unit_decode/n127 ), 
        .QN(\unit_decode/n1330 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][12]  ( .D(
        \unit_decode/RegisterFile/n1344 ), .CK(CLK), .Q(\unit_decode/n130 ), 
        .QN(\unit_decode/n1329 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][11]  ( .D(
        \unit_decode/RegisterFile/n1343 ), .CK(CLK), .Q(\unit_decode/n133 ), 
        .QN(\unit_decode/n1328 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][10]  ( .D(
        \unit_decode/RegisterFile/n1342 ), .CK(CLK), .Q(\unit_decode/n136 ), 
        .QN(\unit_decode/n1327 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][9]  ( .D(
        \unit_decode/RegisterFile/n1341 ), .CK(CLK), .Q(\unit_decode/n139 ), 
        .QN(\unit_decode/n1326 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][8]  ( .D(
        \unit_decode/RegisterFile/n1340 ), .CK(CLK), .Q(\unit_decode/n142 ), 
        .QN(\unit_decode/n1325 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][7]  ( .D(
        \unit_decode/RegisterFile/n1339 ), .CK(CLK), .Q(\unit_decode/n145 ), 
        .QN(\unit_decode/n1324 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][6]  ( .D(
        \unit_decode/RegisterFile/n1338 ), .CK(CLK), .Q(\unit_decode/n148 ), 
        .QN(\unit_decode/n1323 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][5]  ( .D(
        \unit_decode/RegisterFile/n1337 ), .CK(CLK), .Q(\unit_decode/n151 ), 
        .QN(\unit_decode/n1322 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][4]  ( .D(
        \unit_decode/RegisterFile/n1336 ), .CK(CLK), .Q(\unit_decode/n154 ), 
        .QN(\unit_decode/n1321 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][3]  ( .D(
        \unit_decode/RegisterFile/n1335 ), .CK(CLK), .Q(\unit_decode/n157 ), 
        .QN(\unit_decode/n1320 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][2]  ( .D(
        \unit_decode/RegisterFile/n1334 ), .CK(CLK), .Q(\unit_decode/n160 ), 
        .QN(\unit_decode/n1319 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][1]  ( .D(
        \unit_decode/RegisterFile/n1333 ), .CK(CLK), .Q(\unit_decode/n163 ), 
        .QN(\unit_decode/n1318 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][0]  ( .D(
        \unit_decode/RegisterFile/n1332 ), .CK(CLK), .Q(\unit_decode/n166 ), 
        .QN(\unit_decode/n1317 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][23]  ( .D(
        \unit_decode/RegisterFile/n1323 ), .CK(CLK), .QN(\unit_decode/n1316 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][22]  ( .D(
        \unit_decode/RegisterFile/n1322 ), .CK(CLK), .QN(\unit_decode/n1315 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][21]  ( .D(
        \unit_decode/RegisterFile/n1321 ), .CK(CLK), .QN(\unit_decode/n1314 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][20]  ( .D(
        \unit_decode/RegisterFile/n1320 ), .CK(CLK), .QN(\unit_decode/n1313 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][19]  ( .D(
        \unit_decode/RegisterFile/n1319 ), .CK(CLK), .QN(\unit_decode/n1312 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][18]  ( .D(
        \unit_decode/RegisterFile/n1318 ), .CK(CLK), .QN(\unit_decode/n1311 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][17]  ( .D(
        \unit_decode/RegisterFile/n1317 ), .CK(CLK), .QN(\unit_decode/n1310 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][16]  ( .D(
        \unit_decode/RegisterFile/n1316 ), .CK(CLK), .QN(\unit_decode/n1309 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][15]  ( .D(
        \unit_decode/RegisterFile/n1315 ), .CK(CLK), .QN(\unit_decode/n1308 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][14]  ( .D(
        \unit_decode/RegisterFile/n1314 ), .CK(CLK), .QN(\unit_decode/n1307 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][13]  ( .D(
        \unit_decode/RegisterFile/n1313 ), .CK(CLK), .QN(\unit_decode/n1306 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][12]  ( .D(
        \unit_decode/RegisterFile/n1312 ), .CK(CLK), .QN(\unit_decode/n1305 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][11]  ( .D(
        \unit_decode/RegisterFile/n1311 ), .CK(CLK), .QN(\unit_decode/n1304 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][10]  ( .D(
        \unit_decode/RegisterFile/n1310 ), .CK(CLK), .QN(\unit_decode/n1303 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][9]  ( .D(
        \unit_decode/RegisterFile/n1309 ), .CK(CLK), .QN(\unit_decode/n1302 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][8]  ( .D(
        \unit_decode/RegisterFile/n1308 ), .CK(CLK), .QN(\unit_decode/n1301 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][7]  ( .D(
        \unit_decode/RegisterFile/n1307 ), .CK(CLK), .QN(\unit_decode/n1300 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][6]  ( .D(
        \unit_decode/RegisterFile/n1306 ), .CK(CLK), .QN(\unit_decode/n1299 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][5]  ( .D(
        \unit_decode/RegisterFile/n1305 ), .CK(CLK), .QN(\unit_decode/n1298 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][4]  ( .D(
        \unit_decode/RegisterFile/n1304 ), .CK(CLK), .QN(\unit_decode/n1297 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][3]  ( .D(
        \unit_decode/RegisterFile/n1303 ), .CK(CLK), .QN(\unit_decode/n1296 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][2]  ( .D(
        \unit_decode/RegisterFile/n1302 ), .CK(CLK), .QN(\unit_decode/n1295 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][1]  ( .D(
        \unit_decode/RegisterFile/n1301 ), .CK(CLK), .QN(\unit_decode/n1294 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][0]  ( .D(
        \unit_decode/RegisterFile/n1300 ), .CK(CLK), .QN(\unit_decode/n1293 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][23]  ( .D(
        \unit_decode/RegisterFile/n1291 ), .CK(CLK), .QN(\unit_decode/n1292 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][22]  ( .D(
        \unit_decode/RegisterFile/n1290 ), .CK(CLK), .QN(\unit_decode/n1291 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][21]  ( .D(
        \unit_decode/RegisterFile/n1289 ), .CK(CLK), .QN(\unit_decode/n1290 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][20]  ( .D(
        \unit_decode/RegisterFile/n1288 ), .CK(CLK), .QN(\unit_decode/n1289 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][19]  ( .D(
        \unit_decode/RegisterFile/n1287 ), .CK(CLK), .QN(\unit_decode/n1288 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][18]  ( .D(
        \unit_decode/RegisterFile/n1286 ), .CK(CLK), .QN(\unit_decode/n1287 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][17]  ( .D(
        \unit_decode/RegisterFile/n1285 ), .CK(CLK), .QN(\unit_decode/n1286 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][16]  ( .D(
        \unit_decode/RegisterFile/n1284 ), .CK(CLK), .QN(\unit_decode/n1285 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][15]  ( .D(
        \unit_decode/RegisterFile/n1283 ), .CK(CLK), .QN(\unit_decode/n1284 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][14]  ( .D(
        \unit_decode/RegisterFile/n1282 ), .CK(CLK), .QN(\unit_decode/n1283 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][13]  ( .D(
        \unit_decode/RegisterFile/n1281 ), .CK(CLK), .QN(\unit_decode/n1282 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][12]  ( .D(
        \unit_decode/RegisterFile/n1280 ), .CK(CLK), .QN(\unit_decode/n1281 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][11]  ( .D(
        \unit_decode/RegisterFile/n1279 ), .CK(CLK), .QN(\unit_decode/n1280 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][10]  ( .D(
        \unit_decode/RegisterFile/n1278 ), .CK(CLK), .QN(\unit_decode/n1279 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][9]  ( .D(
        \unit_decode/RegisterFile/n1277 ), .CK(CLK), .QN(\unit_decode/n1278 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][8]  ( .D(
        \unit_decode/RegisterFile/n1276 ), .CK(CLK), .QN(\unit_decode/n1277 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][7]  ( .D(
        \unit_decode/RegisterFile/n1275 ), .CK(CLK), .QN(\unit_decode/n1276 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][6]  ( .D(
        \unit_decode/RegisterFile/n1274 ), .CK(CLK), .QN(\unit_decode/n1275 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][5]  ( .D(
        \unit_decode/RegisterFile/n1273 ), .CK(CLK), .QN(\unit_decode/n1274 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][4]  ( .D(
        \unit_decode/RegisterFile/n1272 ), .CK(CLK), .QN(\unit_decode/n1273 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][3]  ( .D(
        \unit_decode/RegisterFile/n1271 ), .CK(CLK), .QN(\unit_decode/n1272 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][2]  ( .D(
        \unit_decode/RegisterFile/n1270 ), .CK(CLK), .QN(\unit_decode/n1271 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][1]  ( .D(
        \unit_decode/RegisterFile/n1269 ), .CK(CLK), .QN(\unit_decode/n1270 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][0]  ( .D(
        \unit_decode/RegisterFile/n1268 ), .CK(CLK), .QN(\unit_decode/n1269 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][23]  ( .D(
        \unit_decode/RegisterFile/n1259 ), .CK(CLK), .QN(\unit_decode/n1268 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][22]  ( .D(
        \unit_decode/RegisterFile/n1258 ), .CK(CLK), .QN(\unit_decode/n1267 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][21]  ( .D(
        \unit_decode/RegisterFile/n1257 ), .CK(CLK), .QN(\unit_decode/n1266 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][20]  ( .D(
        \unit_decode/RegisterFile/n1256 ), .CK(CLK), .QN(\unit_decode/n1265 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][19]  ( .D(
        \unit_decode/RegisterFile/n1255 ), .CK(CLK), .QN(\unit_decode/n1264 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][18]  ( .D(
        \unit_decode/RegisterFile/n1254 ), .CK(CLK), .QN(\unit_decode/n1263 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][17]  ( .D(
        \unit_decode/RegisterFile/n1253 ), .CK(CLK), .QN(\unit_decode/n1262 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][16]  ( .D(
        \unit_decode/RegisterFile/n1252 ), .CK(CLK), .QN(\unit_decode/n1261 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][15]  ( .D(
        \unit_decode/RegisterFile/n1251 ), .CK(CLK), .QN(\unit_decode/n1260 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][14]  ( .D(
        \unit_decode/RegisterFile/n1250 ), .CK(CLK), .QN(\unit_decode/n1259 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][13]  ( .D(
        \unit_decode/RegisterFile/n1249 ), .CK(CLK), .QN(\unit_decode/n1258 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][12]  ( .D(
        \unit_decode/RegisterFile/n1248 ), .CK(CLK), .QN(\unit_decode/n1257 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][11]  ( .D(
        \unit_decode/RegisterFile/n1247 ), .CK(CLK), .QN(\unit_decode/n1256 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][10]  ( .D(
        \unit_decode/RegisterFile/n1246 ), .CK(CLK), .QN(\unit_decode/n1255 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][9]  ( .D(
        \unit_decode/RegisterFile/n1245 ), .CK(CLK), .QN(\unit_decode/n1254 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][8]  ( .D(
        \unit_decode/RegisterFile/n1244 ), .CK(CLK), .QN(\unit_decode/n1253 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][7]  ( .D(
        \unit_decode/RegisterFile/n1243 ), .CK(CLK), .QN(\unit_decode/n1252 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][6]  ( .D(
        \unit_decode/RegisterFile/n1242 ), .CK(CLK), .QN(\unit_decode/n1251 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][5]  ( .D(
        \unit_decode/RegisterFile/n1241 ), .CK(CLK), .QN(\unit_decode/n1250 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][4]  ( .D(
        \unit_decode/RegisterFile/n1240 ), .CK(CLK), .QN(\unit_decode/n1249 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][3]  ( .D(
        \unit_decode/RegisterFile/n1239 ), .CK(CLK), .QN(\unit_decode/n1248 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][2]  ( .D(
        \unit_decode/RegisterFile/n1238 ), .CK(CLK), .QN(\unit_decode/n1247 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][1]  ( .D(
        \unit_decode/RegisterFile/n1237 ), .CK(CLK), .QN(\unit_decode/n1246 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][0]  ( .D(
        \unit_decode/RegisterFile/n1236 ), .CK(CLK), .QN(\unit_decode/n1245 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][23]  ( .D(
        \unit_decode/RegisterFile/n1227 ), .CK(CLK), .QN(\unit_decode/n1244 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][22]  ( .D(
        \unit_decode/RegisterFile/n1226 ), .CK(CLK), .QN(\unit_decode/n1243 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][21]  ( .D(
        \unit_decode/RegisterFile/n1225 ), .CK(CLK), .QN(\unit_decode/n1242 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][20]  ( .D(
        \unit_decode/RegisterFile/n1224 ), .CK(CLK), .QN(\unit_decode/n1241 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][19]  ( .D(
        \unit_decode/RegisterFile/n1223 ), .CK(CLK), .QN(\unit_decode/n1240 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][18]  ( .D(
        \unit_decode/RegisterFile/n1222 ), .CK(CLK), .QN(\unit_decode/n1239 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][17]  ( .D(
        \unit_decode/RegisterFile/n1221 ), .CK(CLK), .QN(\unit_decode/n1238 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][16]  ( .D(
        \unit_decode/RegisterFile/n1220 ), .CK(CLK), .QN(\unit_decode/n1237 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][15]  ( .D(
        \unit_decode/RegisterFile/n1219 ), .CK(CLK), .QN(\unit_decode/n1236 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][14]  ( .D(
        \unit_decode/RegisterFile/n1218 ), .CK(CLK), .QN(\unit_decode/n1235 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][13]  ( .D(
        \unit_decode/RegisterFile/n1217 ), .CK(CLK), .QN(\unit_decode/n1234 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][12]  ( .D(
        \unit_decode/RegisterFile/n1216 ), .CK(CLK), .QN(\unit_decode/n1233 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][11]  ( .D(
        \unit_decode/RegisterFile/n1215 ), .CK(CLK), .QN(\unit_decode/n1232 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][10]  ( .D(
        \unit_decode/RegisterFile/n1214 ), .CK(CLK), .QN(\unit_decode/n1231 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][9]  ( .D(
        \unit_decode/RegisterFile/n1213 ), .CK(CLK), .QN(\unit_decode/n1230 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][8]  ( .D(
        \unit_decode/RegisterFile/n1212 ), .CK(CLK), .QN(\unit_decode/n1229 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][7]  ( .D(
        \unit_decode/RegisterFile/n1211 ), .CK(CLK), .QN(\unit_decode/n1228 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][6]  ( .D(
        \unit_decode/RegisterFile/n1210 ), .CK(CLK), .QN(\unit_decode/n1227 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][5]  ( .D(
        \unit_decode/RegisterFile/n1209 ), .CK(CLK), .QN(\unit_decode/n1226 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][4]  ( .D(
        \unit_decode/RegisterFile/n1208 ), .CK(CLK), .QN(\unit_decode/n1225 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][3]  ( .D(
        \unit_decode/RegisterFile/n1207 ), .CK(CLK), .QN(\unit_decode/n1224 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][2]  ( .D(
        \unit_decode/RegisterFile/n1206 ), .CK(CLK), .QN(\unit_decode/n1223 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][1]  ( .D(
        \unit_decode/RegisterFile/n1205 ), .CK(CLK), .QN(\unit_decode/n1222 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[29][0]  ( .D(
        \unit_decode/RegisterFile/n1204 ), .CK(CLK), .QN(\unit_decode/n1221 )
         );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][23]  ( .D(
        \unit_decode/RegisterFile/n1195 ), .CK(CLK), .Q(\unit_decode/n50 ), 
        .QN(\unit_decode/n1220 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][22]  ( .D(
        \unit_decode/RegisterFile/n1194 ), .CK(CLK), .Q(\unit_decode/n52 ), 
        .QN(\unit_decode/n1219 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][21]  ( .D(
        \unit_decode/RegisterFile/n1193 ), .CK(CLK), .Q(\unit_decode/n54 ), 
        .QN(\unit_decode/n1218 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][20]  ( .D(
        \unit_decode/RegisterFile/n1192 ), .CK(CLK), .Q(\unit_decode/n56 ), 
        .QN(\unit_decode/n1217 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][19]  ( .D(
        \unit_decode/RegisterFile/n1191 ), .CK(CLK), .Q(\unit_decode/n58 ), 
        .QN(\unit_decode/n1216 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][18]  ( .D(
        \unit_decode/RegisterFile/n1190 ), .CK(CLK), .Q(\unit_decode/n60 ), 
        .QN(\unit_decode/n1215 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][17]  ( .D(
        \unit_decode/RegisterFile/n1189 ), .CK(CLK), .Q(\unit_decode/n62 ), 
        .QN(\unit_decode/n1214 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][16]  ( .D(
        \unit_decode/RegisterFile/n1188 ), .CK(CLK), .Q(\unit_decode/n64 ), 
        .QN(\unit_decode/n1213 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][15]  ( .D(
        \unit_decode/RegisterFile/n1187 ), .CK(CLK), .Q(\unit_decode/n66 ), 
        .QN(\unit_decode/n1212 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][14]  ( .D(
        \unit_decode/RegisterFile/n1186 ), .CK(CLK), .Q(\unit_decode/n68 ), 
        .QN(\unit_decode/n1211 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][13]  ( .D(
        \unit_decode/RegisterFile/n1185 ), .CK(CLK), .Q(\unit_decode/n70 ), 
        .QN(\unit_decode/n1210 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][12]  ( .D(
        \unit_decode/RegisterFile/n1184 ), .CK(CLK), .Q(\unit_decode/n72 ), 
        .QN(\unit_decode/n1209 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][11]  ( .D(
        \unit_decode/RegisterFile/n1183 ), .CK(CLK), .Q(\unit_decode/n74 ), 
        .QN(\unit_decode/n1208 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][10]  ( .D(
        \unit_decode/RegisterFile/n1182 ), .CK(CLK), .Q(\unit_decode/n76 ), 
        .QN(\unit_decode/n1207 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][9]  ( .D(
        \unit_decode/RegisterFile/n1181 ), .CK(CLK), .Q(\unit_decode/n78 ), 
        .QN(\unit_decode/n1206 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][8]  ( .D(
        \unit_decode/RegisterFile/n1180 ), .CK(CLK), .Q(\unit_decode/n80 ), 
        .QN(\unit_decode/n1205 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][7]  ( .D(
        \unit_decode/RegisterFile/n1179 ), .CK(CLK), .Q(\unit_decode/n82 ), 
        .QN(\unit_decode/n1204 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][6]  ( .D(
        \unit_decode/RegisterFile/n1178 ), .CK(CLK), .Q(\unit_decode/n84 ), 
        .QN(\unit_decode/n1203 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][5]  ( .D(
        \unit_decode/RegisterFile/n1177 ), .CK(CLK), .Q(\unit_decode/n86 ), 
        .QN(\unit_decode/n1202 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][4]  ( .D(
        \unit_decode/RegisterFile/n1176 ), .CK(CLK), .Q(\unit_decode/n88 ), 
        .QN(\unit_decode/n1201 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][3]  ( .D(
        \unit_decode/RegisterFile/n1175 ), .CK(CLK), .Q(\unit_decode/n90 ), 
        .QN(\unit_decode/n1200 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][2]  ( .D(
        \unit_decode/RegisterFile/n1174 ), .CK(CLK), .Q(\unit_decode/n92 ), 
        .QN(\unit_decode/n1199 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][1]  ( .D(
        \unit_decode/RegisterFile/n1173 ), .CK(CLK), .Q(\unit_decode/n94 ), 
        .QN(\unit_decode/n1198 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[30][0]  ( .D(
        \unit_decode/RegisterFile/n1172 ), .CK(CLK), .Q(\unit_decode/n96 ), 
        .QN(\unit_decode/n1197 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][31]  ( .D(
        \unit_decode/RegisterFile/n1171 ), .CK(CLK), .Q(\unit_decode/n1 ), 
        .QN(\unit_decode/n1196 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][30]  ( .D(
        \unit_decode/RegisterFile/n1170 ), .CK(CLK), .Q(\unit_decode/n2 ), 
        .QN(\unit_decode/n1195 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][29]  ( .D(
        \unit_decode/RegisterFile/n1169 ), .CK(CLK), .Q(\unit_decode/n3 ), 
        .QN(\unit_decode/n1194 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][28]  ( .D(
        \unit_decode/RegisterFile/n1168 ), .CK(CLK), .Q(\unit_decode/n4 ), 
        .QN(\unit_decode/n1193 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][27]  ( .D(
        \unit_decode/RegisterFile/n1167 ), .CK(CLK), .Q(\unit_decode/n5 ), 
        .QN(\unit_decode/n1192 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][26]  ( .D(
        \unit_decode/RegisterFile/n1166 ), .CK(CLK), .Q(\unit_decode/n6 ), 
        .QN(\unit_decode/n1191 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][25]  ( .D(
        \unit_decode/RegisterFile/n1165 ), .CK(CLK), .Q(\unit_decode/n7 ), 
        .QN(\unit_decode/n1190 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][24]  ( .D(
        \unit_decode/RegisterFile/n1164 ), .CK(CLK), .Q(\unit_decode/n8 ), 
        .QN(\unit_decode/n1189 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][23]  ( .D(
        \unit_decode/RegisterFile/n1163 ), .CK(CLK), .Q(\unit_decode/n9 ), 
        .QN(\unit_decode/n1188 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][22]  ( .D(
        \unit_decode/RegisterFile/n1162 ), .CK(CLK), .Q(\unit_decode/n10 ), 
        .QN(\unit_decode/n1187 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][21]  ( .D(
        \unit_decode/RegisterFile/n1161 ), .CK(CLK), .Q(\unit_decode/n11 ), 
        .QN(\unit_decode/n1186 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][20]  ( .D(
        \unit_decode/RegisterFile/n1160 ), .CK(CLK), .Q(\unit_decode/n12 ), 
        .QN(\unit_decode/n1185 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][19]  ( .D(
        \unit_decode/RegisterFile/n1159 ), .CK(CLK), .Q(\unit_decode/n13 ), 
        .QN(\unit_decode/n1184 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][18]  ( .D(
        \unit_decode/RegisterFile/n1158 ), .CK(CLK), .Q(\unit_decode/n14 ), 
        .QN(\unit_decode/n1183 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][17]  ( .D(
        \unit_decode/RegisterFile/n1157 ), .CK(CLK), .Q(\unit_decode/n15 ), 
        .QN(\unit_decode/n1182 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][16]  ( .D(
        \unit_decode/RegisterFile/n1156 ), .CK(CLK), .Q(\unit_decode/n16 ), 
        .QN(\unit_decode/n1181 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][15]  ( .D(
        \unit_decode/RegisterFile/n1155 ), .CK(CLK), .Q(\unit_decode/n17 ), 
        .QN(\unit_decode/n1180 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][14]  ( .D(
        \unit_decode/RegisterFile/n1154 ), .CK(CLK), .Q(\unit_decode/n18 ), 
        .QN(\unit_decode/n1179 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][13]  ( .D(
        \unit_decode/RegisterFile/n1153 ), .CK(CLK), .Q(\unit_decode/n19 ), 
        .QN(\unit_decode/n1178 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][12]  ( .D(
        \unit_decode/RegisterFile/n1152 ), .CK(CLK), .Q(\unit_decode/n20 ), 
        .QN(\unit_decode/n1177 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][11]  ( .D(
        \unit_decode/RegisterFile/n1151 ), .CK(CLK), .Q(\unit_decode/n21 ), 
        .QN(\unit_decode/n1176 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][10]  ( .D(
        \unit_decode/RegisterFile/n1150 ), .CK(CLK), .Q(\unit_decode/n22 ), 
        .QN(\unit_decode/n1175 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][9]  ( .D(
        \unit_decode/RegisterFile/n1149 ), .CK(CLK), .Q(\unit_decode/n23 ), 
        .QN(\unit_decode/n1174 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[31][8]  ( .D(
        \unit_decode/RegisterFile/n1148 ), .CK(CLK), .Q(\unit_decode/n24 ), 
        .QN(\unit_decode/n1173 ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[31]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N410 ), .Q(\unit_decode/registerA[31] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[30]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N409 ), .Q(\unit_decode/registerA[30] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[29]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N408 ), .Q(\unit_decode/registerA[29] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[28]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N407 ), .Q(\unit_decode/registerA[28] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[27]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N406 ), .Q(\unit_decode/registerA[27] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[26]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N405 ), .Q(\unit_decode/registerA[26] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[25]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N404 ), .Q(\unit_decode/registerA[25] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[24]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N403 ), .Q(\unit_decode/registerA[24] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[23]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N402 ), .Q(\unit_decode/registerA[23] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[22]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N401 ), .Q(\unit_decode/registerA[22] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[21]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N400 ), .Q(\unit_decode/registerA[21] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[20]  ( .G(n708), .D(
        \unit_decode/RegisterFile/N399 ), .Q(\unit_decode/registerA[20] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[19]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N398 ), .Q(\unit_decode/registerA[19] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[18]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N397 ), .Q(\unit_decode/registerA[18] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[17]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N396 ), .Q(\unit_decode/registerA[17] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[16]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N395 ), .Q(\unit_decode/registerA[16] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[15]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N394 ), .Q(\unit_decode/registerA[15] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[14]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N393 ), .Q(\unit_decode/registerA[14] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[13]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N392 ), .Q(\unit_decode/registerA[13] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[12]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N391 ), .Q(\unit_decode/registerA[12] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[11]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N390 ), .Q(\unit_decode/registerA[11] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[10]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N389 ), .Q(\unit_decode/registerA[10] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[9]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N388 ), .Q(\unit_decode/registerA[9] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[8]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N387 ), .Q(\unit_decode/registerA[8] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[7]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N386 ), .Q(\unit_decode/registerA[7] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[6]  ( .G(n707), .D(
        \unit_decode/RegisterFile/N385 ), .Q(\unit_decode/registerA[6] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[5]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N384 ), .Q(\unit_decode/registerA[5] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[4]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N383 ), .Q(\unit_decode/registerA[4] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[3]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N382 ), .Q(\unit_decode/registerA[3] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[2]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N381 ), .Q(\unit_decode/registerA[2] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[1]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N380 ), .Q(\unit_decode/registerA[1] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT1_reg[0]  ( .G(n706), .D(
        \unit_decode/RegisterFile/N379 ), .Q(\unit_decode/registerA[0] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[31]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N443 ), .Q(\unit_decode/registerB[31] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[30]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N442 ), .Q(\unit_decode/registerB[30] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[29]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N441 ), .Q(\unit_decode/registerB[29] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[28]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N440 ), .Q(\unit_decode/registerB[28] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[27]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N439 ), .Q(\unit_decode/registerB[27] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[26]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N438 ), .Q(\unit_decode/registerB[26] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[25]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N437 ), .Q(\unit_decode/registerB[25] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[24]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N436 ), .Q(\unit_decode/registerB[24] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[23]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N435 ), .Q(\unit_decode/registerB[23] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[22]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N434 ), .Q(\unit_decode/registerB[22] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[21]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N433 ), .Q(\unit_decode/registerB[21] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[20]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N432 ), .Q(\unit_decode/registerB[20] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[19]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N431 ), .Q(\unit_decode/registerB[19] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[18]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N430 ), .Q(\unit_decode/registerB[18] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[17]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N429 ), .Q(\unit_decode/registerB[17] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[16]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N428 ), .Q(\unit_decode/registerB[16] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[15]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N427 ), .Q(\unit_decode/registerB[15] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[14]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N426 ), .Q(\unit_decode/registerB[14] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[13]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N425 ), .Q(\unit_decode/registerB[13] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[12]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N424 ), .Q(\unit_decode/registerB[12] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[11]  ( .G(n705), .D(
        \unit_decode/RegisterFile/N423 ), .Q(\unit_decode/registerB[11] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[10]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N422 ), .Q(\unit_decode/registerB[10] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[9]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N421 ), .Q(\unit_decode/registerB[9] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[8]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N420 ), .Q(\unit_decode/registerB[8] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[7]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N419 ), .Q(\unit_decode/registerB[7] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[6]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N418 ), .Q(\unit_decode/registerB[6] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[5]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N417 ), .Q(\unit_decode/registerB[5] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[4]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N416 ), .Q(\unit_decode/registerB[4] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[3]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N415 ), .Q(\unit_decode/registerB[3] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[2]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N414 ), .Q(\unit_decode/registerB[2] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[1]  ( .G(n704), .D(
        \unit_decode/RegisterFile/N413 ), .Q(\unit_decode/registerB[1] ) );
  DLH_X1 \unit_decode/RegisterFile/OUT2_reg[0]  ( .G(n703), .D(
        \unit_decode/RegisterFile/N412 ), .Q(\unit_decode/registerB[0] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[0]  ( .G(1'b0), .D(\unit_memory/DRAM/N566 ), .Q(\unit_memory/DataMemOut[0] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[1]  ( .G(1'b0), .D(\unit_memory/DRAM/N567 ), .Q(\unit_memory/DataMemOut[1] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[2]  ( .G(1'b0), .D(\unit_memory/DRAM/N568 ), .Q(\unit_memory/DataMemOut[2] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[3]  ( .G(1'b0), .D(\unit_memory/DRAM/N569 ), .Q(\unit_memory/DataMemOut[3] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[4]  ( .G(1'b0), .D(\unit_memory/DRAM/N570 ), .Q(\unit_memory/DataMemOut[4] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[5]  ( .G(1'b0), .D(\unit_memory/DRAM/N571 ), .Q(\unit_memory/DataMemOut[5] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[6]  ( .G(1'b0), .D(\unit_memory/DRAM/N572 ), .Q(\unit_memory/DataMemOut[6] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[7]  ( .G(1'b0), .D(\unit_memory/DRAM/N573 ), .Q(\unit_memory/DataMemOut[7] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[8]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3398 ), .Q(\unit_memory/DataMemOut[8] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[9]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3397 ), .Q(\unit_memory/DataMemOut[9] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[10]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3396 ), .Q(\unit_memory/DataMemOut[10] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[11]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3395 ), .Q(\unit_memory/DataMemOut[11] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[12]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3394 ), .Q(\unit_memory/DataMemOut[12] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[13]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3393 ), .Q(\unit_memory/DataMemOut[13] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[14]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3392 ), .Q(\unit_memory/DataMemOut[14] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[15]  ( .G(1'b0), .D(
        \unit_memory/DRAM/n3391 ), .Q(\unit_memory/DataMemOut[15] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[16]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N582 ), .Q(\unit_memory/DataMemOut[16] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[17]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N583 ), .Q(\unit_memory/DataMemOut[17] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[18]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N584 ), .Q(\unit_memory/DataMemOut[18] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[19]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N585 ), .Q(\unit_memory/DataMemOut[19] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[20]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N586 ), .Q(\unit_memory/DataMemOut[20] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[21]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N587 ), .Q(\unit_memory/DataMemOut[21] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[22]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N588 ), .Q(\unit_memory/DataMemOut[22] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[23]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N589 ), .Q(\unit_memory/DataMemOut[23] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[24]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N590 ), .Q(\unit_memory/DataMemOut[24] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[25]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N591 ), .Q(\unit_memory/DataMemOut[25] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[26]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N592 ), .Q(\unit_memory/DataMemOut[26] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[27]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N593 ), .Q(\unit_memory/DataMemOut[27] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[28]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N594 ), .Q(\unit_memory/DataMemOut[28] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[29]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N595 ), .Q(\unit_memory/DataMemOut[29] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[30]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N596 ), .Q(\unit_memory/DataMemOut[30] ) );
  DLH_X1 \unit_memory/DRAM/Dout_reg[31]  ( .G(1'b0), .D(
        \unit_memory/DRAM/N597 ), .Q(\unit_memory/DataMemOut[31] ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_12/n5 ), .CK(CLK), .Q(cw_ex[3]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_11/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_11/n5 ), .CK(CLK), .Q(cw_ex[2]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_10/n5 ), .CK(CLK), .Q(cw_ex[1]) );
  DFF_X1 \unit_decode/IMMreg/ffi_7/Q_reg  ( .D(\unit_decode/IMMreg/ffi_7/n5 ), 
        .CK(CLK), .Q(imm_out[7]), .QN(\unit_decode/n209 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_15/Q_reg  ( .D(\unit_decode/IMMreg/ffi_15/n5 ), .CK(CLK), .Q(imm_out[15]), .QN(\unit_decode/n3614 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_14/Q_reg  ( .D(\unit_decode/IMMreg/ffi_14/n5 ), .CK(CLK), .Q(imm_out[14]), .QN(\unit_decode/n3615 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_11/Q_reg  ( .D(\unit_decode/IMMreg/ffi_11/n5 ), .CK(CLK), .Q(imm_out[11]), .QN(\unit_decode/n3618 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_6/Q_reg  ( .D(\unit_decode/IMMreg/ffi_6/n5 ), 
        .CK(CLK), .Q(imm_out[6]), .QN(\unit_decode/n197 ) );
  DFF_X1 \unit_decode/Areg/ffi_11/Q_reg  ( .D(\unit_decode/Areg/ffi_11/n5 ), 
        .CK(CLK), .Q(rega_out[11]), .QN(\unit_decode/n3530 ) );
  DFF_X1 \unit_decode/Areg/ffi_10/Q_reg  ( .D(\unit_decode/Areg/ffi_10/n5 ), 
        .CK(CLK), .Q(rega_out[10]), .QN(\unit_decode/n3531 ) );
  DFF_X1 \unit_decode/Breg/ffi_19/Q_reg  ( .D(\unit_decode/Breg/ffi_19/n5 ), 
        .CK(CLK), .Q(regb_out[19]), .QN(\unit_decode/n3550 ) );
  DFF_X1 \unit_decode/Breg/ffi_18/Q_reg  ( .D(\unit_decode/Breg/ffi_18/n5 ), 
        .CK(CLK), .Q(regb_out[18]), .QN(\unit_decode/n3551 ) );
  DFF_X1 \unit_decode/Breg/ffi_17/Q_reg  ( .D(\unit_decode/Breg/ffi_17/n5 ), 
        .CK(CLK), .Q(regb_out[17]), .QN(\unit_decode/n3552 ) );
  DFF_X1 \unit_decode/Breg/ffi_16/Q_reg  ( .D(\unit_decode/Breg/ffi_16/n5 ), 
        .CK(CLK), .Q(regb_out[16]), .QN(\unit_decode/n3553 ) );
  DFF_X1 \unit_decode/Breg/ffi_15/Q_reg  ( .D(\unit_decode/Breg/ffi_15/n5 ), 
        .CK(CLK), .Q(regb_out[15]), .QN(\unit_decode/n3554 ) );
  DFF_X1 \unit_decode/Breg/ffi_14/Q_reg  ( .D(\unit_decode/Breg/ffi_14/n5 ), 
        .CK(CLK), .Q(regb_out[14]), .QN(\unit_decode/n3555 ) );
  DFF_X1 \unit_decode/Breg/ffi_13/Q_reg  ( .D(\unit_decode/Breg/ffi_13/n5 ), 
        .CK(CLK), .Q(regb_out[13]), .QN(\unit_decode/n3556 ) );
  DFF_X1 \unit_decode/Breg/ffi_12/Q_reg  ( .D(\unit_decode/Breg/ffi_12/n5 ), 
        .CK(CLK), .Q(regb_out[12]), .QN(\unit_decode/n3557 ) );
  DFF_X1 \unit_decode/Breg/ffi_11/Q_reg  ( .D(\unit_decode/Breg/ffi_11/n5 ), 
        .CK(CLK), .Q(regb_out[11]), .QN(\unit_decode/n3558 ) );
  DFF_X1 \unit_decode/Breg/ffi_10/Q_reg  ( .D(\unit_decode/Breg/ffi_10/n5 ), 
        .CK(CLK), .Q(regb_out[10]), .QN(\unit_decode/n3622 ) );
  DFF_X1 \unit_decode/Breg/ffi_1/Q_reg  ( .D(\unit_decode/Breg/ffi_1/n5 ), 
        .CK(CLK), .Q(regb_out[1]), .QN(\unit_decode/n233 ) );
  DFF_X1 \unit_decode/Breg/ffi_0/Q_reg  ( .D(\unit_decode/Breg/ffi_0/n5 ), 
        .CK(CLK), .Q(regb_out[0]), .QN(\unit_decode/n239 ) );
  DFF_X1 \unit_decode/Areg/ffi_31/Q_reg  ( .D(\unit_decode/Areg/ffi_31/n5 ), 
        .CK(CLK), .Q(rega_out[31]), .QN(\unit_decode/n3587 ) );
  DFF_X1 \unit_decode/Areg/ffi_30/Q_reg  ( .D(\unit_decode/Areg/ffi_30/n5 ), 
        .CK(CLK), .Q(rega_out[30]), .QN(\unit_decode/n3588 ) );
  DFF_X1 \unit_decode/Areg/ffi_29/Q_reg  ( .D(\unit_decode/Areg/ffi_29/n5 ), 
        .CK(CLK), .Q(rega_out[29]), .QN(\unit_decode/n3589 ) );
  DFF_X1 \unit_decode/Areg/ffi_28/Q_reg  ( .D(\unit_decode/Areg/ffi_28/n5 ), 
        .CK(CLK), .Q(rega_out[28]), .QN(\unit_decode/n3590 ) );
  DFF_X1 \unit_decode/Areg/ffi_27/Q_reg  ( .D(\unit_decode/Areg/ffi_27/n5 ), 
        .CK(CLK), .Q(rega_out[27]), .QN(\unit_decode/n3591 ) );
  DFF_X1 \unit_decode/Areg/ffi_26/Q_reg  ( .D(\unit_decode/Areg/ffi_26/n5 ), 
        .CK(CLK), .Q(rega_out[26]), .QN(\unit_decode/n3592 ) );
  DFF_X1 \unit_decode/Areg/ffi_25/Q_reg  ( .D(\unit_decode/Areg/ffi_25/n5 ), 
        .CK(CLK), .Q(rega_out[25]), .QN(\unit_decode/n3593 ) );
  DFF_X1 \unit_decode/Areg/ffi_24/Q_reg  ( .D(\unit_decode/Areg/ffi_24/n5 ), 
        .CK(CLK), .Q(rega_out[24]), .QN(\unit_decode/n3594 ) );
  DFF_X1 \unit_decode/Areg/ffi_23/Q_reg  ( .D(\unit_decode/Areg/ffi_23/n5 ), 
        .CK(CLK), .Q(rega_out[23]), .QN(\unit_decode/n3595 ) );
  DFF_X1 \unit_decode/Areg/ffi_22/Q_reg  ( .D(\unit_decode/Areg/ffi_22/n5 ), 
        .CK(CLK), .Q(rega_out[22]), .QN(\unit_decode/n3596 ) );
  DFF_X1 \unit_decode/Areg/ffi_21/Q_reg  ( .D(\unit_decode/Areg/ffi_21/n5 ), 
        .CK(CLK), .Q(rega_out[21]), .QN(\unit_decode/n3597 ) );
  DFF_X1 \unit_decode/Areg/ffi_20/Q_reg  ( .D(\unit_decode/Areg/ffi_20/n5 ), 
        .CK(CLK), .Q(rega_out[20]), .QN(\unit_decode/n3598 ) );
  DFF_X1 \unit_decode/Areg/ffi_19/Q_reg  ( .D(\unit_decode/Areg/ffi_19/n5 ), 
        .CK(CLK), .Q(rega_out[19]), .QN(\unit_decode/n3599 ) );
  DFF_X1 \unit_decode/Areg/ffi_18/Q_reg  ( .D(\unit_decode/Areg/ffi_18/n5 ), 
        .CK(CLK), .Q(rega_out[18]), .QN(\unit_decode/n3523 ) );
  DFF_X1 \unit_decode/Areg/ffi_17/Q_reg  ( .D(\unit_decode/Areg/ffi_17/n5 ), 
        .CK(CLK), .Q(rega_out[17]), .QN(\unit_decode/n3524 ) );
  DFF_X1 \unit_decode/Areg/ffi_16/Q_reg  ( .D(\unit_decode/Areg/ffi_16/n5 ), 
        .CK(CLK), .Q(rega_out[16]), .QN(\unit_decode/n3525 ) );
  DFF_X1 \unit_decode/Areg/ffi_15/Q_reg  ( .D(\unit_decode/Areg/ffi_15/n5 ), 
        .CK(CLK), .Q(rega_out[15]), .QN(\unit_decode/n3526 ) );
  DFF_X1 \unit_decode/Areg/ffi_14/Q_reg  ( .D(\unit_decode/Areg/ffi_14/n5 ), 
        .CK(CLK), .Q(rega_out[14]), .QN(\unit_decode/n3527 ) );
  DFF_X1 \unit_decode/Areg/ffi_6/Q_reg  ( .D(\unit_decode/Areg/ffi_6/n5 ), 
        .CK(CLK), .Q(rega_out[6]), .QN(\unit_decode/n3535 ) );
  DFF_X1 \unit_decode/Breg/ffi_31/Q_reg  ( .D(\unit_decode/Breg/ffi_31/n5 ), 
        .CK(CLK), .Q(regb_out[31]), .QN(\unit_decode/n3538 ) );
  DFF_X1 \unit_decode/Breg/ffi_9/Q_reg  ( .D(\unit_decode/Breg/ffi_9/n5 ), 
        .CK(CLK), .Q(regb_out[9]), .QN(\unit_decode/n3623 ) );
  DFF_X1 \unit_decode/Breg/ffi_8/Q_reg  ( .D(\unit_decode/Breg/ffi_8/n5 ), 
        .CK(CLK), .Q(regb_out[8]), .QN(\unit_decode/n3624 ) );
  DFF_X1 \unit_decode/Breg/ffi_7/Q_reg  ( .D(\unit_decode/Breg/ffi_7/n5 ), 
        .CK(CLK), .Q(regb_out[7]), .QN(\unit_decode/n219 ) );
  DFF_X1 \unit_decode/Breg/ffi_6/Q_reg  ( .D(\unit_decode/Breg/ffi_6/n5 ), 
        .CK(CLK), .Q(regb_out[6]), .QN(\unit_decode/n207 ) );
  DFF_X1 \unit_decode/Breg/ffi_5/Q_reg  ( .D(\unit_decode/Breg/ffi_5/n5 ), 
        .CK(CLK), .Q(regb_out[5]), .QN(\unit_decode/n223 ) );
  DFF_X1 \unit_decode/Breg/ffi_4/Q_reg  ( .D(\unit_decode/Breg/ffi_4/n5 ), 
        .CK(CLK), .Q(regb_out[4]), .QN(\unit_decode/n221 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_4/Q_reg  ( .D(\unit_decode/RD1reg/ffi_4/n5 ), 
        .CK(CLK), .Q(rd1_out[4]), .QN(n1397) );
  DFF_X1 \unit_decode/RD1reg/ffi_3/Q_reg  ( .D(\unit_decode/RD1reg/ffi_3/n5 ), 
        .CK(CLK), .Q(rd1_out[3]), .QN(n1386) );
  DFF_X1 \unit_decode/RD1reg/ffi_2/Q_reg  ( .D(\unit_decode/RD1reg/ffi_2/n5 ), 
        .CK(CLK), .Q(rd1_out[2]), .QN(n1375) );
  DFF_X1 \unit_decode/RD1reg/ffi_1/Q_reg  ( .D(\unit_decode/RD1reg/ffi_1/n5 ), 
        .CK(CLK), .Q(rd1_out[1]), .QN(n1396) );
  DFF_X1 \unit_decode/RD1reg/ffi_0/Q_reg  ( .D(\unit_decode/RD1reg/ffi_0/n5 ), 
        .CK(CLK), .Q(rd1_out[0]), .QN(n1374) );
  DFF_X1 \unit_decode/NPC1reg/ffi_31/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_31/n5 ), .CK(CLK), .Q(npc1_out[31]), .QN(
        \unit_decode/n3626 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_30/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_30/n5 ), .CK(CLK), .Q(npc1_out[30]), .QN(
        \unit_decode/n3560 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_29/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_29/n5 ), .CK(CLK), .Q(npc1_out[29]), .QN(
        \unit_decode/n3561 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_28/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_28/n5 ), .CK(CLK), .Q(npc1_out[28]), .QN(
        \unit_decode/n3562 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_27/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_27/n5 ), .CK(CLK), .Q(npc1_out[27]), .QN(
        \unit_decode/n3563 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_26/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_26/n5 ), .CK(CLK), .Q(npc1_out[26]), .QN(
        \unit_decode/n3564 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_25/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_25/n5 ), .CK(CLK), .Q(npc1_out[25]), .QN(
        \unit_decode/n3565 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_24/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_24/n5 ), .CK(CLK), .Q(npc1_out[24]), .QN(
        \unit_decode/n3566 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_23/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_23/n5 ), .CK(CLK), .Q(npc1_out[23]), .QN(
        \unit_decode/n3567 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_22/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_22/n5 ), .CK(CLK), .Q(npc1_out[22]), .QN(
        \unit_decode/n3568 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_21/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_21/n5 ), .CK(CLK), .Q(npc1_out[21]), .QN(
        \unit_decode/n3569 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_20/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_20/n5 ), .CK(CLK), .Q(npc1_out[20]), .QN(
        \unit_decode/n3570 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_19/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_19/n5 ), .CK(CLK), .Q(npc1_out[19]), .QN(
        \unit_decode/n3571 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_18/Q_reg  ( .D(
        \unit_decode/NPC1reg/ffi_18/n5 ), .CK(CLK), .Q(npc1_out[18]), .QN(
        \unit_decode/n3572 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][31]  ( .D(
        \unit_decode/RegisterFile/n1427 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3708 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][30]  ( .D(
        \unit_decode/RegisterFile/n1426 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3709 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][29]  ( .D(
        \unit_decode/RegisterFile/n1425 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3710 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][28]  ( .D(
        \unit_decode/RegisterFile/n1424 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3711 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][27]  ( .D(
        \unit_decode/RegisterFile/n1423 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3712 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][26]  ( .D(
        \unit_decode/RegisterFile/n1422 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3713 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][25]  ( .D(
        \unit_decode/RegisterFile/n1421 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3714 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][24]  ( .D(
        \unit_decode/RegisterFile/n1420 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3715 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][31]  ( .D(
        \unit_decode/RegisterFile/n1459 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3676 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][30]  ( .D(
        \unit_decode/RegisterFile/n1458 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3677 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][29]  ( .D(
        \unit_decode/RegisterFile/n1457 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3678 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][28]  ( .D(
        \unit_decode/RegisterFile/n1456 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3679 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][27]  ( .D(
        \unit_decode/RegisterFile/n1455 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3680 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][26]  ( .D(
        \unit_decode/RegisterFile/n1454 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3681 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][25]  ( .D(
        \unit_decode/RegisterFile/n1453 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3682 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][24]  ( .D(
        \unit_decode/RegisterFile/n1452 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3683 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][31]  ( .D(
        \unit_decode/RegisterFile/n1491 ), .CK(CLK), .Q(\unit_decode/n1748 ), 
        .QN(\unit_decode/RegisterFile/n3644 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][30]  ( .D(
        \unit_decode/RegisterFile/n1490 ), .CK(CLK), .Q(\unit_decode/n1749 ), 
        .QN(\unit_decode/RegisterFile/n3645 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][29]  ( .D(
        \unit_decode/RegisterFile/n1489 ), .CK(CLK), .Q(\unit_decode/n1750 ), 
        .QN(\unit_decode/RegisterFile/n3646 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][28]  ( .D(
        \unit_decode/RegisterFile/n1488 ), .CK(CLK), .Q(\unit_decode/n1751 ), 
        .QN(\unit_decode/RegisterFile/n3647 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][27]  ( .D(
        \unit_decode/RegisterFile/n1487 ), .CK(CLK), .Q(\unit_decode/n1752 ), 
        .QN(\unit_decode/RegisterFile/n3648 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][26]  ( .D(
        \unit_decode/RegisterFile/n1486 ), .CK(CLK), .Q(\unit_decode/n1753 ), 
        .QN(\unit_decode/RegisterFile/n3649 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][25]  ( .D(
        \unit_decode/RegisterFile/n1485 ), .CK(CLK), .Q(\unit_decode/n1754 ), 
        .QN(\unit_decode/RegisterFile/n3650 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][24]  ( .D(
        \unit_decode/RegisterFile/n1484 ), .CK(CLK), .Q(\unit_decode/n1755 ), 
        .QN(\unit_decode/RegisterFile/n3651 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][31]  ( .D(
        \unit_decode/RegisterFile/n1523 ), .CK(CLK), .Q(\unit_decode/n1756 ), 
        .QN(\unit_decode/RegisterFile/n3612 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][30]  ( .D(
        \unit_decode/RegisterFile/n1522 ), .CK(CLK), .Q(\unit_decode/n1757 ), 
        .QN(\unit_decode/RegisterFile/n3613 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][29]  ( .D(
        \unit_decode/RegisterFile/n1521 ), .CK(CLK), .Q(\unit_decode/n1758 ), 
        .QN(\unit_decode/RegisterFile/n3614 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][28]  ( .D(
        \unit_decode/RegisterFile/n1520 ), .CK(CLK), .Q(\unit_decode/n1759 ), 
        .QN(\unit_decode/RegisterFile/n3615 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][27]  ( .D(
        \unit_decode/RegisterFile/n1519 ), .CK(CLK), .Q(\unit_decode/n1760 ), 
        .QN(\unit_decode/RegisterFile/n3616 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][26]  ( .D(
        \unit_decode/RegisterFile/n1518 ), .CK(CLK), .Q(\unit_decode/n1761 ), 
        .QN(\unit_decode/RegisterFile/n3617 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][25]  ( .D(
        \unit_decode/RegisterFile/n1517 ), .CK(CLK), .Q(\unit_decode/n1762 ), 
        .QN(\unit_decode/RegisterFile/n3618 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][24]  ( .D(
        \unit_decode/RegisterFile/n1516 ), .CK(CLK), .Q(\unit_decode/n1763 ), 
        .QN(\unit_decode/RegisterFile/n3619 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][28]  ( .D(
        \unit_decode/RegisterFile/n1552 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3583 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][27]  ( .D(
        \unit_decode/RegisterFile/n1551 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3584 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][26]  ( .D(
        \unit_decode/RegisterFile/n1550 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3585 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][25]  ( .D(
        \unit_decode/RegisterFile/n1549 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3586 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][24]  ( .D(
        \unit_decode/RegisterFile/n1548 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3587 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][3]  ( .D(
        \unit_decode/RegisterFile/n1623 ), .CK(CLK), .Q(\unit_decode/n2080 ), 
        .QN(\unit_decode/RegisterFile/n3512 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][2]  ( .D(
        \unit_decode/RegisterFile/n1622 ), .CK(CLK), .Q(\unit_decode/n2081 ), 
        .QN(\unit_decode/RegisterFile/n3513 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][23]  ( .D(
        \unit_decode/RegisterFile/n1419 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3716 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][22]  ( .D(
        \unit_decode/RegisterFile/n1418 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3717 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][21]  ( .D(
        \unit_decode/RegisterFile/n1417 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3718 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][20]  ( .D(
        \unit_decode/RegisterFile/n1416 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3719 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][19]  ( .D(
        \unit_decode/RegisterFile/n1415 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3720 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][18]  ( .D(
        \unit_decode/RegisterFile/n1414 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3721 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][17]  ( .D(
        \unit_decode/RegisterFile/n1413 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3722 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][16]  ( .D(
        \unit_decode/RegisterFile/n1412 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3723 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][15]  ( .D(
        \unit_decode/RegisterFile/n1411 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3724 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][14]  ( .D(
        \unit_decode/RegisterFile/n1410 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3725 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][13]  ( .D(
        \unit_decode/RegisterFile/n1409 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3726 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][12]  ( .D(
        \unit_decode/RegisterFile/n1408 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3727 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][11]  ( .D(
        \unit_decode/RegisterFile/n1407 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3728 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][10]  ( .D(
        \unit_decode/RegisterFile/n1406 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3729 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][9]  ( .D(
        \unit_decode/RegisterFile/n1405 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3730 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][8]  ( .D(
        \unit_decode/RegisterFile/n1404 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3731 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][7]  ( .D(
        \unit_decode/RegisterFile/n1403 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3732 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][6]  ( .D(
        \unit_decode/RegisterFile/n1402 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3733 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][5]  ( .D(
        \unit_decode/RegisterFile/n1401 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3734 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][4]  ( .D(
        \unit_decode/RegisterFile/n1400 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3735 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][3]  ( .D(
        \unit_decode/RegisterFile/n1399 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3736 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][2]  ( .D(
        \unit_decode/RegisterFile/n1398 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3737 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][1]  ( .D(
        \unit_decode/RegisterFile/n1397 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3738 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[23][0]  ( .D(
        \unit_decode/RegisterFile/n1396 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3739 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][23]  ( .D(
        \unit_decode/RegisterFile/n1451 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3684 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][22]  ( .D(
        \unit_decode/RegisterFile/n1450 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3685 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][21]  ( .D(
        \unit_decode/RegisterFile/n1449 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3686 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][20]  ( .D(
        \unit_decode/RegisterFile/n1448 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3687 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][19]  ( .D(
        \unit_decode/RegisterFile/n1447 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3688 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][18]  ( .D(
        \unit_decode/RegisterFile/n1446 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3689 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][17]  ( .D(
        \unit_decode/RegisterFile/n1445 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3690 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][16]  ( .D(
        \unit_decode/RegisterFile/n1444 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3691 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][15]  ( .D(
        \unit_decode/RegisterFile/n1443 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3692 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][14]  ( .D(
        \unit_decode/RegisterFile/n1442 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3693 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][13]  ( .D(
        \unit_decode/RegisterFile/n1441 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3694 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][12]  ( .D(
        \unit_decode/RegisterFile/n1440 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3695 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][11]  ( .D(
        \unit_decode/RegisterFile/n1439 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3696 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][10]  ( .D(
        \unit_decode/RegisterFile/n1438 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3697 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][9]  ( .D(
        \unit_decode/RegisterFile/n1437 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3698 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][8]  ( .D(
        \unit_decode/RegisterFile/n1436 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3699 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][7]  ( .D(
        \unit_decode/RegisterFile/n1435 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3700 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][6]  ( .D(
        \unit_decode/RegisterFile/n1434 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3701 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][5]  ( .D(
        \unit_decode/RegisterFile/n1433 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3702 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][4]  ( .D(
        \unit_decode/RegisterFile/n1432 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3703 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][3]  ( .D(
        \unit_decode/RegisterFile/n1431 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3704 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][2]  ( .D(
        \unit_decode/RegisterFile/n1430 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3705 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][1]  ( .D(
        \unit_decode/RegisterFile/n1429 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3706 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[22][0]  ( .D(
        \unit_decode/RegisterFile/n1428 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3707 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][23]  ( .D(
        \unit_decode/RegisterFile/n1483 ), .CK(CLK), .Q(\unit_decode/n1964 ), 
        .QN(\unit_decode/RegisterFile/n3652 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][22]  ( .D(
        \unit_decode/RegisterFile/n1482 ), .CK(CLK), .Q(\unit_decode/n1965 ), 
        .QN(\unit_decode/RegisterFile/n3653 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][21]  ( .D(
        \unit_decode/RegisterFile/n1481 ), .CK(CLK), .Q(\unit_decode/n1966 ), 
        .QN(\unit_decode/RegisterFile/n3654 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][20]  ( .D(
        \unit_decode/RegisterFile/n1480 ), .CK(CLK), .Q(\unit_decode/n1967 ), 
        .QN(\unit_decode/RegisterFile/n3655 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][19]  ( .D(
        \unit_decode/RegisterFile/n1479 ), .CK(CLK), .Q(\unit_decode/n1968 ), 
        .QN(\unit_decode/RegisterFile/n3656 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][18]  ( .D(
        \unit_decode/RegisterFile/n1478 ), .CK(CLK), .Q(\unit_decode/n1969 ), 
        .QN(\unit_decode/RegisterFile/n3657 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][17]  ( .D(
        \unit_decode/RegisterFile/n1477 ), .CK(CLK), .Q(\unit_decode/n1970 ), 
        .QN(\unit_decode/RegisterFile/n3658 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][16]  ( .D(
        \unit_decode/RegisterFile/n1476 ), .CK(CLK), .Q(\unit_decode/n1971 ), 
        .QN(\unit_decode/RegisterFile/n3659 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][15]  ( .D(
        \unit_decode/RegisterFile/n1475 ), .CK(CLK), .Q(\unit_decode/n1972 ), 
        .QN(\unit_decode/RegisterFile/n3660 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][14]  ( .D(
        \unit_decode/RegisterFile/n1474 ), .CK(CLK), .Q(\unit_decode/n1973 ), 
        .QN(\unit_decode/RegisterFile/n3661 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][13]  ( .D(
        \unit_decode/RegisterFile/n1473 ), .CK(CLK), .Q(\unit_decode/n1974 ), 
        .QN(\unit_decode/RegisterFile/n3662 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][12]  ( .D(
        \unit_decode/RegisterFile/n1472 ), .CK(CLK), .Q(\unit_decode/n1975 ), 
        .QN(\unit_decode/RegisterFile/n3663 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][11]  ( .D(
        \unit_decode/RegisterFile/n1471 ), .CK(CLK), .Q(\unit_decode/n1976 ), 
        .QN(\unit_decode/RegisterFile/n3664 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][10]  ( .D(
        \unit_decode/RegisterFile/n1470 ), .CK(CLK), .Q(\unit_decode/n1977 ), 
        .QN(\unit_decode/RegisterFile/n3665 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][9]  ( .D(
        \unit_decode/RegisterFile/n1469 ), .CK(CLK), .Q(\unit_decode/n1978 ), 
        .QN(\unit_decode/RegisterFile/n3666 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][8]  ( .D(
        \unit_decode/RegisterFile/n1468 ), .CK(CLK), .Q(\unit_decode/n1979 ), 
        .QN(\unit_decode/RegisterFile/n3667 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][7]  ( .D(
        \unit_decode/RegisterFile/n1467 ), .CK(CLK), .Q(\unit_decode/n1980 ), 
        .QN(\unit_decode/RegisterFile/n3668 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][6]  ( .D(
        \unit_decode/RegisterFile/n1466 ), .CK(CLK), .Q(\unit_decode/n1981 ), 
        .QN(\unit_decode/RegisterFile/n3669 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][5]  ( .D(
        \unit_decode/RegisterFile/n1465 ), .CK(CLK), .Q(\unit_decode/n1982 ), 
        .QN(\unit_decode/RegisterFile/n3670 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][4]  ( .D(
        \unit_decode/RegisterFile/n1464 ), .CK(CLK), .Q(\unit_decode/n1983 ), 
        .QN(\unit_decode/RegisterFile/n3671 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][3]  ( .D(
        \unit_decode/RegisterFile/n1463 ), .CK(CLK), .Q(\unit_decode/n1984 ), 
        .QN(\unit_decode/RegisterFile/n3672 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][2]  ( .D(
        \unit_decode/RegisterFile/n1462 ), .CK(CLK), .Q(\unit_decode/n1985 ), 
        .QN(\unit_decode/RegisterFile/n3673 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][1]  ( .D(
        \unit_decode/RegisterFile/n1461 ), .CK(CLK), .Q(\unit_decode/n1986 ), 
        .QN(\unit_decode/RegisterFile/n3674 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[21][0]  ( .D(
        \unit_decode/RegisterFile/n1460 ), .CK(CLK), .Q(\unit_decode/n1987 ), 
        .QN(\unit_decode/RegisterFile/n3675 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][23]  ( .D(
        \unit_decode/RegisterFile/n1515 ), .CK(CLK), .Q(\unit_decode/n1988 ), 
        .QN(\unit_decode/RegisterFile/n3620 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][22]  ( .D(
        \unit_decode/RegisterFile/n1514 ), .CK(CLK), .Q(\unit_decode/n1989 ), 
        .QN(\unit_decode/RegisterFile/n3621 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][21]  ( .D(
        \unit_decode/RegisterFile/n1513 ), .CK(CLK), .Q(\unit_decode/n1990 ), 
        .QN(\unit_decode/RegisterFile/n3622 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][20]  ( .D(
        \unit_decode/RegisterFile/n1512 ), .CK(CLK), .Q(\unit_decode/n1991 ), 
        .QN(\unit_decode/RegisterFile/n3623 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][19]  ( .D(
        \unit_decode/RegisterFile/n1511 ), .CK(CLK), .Q(\unit_decode/n1992 ), 
        .QN(\unit_decode/RegisterFile/n3624 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][18]  ( .D(
        \unit_decode/RegisterFile/n1510 ), .CK(CLK), .Q(\unit_decode/n1993 ), 
        .QN(\unit_decode/RegisterFile/n3625 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][17]  ( .D(
        \unit_decode/RegisterFile/n1509 ), .CK(CLK), .Q(\unit_decode/n1994 ), 
        .QN(\unit_decode/RegisterFile/n3626 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][16]  ( .D(
        \unit_decode/RegisterFile/n1508 ), .CK(CLK), .Q(\unit_decode/n1995 ), 
        .QN(\unit_decode/RegisterFile/n3627 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][15]  ( .D(
        \unit_decode/RegisterFile/n1507 ), .CK(CLK), .Q(\unit_decode/n1996 ), 
        .QN(\unit_decode/RegisterFile/n3628 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][14]  ( .D(
        \unit_decode/RegisterFile/n1506 ), .CK(CLK), .Q(\unit_decode/n1997 ), 
        .QN(\unit_decode/RegisterFile/n3629 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][13]  ( .D(
        \unit_decode/RegisterFile/n1505 ), .CK(CLK), .Q(\unit_decode/n1998 ), 
        .QN(\unit_decode/RegisterFile/n3630 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][12]  ( .D(
        \unit_decode/RegisterFile/n1504 ), .CK(CLK), .Q(\unit_decode/n1999 ), 
        .QN(\unit_decode/RegisterFile/n3631 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][11]  ( .D(
        \unit_decode/RegisterFile/n1503 ), .CK(CLK), .Q(\unit_decode/n2000 ), 
        .QN(\unit_decode/RegisterFile/n3632 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][10]  ( .D(
        \unit_decode/RegisterFile/n1502 ), .CK(CLK), .Q(\unit_decode/n2001 ), 
        .QN(\unit_decode/RegisterFile/n3633 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][9]  ( .D(
        \unit_decode/RegisterFile/n1501 ), .CK(CLK), .Q(\unit_decode/n2002 ), 
        .QN(\unit_decode/RegisterFile/n3634 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][8]  ( .D(
        \unit_decode/RegisterFile/n1500 ), .CK(CLK), .Q(\unit_decode/n2003 ), 
        .QN(\unit_decode/RegisterFile/n3635 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][7]  ( .D(
        \unit_decode/RegisterFile/n1499 ), .CK(CLK), .Q(\unit_decode/n2004 ), 
        .QN(\unit_decode/RegisterFile/n3636 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][6]  ( .D(
        \unit_decode/RegisterFile/n1498 ), .CK(CLK), .Q(\unit_decode/n2005 ), 
        .QN(\unit_decode/RegisterFile/n3637 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][5]  ( .D(
        \unit_decode/RegisterFile/n1497 ), .CK(CLK), .Q(\unit_decode/n2006 ), 
        .QN(\unit_decode/RegisterFile/n3638 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][4]  ( .D(
        \unit_decode/RegisterFile/n1496 ), .CK(CLK), .Q(\unit_decode/n2007 ), 
        .QN(\unit_decode/RegisterFile/n3639 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][3]  ( .D(
        \unit_decode/RegisterFile/n1495 ), .CK(CLK), .Q(\unit_decode/n2008 ), 
        .QN(\unit_decode/RegisterFile/n3640 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][2]  ( .D(
        \unit_decode/RegisterFile/n1494 ), .CK(CLK), .Q(\unit_decode/n2009 ), 
        .QN(\unit_decode/RegisterFile/n3641 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][1]  ( .D(
        \unit_decode/RegisterFile/n1493 ), .CK(CLK), .Q(\unit_decode/n2010 ), 
        .QN(\unit_decode/RegisterFile/n3642 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[20][0]  ( .D(
        \unit_decode/RegisterFile/n1492 ), .CK(CLK), .Q(\unit_decode/n2011 ), 
        .QN(\unit_decode/RegisterFile/n3643 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][23]  ( .D(
        \unit_decode/RegisterFile/n1547 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3588 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][22]  ( .D(
        \unit_decode/RegisterFile/n1546 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3589 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][21]  ( .D(
        \unit_decode/RegisterFile/n1545 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3590 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][20]  ( .D(
        \unit_decode/RegisterFile/n1544 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3591 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][19]  ( .D(
        \unit_decode/RegisterFile/n1543 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3592 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][18]  ( .D(
        \unit_decode/RegisterFile/n1542 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3593 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][17]  ( .D(
        \unit_decode/RegisterFile/n1541 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3594 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][16]  ( .D(
        \unit_decode/RegisterFile/n1540 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3595 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][15]  ( .D(
        \unit_decode/RegisterFile/n1539 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3596 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][14]  ( .D(
        \unit_decode/RegisterFile/n1538 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3597 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][13]  ( .D(
        \unit_decode/RegisterFile/n1537 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3598 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][12]  ( .D(
        \unit_decode/RegisterFile/n1536 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3599 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][11]  ( .D(
        \unit_decode/RegisterFile/n1535 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3600 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][10]  ( .D(
        \unit_decode/RegisterFile/n1534 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3601 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][9]  ( .D(
        \unit_decode/RegisterFile/n1533 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3602 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][8]  ( .D(
        \unit_decode/RegisterFile/n1532 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3603 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][7]  ( .D(
        \unit_decode/RegisterFile/n1531 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3604 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][6]  ( .D(
        \unit_decode/RegisterFile/n1530 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3605 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][5]  ( .D(
        \unit_decode/RegisterFile/n1529 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3606 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][4]  ( .D(
        \unit_decode/RegisterFile/n1528 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3607 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][3]  ( .D(
        \unit_decode/RegisterFile/n1527 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3608 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][2]  ( .D(
        \unit_decode/RegisterFile/n1526 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3609 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][1]  ( .D(
        \unit_decode/RegisterFile/n1525 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3610 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[19][0]  ( .D(
        \unit_decode/RegisterFile/n1524 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3611 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][31]  ( .D(
        \unit_decode/RegisterFile/n1651 ), .CK(CLK), .Q(\unit_decode/n1783 ), 
        .QN(\unit_decode/RegisterFile/n3484 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][30]  ( .D(
        \unit_decode/RegisterFile/n1650 ), .CK(CLK), .Q(\unit_decode/n1784 ), 
        .QN(\unit_decode/RegisterFile/n3485 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][29]  ( .D(
        \unit_decode/RegisterFile/n1649 ), .CK(CLK), .Q(\unit_decode/n1785 ), 
        .QN(\unit_decode/RegisterFile/n3486 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][22]  ( .D(
        \unit_decode/RegisterFile/n1642 ), .CK(CLK), .Q(\unit_decode/n2061 ), 
        .QN(\unit_decode/RegisterFile/n3493 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][21]  ( .D(
        \unit_decode/RegisterFile/n1641 ), .CK(CLK), .Q(\unit_decode/n2062 ), 
        .QN(\unit_decode/RegisterFile/n3494 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][20]  ( .D(
        \unit_decode/RegisterFile/n1640 ), .CK(CLK), .Q(\unit_decode/n2063 ), 
        .QN(\unit_decode/RegisterFile/n3495 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][19]  ( .D(
        \unit_decode/RegisterFile/n1639 ), .CK(CLK), .Q(\unit_decode/n2064 ), 
        .QN(\unit_decode/RegisterFile/n3496 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][18]  ( .D(
        \unit_decode/RegisterFile/n1638 ), .CK(CLK), .Q(\unit_decode/n2065 ), 
        .QN(\unit_decode/RegisterFile/n3497 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][17]  ( .D(
        \unit_decode/RegisterFile/n1637 ), .CK(CLK), .Q(\unit_decode/n2066 ), 
        .QN(\unit_decode/RegisterFile/n3498 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][16]  ( .D(
        \unit_decode/RegisterFile/n1636 ), .CK(CLK), .Q(\unit_decode/n2067 ), 
        .QN(\unit_decode/RegisterFile/n3499 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][15]  ( .D(
        \unit_decode/RegisterFile/n1635 ), .CK(CLK), .Q(\unit_decode/n2068 ), 
        .QN(\unit_decode/RegisterFile/n3500 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][14]  ( .D(
        \unit_decode/RegisterFile/n1634 ), .CK(CLK), .Q(\unit_decode/n2069 ), 
        .QN(\unit_decode/RegisterFile/n3501 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][13]  ( .D(
        \unit_decode/RegisterFile/n1633 ), .CK(CLK), .Q(\unit_decode/n2070 ), 
        .QN(\unit_decode/RegisterFile/n3502 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][12]  ( .D(
        \unit_decode/RegisterFile/n1632 ), .CK(CLK), .Q(\unit_decode/n2071 ), 
        .QN(\unit_decode/RegisterFile/n3503 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][11]  ( .D(
        \unit_decode/RegisterFile/n1631 ), .CK(CLK), .Q(\unit_decode/n2072 ), 
        .QN(\unit_decode/RegisterFile/n3504 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][10]  ( .D(
        \unit_decode/RegisterFile/n1630 ), .CK(CLK), .Q(\unit_decode/n2073 ), 
        .QN(\unit_decode/RegisterFile/n3505 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][9]  ( .D(
        \unit_decode/RegisterFile/n1629 ), .CK(CLK), .Q(\unit_decode/n2074 ), 
        .QN(\unit_decode/RegisterFile/n3506 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][8]  ( .D(
        \unit_decode/RegisterFile/n1628 ), .CK(CLK), .Q(\unit_decode/n2075 ), 
        .QN(\unit_decode/RegisterFile/n3507 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][7]  ( .D(
        \unit_decode/RegisterFile/n1627 ), .CK(CLK), .Q(\unit_decode/n2076 ), 
        .QN(\unit_decode/RegisterFile/n3508 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][6]  ( .D(
        \unit_decode/RegisterFile/n1626 ), .CK(CLK), .Q(\unit_decode/n2077 ), 
        .QN(\unit_decode/RegisterFile/n3509 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][5]  ( .D(
        \unit_decode/RegisterFile/n1625 ), .CK(CLK), .Q(\unit_decode/n2078 ), 
        .QN(\unit_decode/RegisterFile/n3510 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][4]  ( .D(
        \unit_decode/RegisterFile/n1624 ), .CK(CLK), .Q(\unit_decode/n2079 ), 
        .QN(\unit_decode/RegisterFile/n3511 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][1]  ( .D(
        \unit_decode/RegisterFile/n1621 ), .CK(CLK), .Q(\unit_decode/n2082 ), 
        .QN(\unit_decode/RegisterFile/n3514 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[16][0]  ( .D(
        \unit_decode/RegisterFile/n1620 ), .CK(CLK), .Q(\unit_decode/n2083 ), 
        .QN(\unit_decode/RegisterFile/n3515 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][31]  ( .D(
        \unit_decode/RegisterFile/n1619 ), .CK(CLK), .Q(\unit_decode/n1775 ), 
        .QN(\unit_decode/RegisterFile/n3516 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][30]  ( .D(
        \unit_decode/RegisterFile/n1618 ), .CK(CLK), .Q(\unit_decode/n1776 ), 
        .QN(\unit_decode/RegisterFile/n3517 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[17][29]  ( .D(
        \unit_decode/RegisterFile/n1617 ), .CK(CLK), .Q(\unit_decode/n1777 ), 
        .QN(\unit_decode/RegisterFile/n3518 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][31]  ( .D(
        \unit_decode/RegisterFile/n1299 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3836 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][30]  ( .D(
        \unit_decode/RegisterFile/n1298 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3837 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][29]  ( .D(
        \unit_decode/RegisterFile/n1297 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3838 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][28]  ( .D(
        \unit_decode/RegisterFile/n1296 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3839 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][27]  ( .D(
        \unit_decode/RegisterFile/n1295 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3840 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][26]  ( .D(
        \unit_decode/RegisterFile/n1294 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3841 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][25]  ( .D(
        \unit_decode/RegisterFile/n1293 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3842 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[27][24]  ( .D(
        \unit_decode/RegisterFile/n1292 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3843 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][31]  ( .D(
        \unit_decode/RegisterFile/n1331 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3804 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][30]  ( .D(
        \unit_decode/RegisterFile/n1330 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3805 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][29]  ( .D(
        \unit_decode/RegisterFile/n1329 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3806 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][28]  ( .D(
        \unit_decode/RegisterFile/n1328 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3807 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][27]  ( .D(
        \unit_decode/RegisterFile/n1327 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3808 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][26]  ( .D(
        \unit_decode/RegisterFile/n1326 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3809 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][25]  ( .D(
        \unit_decode/RegisterFile/n1325 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3810 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[26][24]  ( .D(
        \unit_decode/RegisterFile/n1324 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3811 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][31]  ( .D(
        \unit_decode/RegisterFile/n1363 ), .CK(CLK), .Q(\unit_decode/n1876 ), 
        .QN(\unit_decode/RegisterFile/n3772 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][30]  ( .D(
        \unit_decode/RegisterFile/n1362 ), .CK(CLK), .Q(\unit_decode/n1877 ), 
        .QN(\unit_decode/RegisterFile/n3773 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][29]  ( .D(
        \unit_decode/RegisterFile/n1361 ), .CK(CLK), .Q(\unit_decode/n1878 ), 
        .QN(\unit_decode/RegisterFile/n3774 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][28]  ( .D(
        \unit_decode/RegisterFile/n1360 ), .CK(CLK), .Q(\unit_decode/n1879 ), 
        .QN(\unit_decode/RegisterFile/n3775 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][27]  ( .D(
        \unit_decode/RegisterFile/n1359 ), .CK(CLK), .Q(\unit_decode/n1880 ), 
        .QN(\unit_decode/RegisterFile/n3776 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][26]  ( .D(
        \unit_decode/RegisterFile/n1358 ), .CK(CLK), .Q(\unit_decode/n1881 ), 
        .QN(\unit_decode/RegisterFile/n3777 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][25]  ( .D(
        \unit_decode/RegisterFile/n1357 ), .CK(CLK), .Q(\unit_decode/n1882 ), 
        .QN(\unit_decode/RegisterFile/n3778 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[25][24]  ( .D(
        \unit_decode/RegisterFile/n1356 ), .CK(CLK), .Q(\unit_decode/n1883 ), 
        .QN(\unit_decode/RegisterFile/n3779 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][31]  ( .D(
        \unit_decode/RegisterFile/n1395 ), .CK(CLK), .Q(\unit_decode/n1884 ), 
        .QN(\unit_decode/RegisterFile/n3740 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][30]  ( .D(
        \unit_decode/RegisterFile/n1394 ), .CK(CLK), .Q(\unit_decode/n1885 ), 
        .QN(\unit_decode/RegisterFile/n3741 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][29]  ( .D(
        \unit_decode/RegisterFile/n1393 ), .CK(CLK), .Q(\unit_decode/n1886 ), 
        .QN(\unit_decode/RegisterFile/n3742 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][28]  ( .D(
        \unit_decode/RegisterFile/n1392 ), .CK(CLK), .Q(\unit_decode/n1887 ), 
        .QN(\unit_decode/RegisterFile/n3743 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][27]  ( .D(
        \unit_decode/RegisterFile/n1391 ), .CK(CLK), .Q(\unit_decode/n1888 ), 
        .QN(\unit_decode/RegisterFile/n3744 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][26]  ( .D(
        \unit_decode/RegisterFile/n1390 ), .CK(CLK), .Q(\unit_decode/n1889 ), 
        .QN(\unit_decode/RegisterFile/n3745 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][25]  ( .D(
        \unit_decode/RegisterFile/n1389 ), .CK(CLK), .Q(\unit_decode/n1890 ), 
        .QN(\unit_decode/RegisterFile/n3746 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[24][24]  ( .D(
        \unit_decode/RegisterFile/n1388 ), .CK(CLK), .Q(\unit_decode/n1891 ), 
        .QN(\unit_decode/RegisterFile/n3747 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][31]  ( .D(
        \unit_decode/RegisterFile/n1267 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3868 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][30]  ( .D(
        \unit_decode/RegisterFile/n1266 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3869 ) );
  DFF_X1 \unit_decode/RegisterFile/REGISTERS_reg[28][29]  ( .D(
        \unit_decode/RegisterFile/n1265 ), .CK(CLK), .QN(
        \unit_decode/RegisterFile/n3870 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][31]  ( .D(
        \unit_memory/DRAM/n1316 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n353 ), .QN(\unit_memory/DRAM/n3231 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][30]  ( .D(
        \unit_memory/DRAM/n1315 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n354 ), .QN(\unit_memory/DRAM/n3232 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][29]  ( .D(
        \unit_memory/DRAM/n1314 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n355 ), .QN(\unit_memory/DRAM/n3233 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][28]  ( .D(
        \unit_memory/DRAM/n1313 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n356 ), .QN(\unit_memory/DRAM/n3234 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][27]  ( .D(
        \unit_memory/DRAM/n1312 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n357 ), .QN(\unit_memory/DRAM/n3235 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][26]  ( .D(
        \unit_memory/DRAM/n1311 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n358 ), .QN(\unit_memory/DRAM/n3236 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][25]  ( .D(
        \unit_memory/DRAM/n1310 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n359 ), .QN(\unit_memory/DRAM/n3237 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][24]  ( .D(
        \unit_memory/DRAM/n1309 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n360 ), .QN(\unit_memory/DRAM/n3238 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][31]  ( .D(
        \unit_memory/DRAM/n1444 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n225 ), .QN(\unit_memory/DRAM/n3103 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][30]  ( .D(
        \unit_memory/DRAM/n1443 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n226 ), .QN(\unit_memory/DRAM/n3104 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][29]  ( .D(
        \unit_memory/DRAM/n1442 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n227 ), .QN(\unit_memory/DRAM/n3105 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][28]  ( .D(
        \unit_memory/DRAM/n1441 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n228 ), .QN(\unit_memory/DRAM/n3106 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][27]  ( .D(
        \unit_memory/DRAM/n1440 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n229 ), .QN(\unit_memory/DRAM/n3107 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][26]  ( .D(
        \unit_memory/DRAM/n1439 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n230 ), .QN(\unit_memory/DRAM/n3108 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][25]  ( .D(
        \unit_memory/DRAM/n1438 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n231 ), .QN(\unit_memory/DRAM/n3109 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][24]  ( .D(
        \unit_memory/DRAM/n1437 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n232 ), .QN(\unit_memory/DRAM/n3110 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][31]  ( .D(
        \unit_memory/DRAM/n1572 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n97 ), .QN(\unit_memory/DRAM/n2975 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][30]  ( .D(
        \unit_memory/DRAM/n1571 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n98 ), .QN(\unit_memory/DRAM/n2976 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][29]  ( .D(
        \unit_memory/DRAM/n1570 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n99 ), .QN(\unit_memory/DRAM/n2977 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][28]  ( .D(
        \unit_memory/DRAM/n1569 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n100 ), .QN(\unit_memory/DRAM/n2978 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][27]  ( .D(
        \unit_memory/DRAM/n1568 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n101 ), .QN(\unit_memory/DRAM/n2979 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][26]  ( .D(
        \unit_memory/DRAM/n1567 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n102 ), .QN(\unit_memory/DRAM/n2980 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][25]  ( .D(
        \unit_memory/DRAM/n1566 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n103 ), .QN(\unit_memory/DRAM/n2981 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][24]  ( .D(
        \unit_memory/DRAM/n1565 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n104 ), .QN(\unit_memory/DRAM/n2982 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][31]  ( .D(
        \unit_memory/DRAM/n1700 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2847 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][30]  ( .D(
        \unit_memory/DRAM/n1699 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2848 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][29]  ( .D(
        \unit_memory/DRAM/n1698 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2849 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][28]  ( .D(
        \unit_memory/DRAM/n1697 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2850 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][27]  ( .D(
        \unit_memory/DRAM/n1696 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2851 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][26]  ( .D(
        \unit_memory/DRAM/n1695 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2852 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][25]  ( .D(
        \unit_memory/DRAM/n1694 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2853 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][24]  ( .D(
        \unit_memory/DRAM/n1693 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2854 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][31]  ( .D(
        \unit_memory/DRAM/n1828 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2719 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][30]  ( .D(
        \unit_memory/DRAM/n1827 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2720 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][29]  ( .D(
        \unit_memory/DRAM/n1826 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2721 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][28]  ( .D(
        \unit_memory/DRAM/n1825 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2722 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][27]  ( .D(
        \unit_memory/DRAM/n1824 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2723 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][26]  ( .D(
        \unit_memory/DRAM/n1823 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2724 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][25]  ( .D(
        \unit_memory/DRAM/n1822 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2725 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][24]  ( .D(
        \unit_memory/DRAM/n1821 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2726 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][31]  ( .D(\unit_memory/DRAM/n1956 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2591 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][30]  ( .D(\unit_memory/DRAM/n1955 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2592 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][29]  ( .D(\unit_memory/DRAM/n1954 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2593 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][28]  ( .D(\unit_memory/DRAM/n1953 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2594 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][27]  ( .D(\unit_memory/DRAM/n1952 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2595 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][26]  ( .D(\unit_memory/DRAM/n1951 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2596 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][25]  ( .D(\unit_memory/DRAM/n1950 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2597 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][24]  ( .D(\unit_memory/DRAM/n1949 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2598 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][31]  ( .D(\unit_memory/DRAM/n2084 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2463 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][30]  ( .D(\unit_memory/DRAM/n2083 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2464 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][29]  ( .D(\unit_memory/DRAM/n2082 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2465 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][28]  ( .D(\unit_memory/DRAM/n2081 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2466 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][27]  ( .D(\unit_memory/DRAM/n2080 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2467 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][26]  ( .D(\unit_memory/DRAM/n2079 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2468 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][25]  ( .D(\unit_memory/DRAM/n2078 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2469 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][24]  ( .D(\unit_memory/DRAM/n2077 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2470 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][23]  ( .D(
        \unit_memory/DRAM/n1308 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n361 ), .QN(\unit_memory/DRAM/n3239 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][22]  ( .D(
        \unit_memory/DRAM/n1307 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n362 ), .QN(\unit_memory/DRAM/n3240 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][21]  ( .D(
        \unit_memory/DRAM/n1306 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n363 ), .QN(\unit_memory/DRAM/n3241 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][20]  ( .D(
        \unit_memory/DRAM/n1305 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n364 ), .QN(\unit_memory/DRAM/n3242 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][19]  ( .D(
        \unit_memory/DRAM/n1304 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n365 ), .QN(\unit_memory/DRAM/n3243 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][18]  ( .D(
        \unit_memory/DRAM/n1303 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n366 ), .QN(\unit_memory/DRAM/n3244 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][17]  ( .D(
        \unit_memory/DRAM/n1302 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n367 ), .QN(\unit_memory/DRAM/n3245 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][16]  ( .D(
        \unit_memory/DRAM/n1301 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n368 ), .QN(\unit_memory/DRAM/n3246 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][15]  ( .D(
        \unit_memory/DRAM/n1300 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n369 ), .QN(\unit_memory/DRAM/n3247 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][14]  ( .D(
        \unit_memory/DRAM/n1299 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n370 ), .QN(\unit_memory/DRAM/n3248 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][13]  ( .D(
        \unit_memory/DRAM/n1298 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n371 ), .QN(\unit_memory/DRAM/n3249 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][12]  ( .D(
        \unit_memory/DRAM/n1297 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n372 ), .QN(\unit_memory/DRAM/n3250 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][11]  ( .D(
        \unit_memory/DRAM/n1296 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n373 ), .QN(\unit_memory/DRAM/n3251 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][10]  ( .D(
        \unit_memory/DRAM/n1295 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n374 ), .QN(\unit_memory/DRAM/n3252 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][9]  ( .D(\unit_memory/DRAM/n1294 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n375 ), .QN(
        \unit_memory/DRAM/n3253 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][8]  ( .D(\unit_memory/DRAM/n1293 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n376 ), .QN(
        \unit_memory/DRAM/n3254 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][7]  ( .D(\unit_memory/DRAM/n1292 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n377 ), .QN(
        \unit_memory/DRAM/n3255 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][6]  ( .D(\unit_memory/DRAM/n1291 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n378 ), .QN(
        \unit_memory/DRAM/n3256 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][5]  ( .D(\unit_memory/DRAM/n1290 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n379 ), .QN(
        \unit_memory/DRAM/n3257 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][4]  ( .D(\unit_memory/DRAM/n1289 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n380 ), .QN(
        \unit_memory/DRAM/n3258 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][3]  ( .D(\unit_memory/DRAM/n1288 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n381 ), .QN(
        \unit_memory/DRAM/n3259 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][2]  ( .D(\unit_memory/DRAM/n1287 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n382 ), .QN(
        \unit_memory/DRAM/n3260 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][1]  ( .D(\unit_memory/DRAM/n1286 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n383 ), .QN(
        \unit_memory/DRAM/n3261 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[27][0]  ( .D(\unit_memory/DRAM/n1285 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n384 ), .QN(
        \unit_memory/DRAM/n3262 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][23]  ( .D(
        \unit_memory/DRAM/n1436 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n233 ), .QN(\unit_memory/DRAM/n3111 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][22]  ( .D(
        \unit_memory/DRAM/n1435 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n234 ), .QN(\unit_memory/DRAM/n3112 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][21]  ( .D(
        \unit_memory/DRAM/n1434 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n235 ), .QN(\unit_memory/DRAM/n3113 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][20]  ( .D(
        \unit_memory/DRAM/n1433 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n236 ), .QN(\unit_memory/DRAM/n3114 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][19]  ( .D(
        \unit_memory/DRAM/n1432 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n237 ), .QN(\unit_memory/DRAM/n3115 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][18]  ( .D(
        \unit_memory/DRAM/n1431 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n238 ), .QN(\unit_memory/DRAM/n3116 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][17]  ( .D(
        \unit_memory/DRAM/n1430 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n239 ), .QN(\unit_memory/DRAM/n3117 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][16]  ( .D(
        \unit_memory/DRAM/n1429 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n240 ), .QN(\unit_memory/DRAM/n3118 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][15]  ( .D(
        \unit_memory/DRAM/n1428 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n241 ), .QN(\unit_memory/DRAM/n3119 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][14]  ( .D(
        \unit_memory/DRAM/n1427 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n242 ), .QN(\unit_memory/DRAM/n3120 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][13]  ( .D(
        \unit_memory/DRAM/n1426 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n243 ), .QN(\unit_memory/DRAM/n3121 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][12]  ( .D(
        \unit_memory/DRAM/n1425 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n244 ), .QN(\unit_memory/DRAM/n3122 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][11]  ( .D(
        \unit_memory/DRAM/n1424 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n245 ), .QN(\unit_memory/DRAM/n3123 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][10]  ( .D(
        \unit_memory/DRAM/n1423 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n246 ), .QN(\unit_memory/DRAM/n3124 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][9]  ( .D(\unit_memory/DRAM/n1422 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n247 ), .QN(
        \unit_memory/DRAM/n3125 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][8]  ( .D(\unit_memory/DRAM/n1421 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n248 ), .QN(
        \unit_memory/DRAM/n3126 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][7]  ( .D(\unit_memory/DRAM/n1420 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n249 ), .QN(
        \unit_memory/DRAM/n3127 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][6]  ( .D(\unit_memory/DRAM/n1419 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n250 ), .QN(
        \unit_memory/DRAM/n3128 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][5]  ( .D(\unit_memory/DRAM/n1418 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n251 ), .QN(
        \unit_memory/DRAM/n3129 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][4]  ( .D(\unit_memory/DRAM/n1417 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n252 ), .QN(
        \unit_memory/DRAM/n3130 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][3]  ( .D(\unit_memory/DRAM/n1416 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n253 ), .QN(
        \unit_memory/DRAM/n3131 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][2]  ( .D(\unit_memory/DRAM/n1415 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n254 ), .QN(
        \unit_memory/DRAM/n3132 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][1]  ( .D(\unit_memory/DRAM/n1414 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n255 ), .QN(
        \unit_memory/DRAM/n3133 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[23][0]  ( .D(\unit_memory/DRAM/n1413 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n256 ), .QN(
        \unit_memory/DRAM/n3134 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][23]  ( .D(
        \unit_memory/DRAM/n1564 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n105 ), .QN(\unit_memory/DRAM/n2983 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][22]  ( .D(
        \unit_memory/DRAM/n1563 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n106 ), .QN(\unit_memory/DRAM/n2984 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][21]  ( .D(
        \unit_memory/DRAM/n1562 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n107 ), .QN(\unit_memory/DRAM/n2985 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][20]  ( .D(
        \unit_memory/DRAM/n1561 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n108 ), .QN(\unit_memory/DRAM/n2986 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][19]  ( .D(
        \unit_memory/DRAM/n1560 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n109 ), .QN(\unit_memory/DRAM/n2987 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][18]  ( .D(
        \unit_memory/DRAM/n1559 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n110 ), .QN(\unit_memory/DRAM/n2988 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][17]  ( .D(
        \unit_memory/DRAM/n1558 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n111 ), .QN(\unit_memory/DRAM/n2989 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][16]  ( .D(
        \unit_memory/DRAM/n1557 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n112 ), .QN(\unit_memory/DRAM/n2990 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][15]  ( .D(
        \unit_memory/DRAM/n1556 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n113 ), .QN(\unit_memory/DRAM/n2991 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][14]  ( .D(
        \unit_memory/DRAM/n1555 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n114 ), .QN(\unit_memory/DRAM/n2992 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][13]  ( .D(
        \unit_memory/DRAM/n1554 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n115 ), .QN(\unit_memory/DRAM/n2993 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][12]  ( .D(
        \unit_memory/DRAM/n1553 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n116 ), .QN(\unit_memory/DRAM/n2994 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][11]  ( .D(
        \unit_memory/DRAM/n1552 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n117 ), .QN(\unit_memory/DRAM/n2995 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][10]  ( .D(
        \unit_memory/DRAM/n1551 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n118 ), .QN(\unit_memory/DRAM/n2996 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][9]  ( .D(\unit_memory/DRAM/n1550 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n119 ), .QN(
        \unit_memory/DRAM/n2997 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][8]  ( .D(\unit_memory/DRAM/n1549 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n120 ), .QN(
        \unit_memory/DRAM/n2998 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][7]  ( .D(\unit_memory/DRAM/n1548 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n121 ), .QN(
        \unit_memory/DRAM/n2999 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][6]  ( .D(\unit_memory/DRAM/n1547 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n122 ), .QN(
        \unit_memory/DRAM/n3000 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][5]  ( .D(\unit_memory/DRAM/n1546 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n123 ), .QN(
        \unit_memory/DRAM/n3001 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][4]  ( .D(\unit_memory/DRAM/n1545 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n124 ), .QN(
        \unit_memory/DRAM/n3002 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][3]  ( .D(\unit_memory/DRAM/n1544 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n125 ), .QN(
        \unit_memory/DRAM/n3003 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][2]  ( .D(\unit_memory/DRAM/n1543 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n126 ), .QN(
        \unit_memory/DRAM/n3004 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][1]  ( .D(\unit_memory/DRAM/n1542 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n127 ), .QN(
        \unit_memory/DRAM/n3005 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[19][0]  ( .D(\unit_memory/DRAM/n1541 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n128 ), .QN(
        \unit_memory/DRAM/n3006 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][23]  ( .D(
        \unit_memory/DRAM/n1692 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2855 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][22]  ( .D(
        \unit_memory/DRAM/n1691 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2856 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][21]  ( .D(
        \unit_memory/DRAM/n1690 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2857 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][20]  ( .D(
        \unit_memory/DRAM/n1689 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2858 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][19]  ( .D(
        \unit_memory/DRAM/n1688 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2859 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][18]  ( .D(
        \unit_memory/DRAM/n1687 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2860 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][17]  ( .D(
        \unit_memory/DRAM/n1686 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2861 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][16]  ( .D(
        \unit_memory/DRAM/n1685 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2862 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][15]  ( .D(
        \unit_memory/DRAM/n1684 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2863 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][14]  ( .D(
        \unit_memory/DRAM/n1683 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2864 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][13]  ( .D(
        \unit_memory/DRAM/n1682 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2865 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][12]  ( .D(
        \unit_memory/DRAM/n1681 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2866 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][11]  ( .D(
        \unit_memory/DRAM/n1680 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2867 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][10]  ( .D(
        \unit_memory/DRAM/n1679 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2868 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][9]  ( .D(\unit_memory/DRAM/n1678 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2869 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][8]  ( .D(\unit_memory/DRAM/n1677 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2870 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][7]  ( .D(\unit_memory/DRAM/n1676 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2871 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][6]  ( .D(\unit_memory/DRAM/n1675 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2872 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][5]  ( .D(\unit_memory/DRAM/n1674 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2873 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][4]  ( .D(\unit_memory/DRAM/n1673 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2874 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][3]  ( .D(\unit_memory/DRAM/n1672 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2875 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][2]  ( .D(\unit_memory/DRAM/n1671 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2876 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][1]  ( .D(\unit_memory/DRAM/n1670 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2877 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[15][0]  ( .D(\unit_memory/DRAM/n1669 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2878 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][23]  ( .D(
        \unit_memory/DRAM/n1820 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2727 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][22]  ( .D(
        \unit_memory/DRAM/n1819 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2728 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][21]  ( .D(
        \unit_memory/DRAM/n1818 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2729 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][20]  ( .D(
        \unit_memory/DRAM/n1817 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2730 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][19]  ( .D(
        \unit_memory/DRAM/n1816 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2731 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][18]  ( .D(
        \unit_memory/DRAM/n1815 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2732 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][17]  ( .D(
        \unit_memory/DRAM/n1814 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2733 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][16]  ( .D(
        \unit_memory/DRAM/n1813 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2734 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][15]  ( .D(
        \unit_memory/DRAM/n1812 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2735 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][14]  ( .D(
        \unit_memory/DRAM/n1811 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2736 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][13]  ( .D(
        \unit_memory/DRAM/n1810 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2737 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][12]  ( .D(
        \unit_memory/DRAM/n1809 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2738 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][11]  ( .D(
        \unit_memory/DRAM/n1808 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2739 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][10]  ( .D(
        \unit_memory/DRAM/n1807 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2740 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][9]  ( .D(\unit_memory/DRAM/n1806 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2741 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][8]  ( .D(\unit_memory/DRAM/n1805 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2742 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][7]  ( .D(\unit_memory/DRAM/n1804 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2743 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][6]  ( .D(\unit_memory/DRAM/n1803 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2744 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][5]  ( .D(\unit_memory/DRAM/n1802 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2745 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][4]  ( .D(\unit_memory/DRAM/n1801 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2746 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][3]  ( .D(\unit_memory/DRAM/n1800 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2747 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][2]  ( .D(\unit_memory/DRAM/n1799 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2748 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][1]  ( .D(\unit_memory/DRAM/n1798 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2749 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[11][0]  ( .D(\unit_memory/DRAM/n1797 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2750 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][23]  ( .D(\unit_memory/DRAM/n1948 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2599 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][22]  ( .D(\unit_memory/DRAM/n1947 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2600 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][21]  ( .D(\unit_memory/DRAM/n1946 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2601 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][20]  ( .D(\unit_memory/DRAM/n1945 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2602 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][19]  ( .D(\unit_memory/DRAM/n1944 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2603 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][18]  ( .D(\unit_memory/DRAM/n1943 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2604 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][17]  ( .D(\unit_memory/DRAM/n1942 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2605 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][16]  ( .D(\unit_memory/DRAM/n1941 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2606 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][15]  ( .D(\unit_memory/DRAM/n1940 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2607 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][14]  ( .D(\unit_memory/DRAM/n1939 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2608 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][13]  ( .D(\unit_memory/DRAM/n1938 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2609 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][12]  ( .D(\unit_memory/DRAM/n1937 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2610 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][11]  ( .D(\unit_memory/DRAM/n1936 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2611 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][10]  ( .D(\unit_memory/DRAM/n1935 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2612 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][9]  ( .D(\unit_memory/DRAM/n1934 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2613 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][8]  ( .D(\unit_memory/DRAM/n1933 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2614 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][7]  ( .D(\unit_memory/DRAM/n1932 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2615 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][6]  ( .D(\unit_memory/DRAM/n1931 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2616 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][5]  ( .D(\unit_memory/DRAM/n1930 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2617 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][4]  ( .D(\unit_memory/DRAM/n1929 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2618 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][3]  ( .D(\unit_memory/DRAM/n1928 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2619 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][2]  ( .D(\unit_memory/DRAM/n1927 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2620 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][1]  ( .D(\unit_memory/DRAM/n1926 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2621 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[7][0]  ( .D(\unit_memory/DRAM/n1925 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2622 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][23]  ( .D(\unit_memory/DRAM/n2076 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2471 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][22]  ( .D(\unit_memory/DRAM/n2075 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2472 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][21]  ( .D(\unit_memory/DRAM/n2074 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2473 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][20]  ( .D(\unit_memory/DRAM/n2073 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2474 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][19]  ( .D(\unit_memory/DRAM/n2072 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2475 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][18]  ( .D(\unit_memory/DRAM/n2071 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2476 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][17]  ( .D(\unit_memory/DRAM/n2070 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2477 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][16]  ( .D(\unit_memory/DRAM/n2069 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2478 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][15]  ( .D(\unit_memory/DRAM/n2068 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2479 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][14]  ( .D(\unit_memory/DRAM/n2067 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2480 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][13]  ( .D(\unit_memory/DRAM/n2066 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2481 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][12]  ( .D(\unit_memory/DRAM/n2065 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2482 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][11]  ( .D(\unit_memory/DRAM/n2064 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2483 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][10]  ( .D(\unit_memory/DRAM/n2063 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2484 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][9]  ( .D(\unit_memory/DRAM/n2062 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2485 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][8]  ( .D(\unit_memory/DRAM/n2061 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2486 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][7]  ( .D(\unit_memory/DRAM/n2060 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2487 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][6]  ( .D(\unit_memory/DRAM/n2059 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2488 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][5]  ( .D(\unit_memory/DRAM/n2058 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2489 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][4]  ( .D(\unit_memory/DRAM/n2057 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2490 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][3]  ( .D(\unit_memory/DRAM/n2056 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2491 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][2]  ( .D(\unit_memory/DRAM/n2055 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2492 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][1]  ( .D(\unit_memory/DRAM/n2054 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2493 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[3][0]  ( .D(\unit_memory/DRAM/n2053 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2494 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][7]  ( .D(\unit_memory/DRAM/n1164 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n505 ), .QN(
        \unit_memory/DRAM/n3383 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][6]  ( .D(\unit_memory/DRAM/n1163 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n506 ), .QN(
        \unit_memory/DRAM/n3384 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][5]  ( .D(\unit_memory/DRAM/n1162 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n507 ), .QN(
        \unit_memory/DRAM/n3385 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][4]  ( .D(\unit_memory/DRAM/n1161 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n508 ), .QN(
        \unit_memory/DRAM/n3386 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][3]  ( .D(\unit_memory/DRAM/n1160 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n509 ), .QN(
        \unit_memory/DRAM/n3387 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][2]  ( .D(\unit_memory/DRAM/n1159 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n510 ), .QN(
        \unit_memory/DRAM/n3388 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][1]  ( .D(\unit_memory/DRAM/n1158 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n511 ), .QN(
        \unit_memory/DRAM/n3389 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][0]  ( .D(\unit_memory/DRAM/n1157 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n512 ), .QN(
        \unit_memory/DRAM/n3390 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][31]  ( .D(
        \unit_memory/DRAM/n1284 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n385 ), .QN(\unit_memory/DRAM/n3263 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][30]  ( .D(
        \unit_memory/DRAM/n1283 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n386 ), .QN(\unit_memory/DRAM/n3264 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][29]  ( .D(
        \unit_memory/DRAM/n1282 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n387 ), .QN(\unit_memory/DRAM/n3265 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][28]  ( .D(
        \unit_memory/DRAM/n1281 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n388 ), .QN(\unit_memory/DRAM/n3266 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][27]  ( .D(
        \unit_memory/DRAM/n1280 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n389 ), .QN(\unit_memory/DRAM/n3267 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][26]  ( .D(
        \unit_memory/DRAM/n1279 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n390 ), .QN(\unit_memory/DRAM/n3268 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][25]  ( .D(
        \unit_memory/DRAM/n1278 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n391 ), .QN(\unit_memory/DRAM/n3269 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][24]  ( .D(
        \unit_memory/DRAM/n1277 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n392 ), .QN(\unit_memory/DRAM/n3270 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][31]  ( .D(
        \unit_memory/DRAM/n1412 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n257 ), .QN(\unit_memory/DRAM/n3135 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][30]  ( .D(
        \unit_memory/DRAM/n1411 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n258 ), .QN(\unit_memory/DRAM/n3136 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][29]  ( .D(
        \unit_memory/DRAM/n1410 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n259 ), .QN(\unit_memory/DRAM/n3137 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][28]  ( .D(
        \unit_memory/DRAM/n1409 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n260 ), .QN(\unit_memory/DRAM/n3138 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][27]  ( .D(
        \unit_memory/DRAM/n1408 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n261 ), .QN(\unit_memory/DRAM/n3139 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][26]  ( .D(
        \unit_memory/DRAM/n1407 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n262 ), .QN(\unit_memory/DRAM/n3140 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][25]  ( .D(
        \unit_memory/DRAM/n1406 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n263 ), .QN(\unit_memory/DRAM/n3141 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][24]  ( .D(
        \unit_memory/DRAM/n1405 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n264 ), .QN(\unit_memory/DRAM/n3142 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][31]  ( .D(
        \unit_memory/DRAM/n1540 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n129 ), .QN(\unit_memory/DRAM/n3007 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][30]  ( .D(
        \unit_memory/DRAM/n1539 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n130 ), .QN(\unit_memory/DRAM/n3008 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][29]  ( .D(
        \unit_memory/DRAM/n1538 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n131 ), .QN(\unit_memory/DRAM/n3009 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][28]  ( .D(
        \unit_memory/DRAM/n1537 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n132 ), .QN(\unit_memory/DRAM/n3010 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][27]  ( .D(
        \unit_memory/DRAM/n1536 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n133 ), .QN(\unit_memory/DRAM/n3011 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][26]  ( .D(
        \unit_memory/DRAM/n1535 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n134 ), .QN(\unit_memory/DRAM/n3012 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][25]  ( .D(
        \unit_memory/DRAM/n1534 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n135 ), .QN(\unit_memory/DRAM/n3013 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][24]  ( .D(
        \unit_memory/DRAM/n1533 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n136 ), .QN(\unit_memory/DRAM/n3014 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][31]  ( .D(
        \unit_memory/DRAM/n1668 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n1 ), .QN(\unit_memory/DRAM/n2879 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][30]  ( .D(
        \unit_memory/DRAM/n1667 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n2 ), .QN(\unit_memory/DRAM/n2880 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][29]  ( .D(
        \unit_memory/DRAM/n1666 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n3 ), .QN(\unit_memory/DRAM/n2881 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][28]  ( .D(
        \unit_memory/DRAM/n1665 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n4 ), .QN(\unit_memory/DRAM/n2882 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][27]  ( .D(
        \unit_memory/DRAM/n1664 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n5 ), .QN(\unit_memory/DRAM/n2883 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][26]  ( .D(
        \unit_memory/DRAM/n1663 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n6 ), .QN(\unit_memory/DRAM/n2884 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][25]  ( .D(
        \unit_memory/DRAM/n1662 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n7 ), .QN(\unit_memory/DRAM/n2885 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][24]  ( .D(
        \unit_memory/DRAM/n1661 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n8 ), .QN(\unit_memory/DRAM/n2886 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][31]  ( .D(
        \unit_memory/DRAM/n1796 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2751 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][30]  ( .D(
        \unit_memory/DRAM/n1795 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2752 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][29]  ( .D(
        \unit_memory/DRAM/n1794 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2753 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][28]  ( .D(
        \unit_memory/DRAM/n1793 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2754 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][27]  ( .D(
        \unit_memory/DRAM/n1792 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2755 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][26]  ( .D(
        \unit_memory/DRAM/n1791 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2756 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][25]  ( .D(
        \unit_memory/DRAM/n1790 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2757 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][24]  ( .D(
        \unit_memory/DRAM/n1789 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2758 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][31]  ( .D(\unit_memory/DRAM/n1924 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2623 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][30]  ( .D(\unit_memory/DRAM/n1923 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2624 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][29]  ( .D(\unit_memory/DRAM/n1922 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2625 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][28]  ( .D(\unit_memory/DRAM/n1921 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2626 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][27]  ( .D(\unit_memory/DRAM/n1920 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2627 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][26]  ( .D(\unit_memory/DRAM/n1919 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2628 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][25]  ( .D(\unit_memory/DRAM/n1918 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2629 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][24]  ( .D(\unit_memory/DRAM/n1917 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2630 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][31]  ( .D(\unit_memory/DRAM/n2052 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2495 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][30]  ( .D(\unit_memory/DRAM/n2051 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2496 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][29]  ( .D(\unit_memory/DRAM/n2050 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2497 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][28]  ( .D(\unit_memory/DRAM/n2049 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2498 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][27]  ( .D(\unit_memory/DRAM/n2048 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2499 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][26]  ( .D(\unit_memory/DRAM/n2047 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2500 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][25]  ( .D(\unit_memory/DRAM/n2046 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2501 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][24]  ( .D(\unit_memory/DRAM/n2045 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2502 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][23]  ( .D(
        \unit_memory/DRAM/n1276 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n393 ), .QN(\unit_memory/DRAM/n3271 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][22]  ( .D(
        \unit_memory/DRAM/n1275 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n394 ), .QN(\unit_memory/DRAM/n3272 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][21]  ( .D(
        \unit_memory/DRAM/n1274 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n395 ), .QN(\unit_memory/DRAM/n3273 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][20]  ( .D(
        \unit_memory/DRAM/n1273 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n396 ), .QN(\unit_memory/DRAM/n3274 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][19]  ( .D(
        \unit_memory/DRAM/n1272 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n397 ), .QN(\unit_memory/DRAM/n3275 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][18]  ( .D(
        \unit_memory/DRAM/n1271 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n398 ), .QN(\unit_memory/DRAM/n3276 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][17]  ( .D(
        \unit_memory/DRAM/n1270 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n399 ), .QN(\unit_memory/DRAM/n3277 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][16]  ( .D(
        \unit_memory/DRAM/n1269 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n400 ), .QN(\unit_memory/DRAM/n3278 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][15]  ( .D(
        \unit_memory/DRAM/n1268 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n401 ), .QN(\unit_memory/DRAM/n3279 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][14]  ( .D(
        \unit_memory/DRAM/n1267 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n402 ), .QN(\unit_memory/DRAM/n3280 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][13]  ( .D(
        \unit_memory/DRAM/n1266 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n403 ), .QN(\unit_memory/DRAM/n3281 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][12]  ( .D(
        \unit_memory/DRAM/n1265 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n404 ), .QN(\unit_memory/DRAM/n3282 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][11]  ( .D(
        \unit_memory/DRAM/n1264 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n405 ), .QN(\unit_memory/DRAM/n3283 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][10]  ( .D(
        \unit_memory/DRAM/n1263 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n406 ), .QN(\unit_memory/DRAM/n3284 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][9]  ( .D(\unit_memory/DRAM/n1262 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n407 ), .QN(
        \unit_memory/DRAM/n3285 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][8]  ( .D(\unit_memory/DRAM/n1261 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n408 ), .QN(
        \unit_memory/DRAM/n3286 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][7]  ( .D(\unit_memory/DRAM/n1260 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n409 ), .QN(
        \unit_memory/DRAM/n3287 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][6]  ( .D(\unit_memory/DRAM/n1259 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n410 ), .QN(
        \unit_memory/DRAM/n3288 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][5]  ( .D(\unit_memory/DRAM/n1258 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n411 ), .QN(
        \unit_memory/DRAM/n3289 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][4]  ( .D(\unit_memory/DRAM/n1257 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n412 ), .QN(
        \unit_memory/DRAM/n3290 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][3]  ( .D(\unit_memory/DRAM/n1256 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n413 ), .QN(
        \unit_memory/DRAM/n3291 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][2]  ( .D(\unit_memory/DRAM/n1255 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n414 ), .QN(
        \unit_memory/DRAM/n3292 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][1]  ( .D(\unit_memory/DRAM/n1254 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n415 ), .QN(
        \unit_memory/DRAM/n3293 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[28][0]  ( .D(\unit_memory/DRAM/n1253 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n416 ), .QN(
        \unit_memory/DRAM/n3294 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][23]  ( .D(
        \unit_memory/DRAM/n1404 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n265 ), .QN(\unit_memory/DRAM/n3143 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][22]  ( .D(
        \unit_memory/DRAM/n1403 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n266 ), .QN(\unit_memory/DRAM/n3144 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][21]  ( .D(
        \unit_memory/DRAM/n1402 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n267 ), .QN(\unit_memory/DRAM/n3145 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][20]  ( .D(
        \unit_memory/DRAM/n1401 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n268 ), .QN(\unit_memory/DRAM/n3146 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][19]  ( .D(
        \unit_memory/DRAM/n1400 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n269 ), .QN(\unit_memory/DRAM/n3147 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][18]  ( .D(
        \unit_memory/DRAM/n1399 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n270 ), .QN(\unit_memory/DRAM/n3148 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][17]  ( .D(
        \unit_memory/DRAM/n1398 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n271 ), .QN(\unit_memory/DRAM/n3149 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][16]  ( .D(
        \unit_memory/DRAM/n1397 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n272 ), .QN(\unit_memory/DRAM/n3150 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][15]  ( .D(
        \unit_memory/DRAM/n1396 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n273 ), .QN(\unit_memory/DRAM/n3151 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][14]  ( .D(
        \unit_memory/DRAM/n1395 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n274 ), .QN(\unit_memory/DRAM/n3152 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][13]  ( .D(
        \unit_memory/DRAM/n1394 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n275 ), .QN(\unit_memory/DRAM/n3153 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][12]  ( .D(
        \unit_memory/DRAM/n1393 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n276 ), .QN(\unit_memory/DRAM/n3154 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][11]  ( .D(
        \unit_memory/DRAM/n1392 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n277 ), .QN(\unit_memory/DRAM/n3155 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][10]  ( .D(
        \unit_memory/DRAM/n1391 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n278 ), .QN(\unit_memory/DRAM/n3156 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][9]  ( .D(\unit_memory/DRAM/n1390 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n279 ), .QN(
        \unit_memory/DRAM/n3157 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][8]  ( .D(\unit_memory/DRAM/n1389 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n280 ), .QN(
        \unit_memory/DRAM/n3158 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][7]  ( .D(\unit_memory/DRAM/n1388 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n281 ), .QN(
        \unit_memory/DRAM/n3159 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][6]  ( .D(\unit_memory/DRAM/n1387 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n282 ), .QN(
        \unit_memory/DRAM/n3160 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][5]  ( .D(\unit_memory/DRAM/n1386 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n283 ), .QN(
        \unit_memory/DRAM/n3161 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][4]  ( .D(\unit_memory/DRAM/n1385 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n284 ), .QN(
        \unit_memory/DRAM/n3162 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][3]  ( .D(\unit_memory/DRAM/n1384 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n285 ), .QN(
        \unit_memory/DRAM/n3163 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][2]  ( .D(\unit_memory/DRAM/n1383 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n286 ), .QN(
        \unit_memory/DRAM/n3164 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][1]  ( .D(\unit_memory/DRAM/n1382 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n287 ), .QN(
        \unit_memory/DRAM/n3165 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[24][0]  ( .D(\unit_memory/DRAM/n1381 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n288 ), .QN(
        \unit_memory/DRAM/n3166 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][23]  ( .D(
        \unit_memory/DRAM/n1532 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n137 ), .QN(\unit_memory/DRAM/n3015 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][22]  ( .D(
        \unit_memory/DRAM/n1531 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n138 ), .QN(\unit_memory/DRAM/n3016 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][21]  ( .D(
        \unit_memory/DRAM/n1530 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n139 ), .QN(\unit_memory/DRAM/n3017 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][20]  ( .D(
        \unit_memory/DRAM/n1529 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n140 ), .QN(\unit_memory/DRAM/n3018 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][19]  ( .D(
        \unit_memory/DRAM/n1528 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n141 ), .QN(\unit_memory/DRAM/n3019 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][18]  ( .D(
        \unit_memory/DRAM/n1527 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n142 ), .QN(\unit_memory/DRAM/n3020 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][17]  ( .D(
        \unit_memory/DRAM/n1526 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n143 ), .QN(\unit_memory/DRAM/n3021 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][16]  ( .D(
        \unit_memory/DRAM/n1525 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n144 ), .QN(\unit_memory/DRAM/n3022 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][15]  ( .D(
        \unit_memory/DRAM/n1524 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n145 ), .QN(\unit_memory/DRAM/n3023 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][14]  ( .D(
        \unit_memory/DRAM/n1523 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n146 ), .QN(\unit_memory/DRAM/n3024 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][13]  ( .D(
        \unit_memory/DRAM/n1522 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n147 ), .QN(\unit_memory/DRAM/n3025 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][12]  ( .D(
        \unit_memory/DRAM/n1521 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n148 ), .QN(\unit_memory/DRAM/n3026 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][11]  ( .D(
        \unit_memory/DRAM/n1520 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n149 ), .QN(\unit_memory/DRAM/n3027 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][10]  ( .D(
        \unit_memory/DRAM/n1519 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n150 ), .QN(\unit_memory/DRAM/n3028 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][9]  ( .D(\unit_memory/DRAM/n1518 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n151 ), .QN(
        \unit_memory/DRAM/n3029 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][8]  ( .D(\unit_memory/DRAM/n1517 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n152 ), .QN(
        \unit_memory/DRAM/n3030 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][7]  ( .D(\unit_memory/DRAM/n1516 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n153 ), .QN(
        \unit_memory/DRAM/n3031 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][6]  ( .D(\unit_memory/DRAM/n1515 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n154 ), .QN(
        \unit_memory/DRAM/n3032 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][5]  ( .D(\unit_memory/DRAM/n1514 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n155 ), .QN(
        \unit_memory/DRAM/n3033 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][4]  ( .D(\unit_memory/DRAM/n1513 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n156 ), .QN(
        \unit_memory/DRAM/n3034 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][3]  ( .D(\unit_memory/DRAM/n1512 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n157 ), .QN(
        \unit_memory/DRAM/n3035 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][2]  ( .D(\unit_memory/DRAM/n1511 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n158 ), .QN(
        \unit_memory/DRAM/n3036 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][1]  ( .D(\unit_memory/DRAM/n1510 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n159 ), .QN(
        \unit_memory/DRAM/n3037 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[20][0]  ( .D(\unit_memory/DRAM/n1509 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n160 ), .QN(
        \unit_memory/DRAM/n3038 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][23]  ( .D(
        \unit_memory/DRAM/n1660 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n9 ), .QN(\unit_memory/DRAM/n2887 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][22]  ( .D(
        \unit_memory/DRAM/n1659 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n10 ), .QN(\unit_memory/DRAM/n2888 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][21]  ( .D(
        \unit_memory/DRAM/n1658 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n11 ), .QN(\unit_memory/DRAM/n2889 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][20]  ( .D(
        \unit_memory/DRAM/n1657 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n12 ), .QN(\unit_memory/DRAM/n2890 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][19]  ( .D(
        \unit_memory/DRAM/n1656 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n13 ), .QN(\unit_memory/DRAM/n2891 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][18]  ( .D(
        \unit_memory/DRAM/n1655 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n14 ), .QN(\unit_memory/DRAM/n2892 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][17]  ( .D(
        \unit_memory/DRAM/n1654 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n15 ), .QN(\unit_memory/DRAM/n2893 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][16]  ( .D(
        \unit_memory/DRAM/n1653 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n16 ), .QN(\unit_memory/DRAM/n2894 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][15]  ( .D(
        \unit_memory/DRAM/n1652 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n17 ), .QN(\unit_memory/DRAM/n2895 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][14]  ( .D(
        \unit_memory/DRAM/n1651 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n18 ), .QN(\unit_memory/DRAM/n2896 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][13]  ( .D(
        \unit_memory/DRAM/n1650 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n19 ), .QN(\unit_memory/DRAM/n2897 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][12]  ( .D(
        \unit_memory/DRAM/n1649 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n20 ), .QN(\unit_memory/DRAM/n2898 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][11]  ( .D(
        \unit_memory/DRAM/n1648 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n21 ), .QN(\unit_memory/DRAM/n2899 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][10]  ( .D(
        \unit_memory/DRAM/n1647 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n22 ), .QN(\unit_memory/DRAM/n2900 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][9]  ( .D(\unit_memory/DRAM/n1646 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n23 ), .QN(\unit_memory/DRAM/n2901 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][8]  ( .D(\unit_memory/DRAM/n1645 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n24 ), .QN(\unit_memory/DRAM/n2902 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][7]  ( .D(\unit_memory/DRAM/n1644 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n25 ), .QN(\unit_memory/DRAM/n2903 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][6]  ( .D(\unit_memory/DRAM/n1643 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n26 ), .QN(\unit_memory/DRAM/n2904 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][5]  ( .D(\unit_memory/DRAM/n1642 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n27 ), .QN(\unit_memory/DRAM/n2905 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][4]  ( .D(\unit_memory/DRAM/n1641 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n28 ), .QN(\unit_memory/DRAM/n2906 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][3]  ( .D(\unit_memory/DRAM/n1640 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n29 ), .QN(\unit_memory/DRAM/n2907 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][2]  ( .D(\unit_memory/DRAM/n1639 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n30 ), .QN(\unit_memory/DRAM/n2908 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][1]  ( .D(\unit_memory/DRAM/n1638 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n31 ), .QN(\unit_memory/DRAM/n2909 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[16][0]  ( .D(\unit_memory/DRAM/n1637 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n32 ), .QN(\unit_memory/DRAM/n2910 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][23]  ( .D(
        \unit_memory/DRAM/n1788 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2759 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][22]  ( .D(
        \unit_memory/DRAM/n1787 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2760 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][21]  ( .D(
        \unit_memory/DRAM/n1786 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2761 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][20]  ( .D(
        \unit_memory/DRAM/n1785 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2762 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][19]  ( .D(
        \unit_memory/DRAM/n1784 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2763 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][18]  ( .D(
        \unit_memory/DRAM/n1783 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2764 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][17]  ( .D(
        \unit_memory/DRAM/n1782 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2765 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][16]  ( .D(
        \unit_memory/DRAM/n1781 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2766 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][15]  ( .D(
        \unit_memory/DRAM/n1780 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2767 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][14]  ( .D(
        \unit_memory/DRAM/n1779 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2768 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][13]  ( .D(
        \unit_memory/DRAM/n1778 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2769 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][12]  ( .D(
        \unit_memory/DRAM/n1777 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2770 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][11]  ( .D(
        \unit_memory/DRAM/n1776 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2771 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][10]  ( .D(
        \unit_memory/DRAM/n1775 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2772 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][9]  ( .D(\unit_memory/DRAM/n1774 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2773 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][8]  ( .D(\unit_memory/DRAM/n1773 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2774 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][7]  ( .D(\unit_memory/DRAM/n1772 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2775 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][6]  ( .D(\unit_memory/DRAM/n1771 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2776 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][5]  ( .D(\unit_memory/DRAM/n1770 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2777 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][4]  ( .D(\unit_memory/DRAM/n1769 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2778 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][3]  ( .D(\unit_memory/DRAM/n1768 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2779 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][2]  ( .D(\unit_memory/DRAM/n1767 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2780 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][1]  ( .D(\unit_memory/DRAM/n1766 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2781 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[12][0]  ( .D(\unit_memory/DRAM/n1765 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2782 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][23]  ( .D(\unit_memory/DRAM/n1916 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2631 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][22]  ( .D(\unit_memory/DRAM/n1915 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2632 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][21]  ( .D(\unit_memory/DRAM/n1914 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2633 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][20]  ( .D(\unit_memory/DRAM/n1913 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2634 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][19]  ( .D(\unit_memory/DRAM/n1912 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2635 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][18]  ( .D(\unit_memory/DRAM/n1911 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2636 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][17]  ( .D(\unit_memory/DRAM/n1910 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2637 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][16]  ( .D(\unit_memory/DRAM/n1909 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2638 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][15]  ( .D(\unit_memory/DRAM/n1908 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2639 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][14]  ( .D(\unit_memory/DRAM/n1907 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2640 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][13]  ( .D(\unit_memory/DRAM/n1906 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2641 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][12]  ( .D(\unit_memory/DRAM/n1905 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2642 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][11]  ( .D(\unit_memory/DRAM/n1904 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2643 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][10]  ( .D(\unit_memory/DRAM/n1903 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2644 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][9]  ( .D(\unit_memory/DRAM/n1902 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2645 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][8]  ( .D(\unit_memory/DRAM/n1901 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2646 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][7]  ( .D(\unit_memory/DRAM/n1900 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2647 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][6]  ( .D(\unit_memory/DRAM/n1899 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2648 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][5]  ( .D(\unit_memory/DRAM/n1898 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2649 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][4]  ( .D(\unit_memory/DRAM/n1897 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2650 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][3]  ( .D(\unit_memory/DRAM/n1896 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2651 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][2]  ( .D(\unit_memory/DRAM/n1895 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2652 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][1]  ( .D(\unit_memory/DRAM/n1894 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2653 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[8][0]  ( .D(\unit_memory/DRAM/n1893 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2654 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][23]  ( .D(\unit_memory/DRAM/n2044 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2503 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][22]  ( .D(\unit_memory/DRAM/n2043 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2504 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][21]  ( .D(\unit_memory/DRAM/n2042 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2505 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][20]  ( .D(\unit_memory/DRAM/n2041 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2506 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][19]  ( .D(\unit_memory/DRAM/n2040 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2507 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][18]  ( .D(\unit_memory/DRAM/n2039 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2508 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][17]  ( .D(\unit_memory/DRAM/n2038 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2509 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][16]  ( .D(\unit_memory/DRAM/n2037 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2510 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][15]  ( .D(\unit_memory/DRAM/n2036 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2511 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][14]  ( .D(\unit_memory/DRAM/n2035 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2512 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][13]  ( .D(\unit_memory/DRAM/n2034 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2513 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][12]  ( .D(\unit_memory/DRAM/n2033 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2514 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][11]  ( .D(\unit_memory/DRAM/n2032 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2515 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][10]  ( .D(\unit_memory/DRAM/n2031 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2516 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][9]  ( .D(\unit_memory/DRAM/n2030 ), 
        .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2517 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][8]  ( .D(\unit_memory/DRAM/n2029 ), 
        .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2518 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][7]  ( .D(\unit_memory/DRAM/n2028 ), 
        .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2519 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][6]  ( .D(\unit_memory/DRAM/n2027 ), 
        .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2520 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][5]  ( .D(\unit_memory/DRAM/n2026 ), 
        .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2521 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][4]  ( .D(\unit_memory/DRAM/n2025 ), 
        .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2522 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][3]  ( .D(\unit_memory/DRAM/n2024 ), 
        .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2523 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][2]  ( .D(\unit_memory/DRAM/n2023 ), 
        .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2524 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][1]  ( .D(\unit_memory/DRAM/n2022 ), 
        .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2525 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[4][0]  ( .D(\unit_memory/DRAM/n2021 ), 
        .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2526 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][31]  ( .D(
        \unit_memory/DRAM/n1188 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n481 ), .QN(\unit_memory/DRAM/n3359 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][30]  ( .D(
        \unit_memory/DRAM/n1187 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n482 ), .QN(\unit_memory/DRAM/n3360 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][29]  ( .D(
        \unit_memory/DRAM/n1186 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n483 ), .QN(\unit_memory/DRAM/n3361 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][28]  ( .D(
        \unit_memory/DRAM/n1185 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n484 ), .QN(\unit_memory/DRAM/n3362 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][27]  ( .D(
        \unit_memory/DRAM/n1184 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n485 ), .QN(\unit_memory/DRAM/n3363 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][26]  ( .D(
        \unit_memory/DRAM/n1183 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n486 ), .QN(\unit_memory/DRAM/n3364 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][25]  ( .D(
        \unit_memory/DRAM/n1182 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n487 ), .QN(\unit_memory/DRAM/n3365 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][24]  ( .D(
        \unit_memory/DRAM/n1181 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n488 ), .QN(\unit_memory/DRAM/n3366 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][23]  ( .D(
        \unit_memory/DRAM/n1180 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n489 ), .QN(\unit_memory/DRAM/n3367 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][22]  ( .D(
        \unit_memory/DRAM/n1179 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n490 ), .QN(\unit_memory/DRAM/n3368 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][21]  ( .D(
        \unit_memory/DRAM/n1178 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n491 ), .QN(\unit_memory/DRAM/n3369 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][20]  ( .D(
        \unit_memory/DRAM/n1177 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n492 ), .QN(\unit_memory/DRAM/n3370 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][19]  ( .D(
        \unit_memory/DRAM/n1176 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n493 ), .QN(\unit_memory/DRAM/n3371 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][18]  ( .D(
        \unit_memory/DRAM/n1175 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n494 ), .QN(\unit_memory/DRAM/n3372 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][17]  ( .D(
        \unit_memory/DRAM/n1174 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n495 ), .QN(\unit_memory/DRAM/n3373 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][16]  ( .D(
        \unit_memory/DRAM/n1173 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n496 ), .QN(\unit_memory/DRAM/n3374 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][15]  ( .D(
        \unit_memory/DRAM/n1172 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n497 ), .QN(\unit_memory/DRAM/n3375 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][14]  ( .D(
        \unit_memory/DRAM/n1171 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n498 ), .QN(\unit_memory/DRAM/n3376 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][13]  ( .D(
        \unit_memory/DRAM/n1170 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n499 ), .QN(\unit_memory/DRAM/n3377 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][12]  ( .D(
        \unit_memory/DRAM/n1169 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n500 ), .QN(\unit_memory/DRAM/n3378 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][11]  ( .D(
        \unit_memory/DRAM/n1168 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n501 ), .QN(\unit_memory/DRAM/n3379 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][10]  ( .D(
        \unit_memory/DRAM/n1167 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n502 ), .QN(\unit_memory/DRAM/n3380 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][9]  ( .D(\unit_memory/DRAM/n1166 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n503 ), .QN(
        \unit_memory/DRAM/n3381 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[31][8]  ( .D(\unit_memory/DRAM/n1165 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n504 ), .QN(
        \unit_memory/DRAM/n3382 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][31]  ( .D(\unit_memory/DRAM/n2180 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2367 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][30]  ( .D(\unit_memory/DRAM/n2179 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2368 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][29]  ( .D(\unit_memory/DRAM/n2178 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2369 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][28]  ( .D(\unit_memory/DRAM/n2177 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2370 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][27]  ( .D(\unit_memory/DRAM/n2176 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2371 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][26]  ( .D(\unit_memory/DRAM/n2175 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2372 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][25]  ( .D(\unit_memory/DRAM/n2174 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2373 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][24]  ( .D(\unit_memory/DRAM/n2173 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2374 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][31]  ( .D(
        \unit_memory/DRAM/n1220 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n449 ), .QN(\unit_memory/DRAM/n3327 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][30]  ( .D(
        \unit_memory/DRAM/n1219 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n450 ), .QN(\unit_memory/DRAM/n3328 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][29]  ( .D(
        \unit_memory/DRAM/n1218 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n451 ), .QN(\unit_memory/DRAM/n3329 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][28]  ( .D(
        \unit_memory/DRAM/n1217 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n452 ), .QN(\unit_memory/DRAM/n3330 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][27]  ( .D(
        \unit_memory/DRAM/n1216 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n453 ), .QN(\unit_memory/DRAM/n3331 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][26]  ( .D(
        \unit_memory/DRAM/n1215 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n454 ), .QN(\unit_memory/DRAM/n3332 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][25]  ( .D(
        \unit_memory/DRAM/n1214 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n455 ), .QN(\unit_memory/DRAM/n3333 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][24]  ( .D(
        \unit_memory/DRAM/n1213 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n456 ), .QN(\unit_memory/DRAM/n3334 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][31]  ( .D(
        \unit_memory/DRAM/n1348 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n321 ), .QN(\unit_memory/DRAM/n3199 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][30]  ( .D(
        \unit_memory/DRAM/n1347 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n322 ), .QN(\unit_memory/DRAM/n3200 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][29]  ( .D(
        \unit_memory/DRAM/n1346 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n323 ), .QN(\unit_memory/DRAM/n3201 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][28]  ( .D(
        \unit_memory/DRAM/n1345 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n324 ), .QN(\unit_memory/DRAM/n3202 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][27]  ( .D(
        \unit_memory/DRAM/n1344 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n325 ), .QN(\unit_memory/DRAM/n3203 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][26]  ( .D(
        \unit_memory/DRAM/n1343 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n326 ), .QN(\unit_memory/DRAM/n3204 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][25]  ( .D(
        \unit_memory/DRAM/n1342 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n327 ), .QN(\unit_memory/DRAM/n3205 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][24]  ( .D(
        \unit_memory/DRAM/n1341 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n328 ), .QN(\unit_memory/DRAM/n3206 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][31]  ( .D(
        \unit_memory/DRAM/n1476 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n193 ), .QN(\unit_memory/DRAM/n3071 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][30]  ( .D(
        \unit_memory/DRAM/n1475 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n194 ), .QN(\unit_memory/DRAM/n3072 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][29]  ( .D(
        \unit_memory/DRAM/n1474 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n195 ), .QN(\unit_memory/DRAM/n3073 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][28]  ( .D(
        \unit_memory/DRAM/n1473 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n196 ), .QN(\unit_memory/DRAM/n3074 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][27]  ( .D(
        \unit_memory/DRAM/n1472 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n197 ), .QN(\unit_memory/DRAM/n3075 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][26]  ( .D(
        \unit_memory/DRAM/n1471 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n198 ), .QN(\unit_memory/DRAM/n3076 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][25]  ( .D(
        \unit_memory/DRAM/n1470 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n199 ), .QN(\unit_memory/DRAM/n3077 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][24]  ( .D(
        \unit_memory/DRAM/n1469 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n200 ), .QN(\unit_memory/DRAM/n3078 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][31]  ( .D(
        \unit_memory/DRAM/n1604 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n65 ), .QN(\unit_memory/DRAM/n2943 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][30]  ( .D(
        \unit_memory/DRAM/n1603 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n66 ), .QN(\unit_memory/DRAM/n2944 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][29]  ( .D(
        \unit_memory/DRAM/n1602 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n67 ), .QN(\unit_memory/DRAM/n2945 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][28]  ( .D(
        \unit_memory/DRAM/n1601 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n68 ), .QN(\unit_memory/DRAM/n2946 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][27]  ( .D(
        \unit_memory/DRAM/n1600 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n69 ), .QN(\unit_memory/DRAM/n2947 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][26]  ( .D(
        \unit_memory/DRAM/n1599 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n70 ), .QN(\unit_memory/DRAM/n2948 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][25]  ( .D(
        \unit_memory/DRAM/n1598 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n71 ), .QN(\unit_memory/DRAM/n2949 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][24]  ( .D(
        \unit_memory/DRAM/n1597 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n72 ), .QN(\unit_memory/DRAM/n2950 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][31]  ( .D(
        \unit_memory/DRAM/n1732 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2815 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][30]  ( .D(
        \unit_memory/DRAM/n1731 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2816 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][29]  ( .D(
        \unit_memory/DRAM/n1730 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2817 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][28]  ( .D(
        \unit_memory/DRAM/n1729 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2818 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][27]  ( .D(
        \unit_memory/DRAM/n1728 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2819 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][26]  ( .D(
        \unit_memory/DRAM/n1727 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2820 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][25]  ( .D(
        \unit_memory/DRAM/n1726 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2821 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][24]  ( .D(
        \unit_memory/DRAM/n1725 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2822 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][31]  ( .D(
        \unit_memory/DRAM/n1860 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2687 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][30]  ( .D(
        \unit_memory/DRAM/n1859 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2688 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][29]  ( .D(
        \unit_memory/DRAM/n1858 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2689 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][28]  ( .D(
        \unit_memory/DRAM/n1857 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2690 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][27]  ( .D(
        \unit_memory/DRAM/n1856 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2691 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][26]  ( .D(
        \unit_memory/DRAM/n1855 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2692 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][25]  ( .D(
        \unit_memory/DRAM/n1854 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2693 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][24]  ( .D(
        \unit_memory/DRAM/n1853 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2694 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][31]  ( .D(\unit_memory/DRAM/n1988 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2559 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][30]  ( .D(\unit_memory/DRAM/n1987 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2560 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][29]  ( .D(\unit_memory/DRAM/n1986 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2561 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][28]  ( .D(\unit_memory/DRAM/n1985 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2562 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][27]  ( .D(\unit_memory/DRAM/n1984 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2563 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][26]  ( .D(\unit_memory/DRAM/n1983 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2564 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][25]  ( .D(\unit_memory/DRAM/n1982 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2565 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][24]  ( .D(\unit_memory/DRAM/n1981 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2566 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][31]  ( .D(\unit_memory/DRAM/n2116 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2431 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][30]  ( .D(\unit_memory/DRAM/n2115 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2432 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][29]  ( .D(\unit_memory/DRAM/n2114 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2433 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][28]  ( .D(\unit_memory/DRAM/n2113 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2434 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][27]  ( .D(\unit_memory/DRAM/n2112 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2435 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][26]  ( .D(\unit_memory/DRAM/n2111 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2436 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][25]  ( .D(\unit_memory/DRAM/n2110 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2437 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][24]  ( .D(\unit_memory/DRAM/n2109 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2438 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][31]  ( .D(
        \unit_memory/DRAM/n1252 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n417 ), .QN(\unit_memory/DRAM/n3295 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][30]  ( .D(
        \unit_memory/DRAM/n1251 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n418 ), .QN(\unit_memory/DRAM/n3296 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][29]  ( .D(
        \unit_memory/DRAM/n1250 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n419 ), .QN(\unit_memory/DRAM/n3297 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][28]  ( .D(
        \unit_memory/DRAM/n1249 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n420 ), .QN(\unit_memory/DRAM/n3298 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][27]  ( .D(
        \unit_memory/DRAM/n1248 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n421 ), .QN(\unit_memory/DRAM/n3299 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][26]  ( .D(
        \unit_memory/DRAM/n1247 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n422 ), .QN(\unit_memory/DRAM/n3300 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][25]  ( .D(
        \unit_memory/DRAM/n1246 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n423 ), .QN(\unit_memory/DRAM/n3301 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][24]  ( .D(
        \unit_memory/DRAM/n1245 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n424 ), .QN(\unit_memory/DRAM/n3302 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][31]  ( .D(
        \unit_memory/DRAM/n1380 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n289 ), .QN(\unit_memory/DRAM/n3167 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][30]  ( .D(
        \unit_memory/DRAM/n1379 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n290 ), .QN(\unit_memory/DRAM/n3168 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][29]  ( .D(
        \unit_memory/DRAM/n1378 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n291 ), .QN(\unit_memory/DRAM/n3169 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][28]  ( .D(
        \unit_memory/DRAM/n1377 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n292 ), .QN(\unit_memory/DRAM/n3170 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][27]  ( .D(
        \unit_memory/DRAM/n1376 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n293 ), .QN(\unit_memory/DRAM/n3171 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][26]  ( .D(
        \unit_memory/DRAM/n1375 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n294 ), .QN(\unit_memory/DRAM/n3172 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][25]  ( .D(
        \unit_memory/DRAM/n1374 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n295 ), .QN(\unit_memory/DRAM/n3173 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][24]  ( .D(
        \unit_memory/DRAM/n1373 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n296 ), .QN(\unit_memory/DRAM/n3174 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][31]  ( .D(
        \unit_memory/DRAM/n1508 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n161 ), .QN(\unit_memory/DRAM/n3039 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][30]  ( .D(
        \unit_memory/DRAM/n1507 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n162 ), .QN(\unit_memory/DRAM/n3040 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][29]  ( .D(
        \unit_memory/DRAM/n1506 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n163 ), .QN(\unit_memory/DRAM/n3041 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][28]  ( .D(
        \unit_memory/DRAM/n1505 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n164 ), .QN(\unit_memory/DRAM/n3042 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][27]  ( .D(
        \unit_memory/DRAM/n1504 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n165 ), .QN(\unit_memory/DRAM/n3043 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][26]  ( .D(
        \unit_memory/DRAM/n1503 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n166 ), .QN(\unit_memory/DRAM/n3044 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][25]  ( .D(
        \unit_memory/DRAM/n1502 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n167 ), .QN(\unit_memory/DRAM/n3045 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][24]  ( .D(
        \unit_memory/DRAM/n1501 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n168 ), .QN(\unit_memory/DRAM/n3046 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][31]  ( .D(
        \unit_memory/DRAM/n1636 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n33 ), .QN(\unit_memory/DRAM/n2911 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][30]  ( .D(
        \unit_memory/DRAM/n1635 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n34 ), .QN(\unit_memory/DRAM/n2912 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][29]  ( .D(
        \unit_memory/DRAM/n1634 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n35 ), .QN(\unit_memory/DRAM/n2913 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][28]  ( .D(
        \unit_memory/DRAM/n1633 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n36 ), .QN(\unit_memory/DRAM/n2914 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][27]  ( .D(
        \unit_memory/DRAM/n1632 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n37 ), .QN(\unit_memory/DRAM/n2915 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][26]  ( .D(
        \unit_memory/DRAM/n1631 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n38 ), .QN(\unit_memory/DRAM/n2916 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][25]  ( .D(
        \unit_memory/DRAM/n1630 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n39 ), .QN(\unit_memory/DRAM/n2917 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][24]  ( .D(
        \unit_memory/DRAM/n1629 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n40 ), .QN(\unit_memory/DRAM/n2918 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][31]  ( .D(
        \unit_memory/DRAM/n1764 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2783 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][30]  ( .D(
        \unit_memory/DRAM/n1763 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2784 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][29]  ( .D(
        \unit_memory/DRAM/n1762 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2785 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][28]  ( .D(
        \unit_memory/DRAM/n1761 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2786 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][27]  ( .D(
        \unit_memory/DRAM/n1760 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2787 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][26]  ( .D(
        \unit_memory/DRAM/n1759 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2788 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][25]  ( .D(
        \unit_memory/DRAM/n1758 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2789 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][24]  ( .D(
        \unit_memory/DRAM/n1757 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2790 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][31]  ( .D(\unit_memory/DRAM/n1892 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2655 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][30]  ( .D(\unit_memory/DRAM/n1891 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2656 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][29]  ( .D(\unit_memory/DRAM/n1890 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2657 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][28]  ( .D(\unit_memory/DRAM/n1889 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2658 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][27]  ( .D(\unit_memory/DRAM/n1888 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2659 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][26]  ( .D(\unit_memory/DRAM/n1887 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2660 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][25]  ( .D(\unit_memory/DRAM/n1886 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2661 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][24]  ( .D(\unit_memory/DRAM/n1885 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2662 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][31]  ( .D(\unit_memory/DRAM/n2020 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2527 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][30]  ( .D(\unit_memory/DRAM/n2019 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2528 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][29]  ( .D(\unit_memory/DRAM/n2018 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2529 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][28]  ( .D(\unit_memory/DRAM/n2017 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2530 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][27]  ( .D(\unit_memory/DRAM/n2016 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2531 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][26]  ( .D(\unit_memory/DRAM/n2015 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2532 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][25]  ( .D(\unit_memory/DRAM/n2014 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2533 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][24]  ( .D(\unit_memory/DRAM/n2013 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2534 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][31]  ( .D(\unit_memory/DRAM/n2148 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2399 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][30]  ( .D(\unit_memory/DRAM/n2147 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2400 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][29]  ( .D(\unit_memory/DRAM/n2146 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2401 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][28]  ( .D(\unit_memory/DRAM/n2145 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2402 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][27]  ( .D(\unit_memory/DRAM/n2144 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2403 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][26]  ( .D(\unit_memory/DRAM/n2143 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2404 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][25]  ( .D(\unit_memory/DRAM/n2142 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2405 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][24]  ( .D(\unit_memory/DRAM/n2141 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2406 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][23]  ( .D(
        \unit_memory/DRAM/n1212 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n457 ), .QN(\unit_memory/DRAM/n3335 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][22]  ( .D(
        \unit_memory/DRAM/n1211 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n458 ), .QN(\unit_memory/DRAM/n3336 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][21]  ( .D(
        \unit_memory/DRAM/n1210 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n459 ), .QN(\unit_memory/DRAM/n3337 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][20]  ( .D(
        \unit_memory/DRAM/n1209 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n460 ), .QN(\unit_memory/DRAM/n3338 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][19]  ( .D(
        \unit_memory/DRAM/n1208 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n461 ), .QN(\unit_memory/DRAM/n3339 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][18]  ( .D(
        \unit_memory/DRAM/n1207 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n462 ), .QN(\unit_memory/DRAM/n3340 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][17]  ( .D(
        \unit_memory/DRAM/n1206 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n463 ), .QN(\unit_memory/DRAM/n3341 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][16]  ( .D(
        \unit_memory/DRAM/n1205 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n464 ), .QN(\unit_memory/DRAM/n3342 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][15]  ( .D(
        \unit_memory/DRAM/n1204 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n465 ), .QN(\unit_memory/DRAM/n3343 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][14]  ( .D(
        \unit_memory/DRAM/n1203 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n466 ), .QN(\unit_memory/DRAM/n3344 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][13]  ( .D(
        \unit_memory/DRAM/n1202 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n467 ), .QN(\unit_memory/DRAM/n3345 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][12]  ( .D(
        \unit_memory/DRAM/n1201 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n468 ), .QN(\unit_memory/DRAM/n3346 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][11]  ( .D(
        \unit_memory/DRAM/n1200 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n469 ), .QN(\unit_memory/DRAM/n3347 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][10]  ( .D(
        \unit_memory/DRAM/n1199 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n470 ), .QN(\unit_memory/DRAM/n3348 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][9]  ( .D(\unit_memory/DRAM/n1198 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n471 ), .QN(
        \unit_memory/DRAM/n3349 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][8]  ( .D(\unit_memory/DRAM/n1197 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n472 ), .QN(
        \unit_memory/DRAM/n3350 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][7]  ( .D(\unit_memory/DRAM/n1196 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n473 ), .QN(
        \unit_memory/DRAM/n3351 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][6]  ( .D(\unit_memory/DRAM/n1195 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n474 ), .QN(
        \unit_memory/DRAM/n3352 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][5]  ( .D(\unit_memory/DRAM/n1194 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n475 ), .QN(
        \unit_memory/DRAM/n3353 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][4]  ( .D(\unit_memory/DRAM/n1193 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n476 ), .QN(
        \unit_memory/DRAM/n3354 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][3]  ( .D(\unit_memory/DRAM/n1192 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n477 ), .QN(
        \unit_memory/DRAM/n3355 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][2]  ( .D(\unit_memory/DRAM/n1191 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n478 ), .QN(
        \unit_memory/DRAM/n3356 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][1]  ( .D(\unit_memory/DRAM/n1190 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n479 ), .QN(
        \unit_memory/DRAM/n3357 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[30][0]  ( .D(\unit_memory/DRAM/n1189 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n480 ), .QN(
        \unit_memory/DRAM/n3358 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][23]  ( .D(
        \unit_memory/DRAM/n1340 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n329 ), .QN(\unit_memory/DRAM/n3207 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][22]  ( .D(
        \unit_memory/DRAM/n1339 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n330 ), .QN(\unit_memory/DRAM/n3208 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][21]  ( .D(
        \unit_memory/DRAM/n1338 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n331 ), .QN(\unit_memory/DRAM/n3209 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][20]  ( .D(
        \unit_memory/DRAM/n1337 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n332 ), .QN(\unit_memory/DRAM/n3210 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][19]  ( .D(
        \unit_memory/DRAM/n1336 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n333 ), .QN(\unit_memory/DRAM/n3211 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][18]  ( .D(
        \unit_memory/DRAM/n1335 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n334 ), .QN(\unit_memory/DRAM/n3212 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][17]  ( .D(
        \unit_memory/DRAM/n1334 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n335 ), .QN(\unit_memory/DRAM/n3213 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][16]  ( .D(
        \unit_memory/DRAM/n1333 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n336 ), .QN(\unit_memory/DRAM/n3214 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][15]  ( .D(
        \unit_memory/DRAM/n1332 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n337 ), .QN(\unit_memory/DRAM/n3215 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][14]  ( .D(
        \unit_memory/DRAM/n1331 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n338 ), .QN(\unit_memory/DRAM/n3216 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][13]  ( .D(
        \unit_memory/DRAM/n1330 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n339 ), .QN(\unit_memory/DRAM/n3217 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][12]  ( .D(
        \unit_memory/DRAM/n1329 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n340 ), .QN(\unit_memory/DRAM/n3218 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][11]  ( .D(
        \unit_memory/DRAM/n1328 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n341 ), .QN(\unit_memory/DRAM/n3219 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][10]  ( .D(
        \unit_memory/DRAM/n1327 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n342 ), .QN(\unit_memory/DRAM/n3220 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][9]  ( .D(\unit_memory/DRAM/n1326 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n343 ), .QN(
        \unit_memory/DRAM/n3221 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][8]  ( .D(\unit_memory/DRAM/n1325 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n344 ), .QN(
        \unit_memory/DRAM/n3222 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][7]  ( .D(\unit_memory/DRAM/n1324 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n345 ), .QN(
        \unit_memory/DRAM/n3223 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][6]  ( .D(\unit_memory/DRAM/n1323 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n346 ), .QN(
        \unit_memory/DRAM/n3224 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][5]  ( .D(\unit_memory/DRAM/n1322 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n347 ), .QN(
        \unit_memory/DRAM/n3225 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][4]  ( .D(\unit_memory/DRAM/n1321 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n348 ), .QN(
        \unit_memory/DRAM/n3226 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][3]  ( .D(\unit_memory/DRAM/n1320 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n349 ), .QN(
        \unit_memory/DRAM/n3227 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][2]  ( .D(\unit_memory/DRAM/n1319 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n350 ), .QN(
        \unit_memory/DRAM/n3228 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][1]  ( .D(\unit_memory/DRAM/n1318 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n351 ), .QN(
        \unit_memory/DRAM/n3229 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[26][0]  ( .D(\unit_memory/DRAM/n1317 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n352 ), .QN(
        \unit_memory/DRAM/n3230 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][23]  ( .D(
        \unit_memory/DRAM/n1468 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n201 ), .QN(\unit_memory/DRAM/n3079 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][22]  ( .D(
        \unit_memory/DRAM/n1467 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n202 ), .QN(\unit_memory/DRAM/n3080 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][21]  ( .D(
        \unit_memory/DRAM/n1466 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n203 ), .QN(\unit_memory/DRAM/n3081 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][20]  ( .D(
        \unit_memory/DRAM/n1465 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n204 ), .QN(\unit_memory/DRAM/n3082 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][19]  ( .D(
        \unit_memory/DRAM/n1464 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n205 ), .QN(\unit_memory/DRAM/n3083 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][18]  ( .D(
        \unit_memory/DRAM/n1463 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n206 ), .QN(\unit_memory/DRAM/n3084 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][17]  ( .D(
        \unit_memory/DRAM/n1462 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n207 ), .QN(\unit_memory/DRAM/n3085 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][16]  ( .D(
        \unit_memory/DRAM/n1461 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n208 ), .QN(\unit_memory/DRAM/n3086 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][15]  ( .D(
        \unit_memory/DRAM/n1460 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n209 ), .QN(\unit_memory/DRAM/n3087 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][14]  ( .D(
        \unit_memory/DRAM/n1459 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n210 ), .QN(\unit_memory/DRAM/n3088 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][13]  ( .D(
        \unit_memory/DRAM/n1458 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n211 ), .QN(\unit_memory/DRAM/n3089 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][12]  ( .D(
        \unit_memory/DRAM/n1457 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n212 ), .QN(\unit_memory/DRAM/n3090 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][11]  ( .D(
        \unit_memory/DRAM/n1456 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n213 ), .QN(\unit_memory/DRAM/n3091 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][10]  ( .D(
        \unit_memory/DRAM/n1455 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n214 ), .QN(\unit_memory/DRAM/n3092 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][9]  ( .D(\unit_memory/DRAM/n1454 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n215 ), .QN(
        \unit_memory/DRAM/n3093 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][8]  ( .D(\unit_memory/DRAM/n1453 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n216 ), .QN(
        \unit_memory/DRAM/n3094 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][7]  ( .D(\unit_memory/DRAM/n1452 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n217 ), .QN(
        \unit_memory/DRAM/n3095 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][6]  ( .D(\unit_memory/DRAM/n1451 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n218 ), .QN(
        \unit_memory/DRAM/n3096 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][5]  ( .D(\unit_memory/DRAM/n1450 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n219 ), .QN(
        \unit_memory/DRAM/n3097 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][4]  ( .D(\unit_memory/DRAM/n1449 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n220 ), .QN(
        \unit_memory/DRAM/n3098 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][3]  ( .D(\unit_memory/DRAM/n1448 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n221 ), .QN(
        \unit_memory/DRAM/n3099 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][2]  ( .D(\unit_memory/DRAM/n1447 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n222 ), .QN(
        \unit_memory/DRAM/n3100 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][1]  ( .D(\unit_memory/DRAM/n1446 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n223 ), .QN(
        \unit_memory/DRAM/n3101 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[22][0]  ( .D(\unit_memory/DRAM/n1445 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n224 ), .QN(
        \unit_memory/DRAM/n3102 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][23]  ( .D(
        \unit_memory/DRAM/n1596 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n73 ), .QN(\unit_memory/DRAM/n2951 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][22]  ( .D(
        \unit_memory/DRAM/n1595 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n74 ), .QN(\unit_memory/DRAM/n2952 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][21]  ( .D(
        \unit_memory/DRAM/n1594 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n75 ), .QN(\unit_memory/DRAM/n2953 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][20]  ( .D(
        \unit_memory/DRAM/n1593 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n76 ), .QN(\unit_memory/DRAM/n2954 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][19]  ( .D(
        \unit_memory/DRAM/n1592 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n77 ), .QN(\unit_memory/DRAM/n2955 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][18]  ( .D(
        \unit_memory/DRAM/n1591 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n78 ), .QN(\unit_memory/DRAM/n2956 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][17]  ( .D(
        \unit_memory/DRAM/n1590 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n79 ), .QN(\unit_memory/DRAM/n2957 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][16]  ( .D(
        \unit_memory/DRAM/n1589 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n80 ), .QN(\unit_memory/DRAM/n2958 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][15]  ( .D(
        \unit_memory/DRAM/n1588 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n81 ), .QN(\unit_memory/DRAM/n2959 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][14]  ( .D(
        \unit_memory/DRAM/n1587 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n82 ), .QN(\unit_memory/DRAM/n2960 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][13]  ( .D(
        \unit_memory/DRAM/n1586 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n83 ), .QN(\unit_memory/DRAM/n2961 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][12]  ( .D(
        \unit_memory/DRAM/n1585 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n84 ), .QN(\unit_memory/DRAM/n2962 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][11]  ( .D(
        \unit_memory/DRAM/n1584 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n85 ), .QN(\unit_memory/DRAM/n2963 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][10]  ( .D(
        \unit_memory/DRAM/n1583 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n86 ), .QN(\unit_memory/DRAM/n2964 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][9]  ( .D(\unit_memory/DRAM/n1582 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n87 ), .QN(\unit_memory/DRAM/n2965 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][8]  ( .D(\unit_memory/DRAM/n1581 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n88 ), .QN(\unit_memory/DRAM/n2966 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][7]  ( .D(\unit_memory/DRAM/n1580 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n89 ), .QN(\unit_memory/DRAM/n2967 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][6]  ( .D(\unit_memory/DRAM/n1579 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n90 ), .QN(\unit_memory/DRAM/n2968 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][5]  ( .D(\unit_memory/DRAM/n1578 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n91 ), .QN(\unit_memory/DRAM/n2969 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][4]  ( .D(\unit_memory/DRAM/n1577 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n92 ), .QN(\unit_memory/DRAM/n2970 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][3]  ( .D(\unit_memory/DRAM/n1576 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n93 ), .QN(\unit_memory/DRAM/n2971 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][2]  ( .D(\unit_memory/DRAM/n1575 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n94 ), .QN(\unit_memory/DRAM/n2972 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][1]  ( .D(\unit_memory/DRAM/n1574 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n95 ), .QN(\unit_memory/DRAM/n2973 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[18][0]  ( .D(\unit_memory/DRAM/n1573 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n96 ), .QN(\unit_memory/DRAM/n2974 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][23]  ( .D(
        \unit_memory/DRAM/n1724 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2823 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][22]  ( .D(
        \unit_memory/DRAM/n1723 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2824 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][21]  ( .D(
        \unit_memory/DRAM/n1722 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2825 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][20]  ( .D(
        \unit_memory/DRAM/n1721 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2826 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][19]  ( .D(
        \unit_memory/DRAM/n1720 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2827 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][18]  ( .D(
        \unit_memory/DRAM/n1719 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2828 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][17]  ( .D(
        \unit_memory/DRAM/n1718 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2829 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][16]  ( .D(
        \unit_memory/DRAM/n1717 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2830 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][15]  ( .D(
        \unit_memory/DRAM/n1716 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2831 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][14]  ( .D(
        \unit_memory/DRAM/n1715 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2832 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][13]  ( .D(
        \unit_memory/DRAM/n1714 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2833 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][12]  ( .D(
        \unit_memory/DRAM/n1713 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2834 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][11]  ( .D(
        \unit_memory/DRAM/n1712 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2835 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][10]  ( .D(
        \unit_memory/DRAM/n1711 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2836 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][9]  ( .D(\unit_memory/DRAM/n1710 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2837 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][8]  ( .D(\unit_memory/DRAM/n1709 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2838 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][7]  ( .D(\unit_memory/DRAM/n1708 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2839 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][6]  ( .D(\unit_memory/DRAM/n1707 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2840 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][5]  ( .D(\unit_memory/DRAM/n1706 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2841 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][4]  ( .D(\unit_memory/DRAM/n1705 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2842 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][3]  ( .D(\unit_memory/DRAM/n1704 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2843 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][2]  ( .D(\unit_memory/DRAM/n1703 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2844 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][1]  ( .D(\unit_memory/DRAM/n1702 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2845 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[14][0]  ( .D(\unit_memory/DRAM/n1701 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2846 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][23]  ( .D(
        \unit_memory/DRAM/n1852 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2695 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][22]  ( .D(
        \unit_memory/DRAM/n1851 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2696 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][21]  ( .D(
        \unit_memory/DRAM/n1850 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2697 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][20]  ( .D(
        \unit_memory/DRAM/n1849 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2698 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][19]  ( .D(
        \unit_memory/DRAM/n1848 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2699 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][18]  ( .D(
        \unit_memory/DRAM/n1847 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2700 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][17]  ( .D(
        \unit_memory/DRAM/n1846 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2701 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][16]  ( .D(
        \unit_memory/DRAM/n1845 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2702 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][15]  ( .D(
        \unit_memory/DRAM/n1844 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2703 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][14]  ( .D(
        \unit_memory/DRAM/n1843 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2704 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][13]  ( .D(
        \unit_memory/DRAM/n1842 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2705 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][12]  ( .D(
        \unit_memory/DRAM/n1841 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2706 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][11]  ( .D(
        \unit_memory/DRAM/n1840 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2707 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][10]  ( .D(
        \unit_memory/DRAM/n1839 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2708 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][9]  ( .D(\unit_memory/DRAM/n1838 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2709 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][8]  ( .D(\unit_memory/DRAM/n1837 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2710 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][7]  ( .D(\unit_memory/DRAM/n1836 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2711 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][6]  ( .D(\unit_memory/DRAM/n1835 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2712 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][5]  ( .D(\unit_memory/DRAM/n1834 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2713 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][4]  ( .D(\unit_memory/DRAM/n1833 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2714 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][3]  ( .D(\unit_memory/DRAM/n1832 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2715 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][2]  ( .D(\unit_memory/DRAM/n1831 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2716 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][1]  ( .D(\unit_memory/DRAM/n1830 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2717 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[10][0]  ( .D(\unit_memory/DRAM/n1829 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2718 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][23]  ( .D(\unit_memory/DRAM/n1980 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2567 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][22]  ( .D(\unit_memory/DRAM/n1979 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2568 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][21]  ( .D(\unit_memory/DRAM/n1978 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2569 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][20]  ( .D(\unit_memory/DRAM/n1977 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2570 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][19]  ( .D(\unit_memory/DRAM/n1976 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2571 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][18]  ( .D(\unit_memory/DRAM/n1975 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2572 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][17]  ( .D(\unit_memory/DRAM/n1974 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2573 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][16]  ( .D(\unit_memory/DRAM/n1973 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2574 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][15]  ( .D(\unit_memory/DRAM/n1972 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2575 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][14]  ( .D(\unit_memory/DRAM/n1971 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2576 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][13]  ( .D(\unit_memory/DRAM/n1970 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2577 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][12]  ( .D(\unit_memory/DRAM/n1969 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2578 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][11]  ( .D(\unit_memory/DRAM/n1968 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2579 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][10]  ( .D(\unit_memory/DRAM/n1967 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2580 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][9]  ( .D(\unit_memory/DRAM/n1966 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2581 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][8]  ( .D(\unit_memory/DRAM/n1965 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2582 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][7]  ( .D(\unit_memory/DRAM/n1964 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2583 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][6]  ( .D(\unit_memory/DRAM/n1963 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2584 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][5]  ( .D(\unit_memory/DRAM/n1962 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2585 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][4]  ( .D(\unit_memory/DRAM/n1961 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2586 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][3]  ( .D(\unit_memory/DRAM/n1960 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2587 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][2]  ( .D(\unit_memory/DRAM/n1959 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2588 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][1]  ( .D(\unit_memory/DRAM/n1958 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2589 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[6][0]  ( .D(\unit_memory/DRAM/n1957 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2590 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][23]  ( .D(\unit_memory/DRAM/n2108 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2439 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][22]  ( .D(\unit_memory/DRAM/n2107 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2440 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][21]  ( .D(\unit_memory/DRAM/n2106 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2441 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][20]  ( .D(\unit_memory/DRAM/n2105 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2442 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][19]  ( .D(\unit_memory/DRAM/n2104 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2443 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][18]  ( .D(\unit_memory/DRAM/n2103 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2444 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][17]  ( .D(\unit_memory/DRAM/n2102 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2445 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][16]  ( .D(\unit_memory/DRAM/n2101 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2446 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][15]  ( .D(\unit_memory/DRAM/n2100 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2447 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][14]  ( .D(\unit_memory/DRAM/n2099 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2448 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][13]  ( .D(\unit_memory/DRAM/n2098 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2449 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][12]  ( .D(\unit_memory/DRAM/n2097 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2450 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][11]  ( .D(\unit_memory/DRAM/n2096 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2451 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][10]  ( .D(\unit_memory/DRAM/n2095 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2452 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][9]  ( .D(\unit_memory/DRAM/n2094 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2453 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][8]  ( .D(\unit_memory/DRAM/n2093 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2454 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][7]  ( .D(\unit_memory/DRAM/n2092 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2455 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][6]  ( .D(\unit_memory/DRAM/n2091 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2456 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][5]  ( .D(\unit_memory/DRAM/n2090 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2457 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][4]  ( .D(\unit_memory/DRAM/n2089 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2458 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][3]  ( .D(\unit_memory/DRAM/n2088 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2459 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][2]  ( .D(\unit_memory/DRAM/n2087 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2460 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][1]  ( .D(\unit_memory/DRAM/n2086 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2461 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[2][0]  ( .D(\unit_memory/DRAM/n2085 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2462 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][7]  ( .D(\unit_memory/DRAM/n2156 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2391 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][6]  ( .D(\unit_memory/DRAM/n2155 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2392 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][5]  ( .D(\unit_memory/DRAM/n2154 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2393 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][4]  ( .D(\unit_memory/DRAM/n2153 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2394 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][3]  ( .D(\unit_memory/DRAM/n2152 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2395 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][2]  ( .D(\unit_memory/DRAM/n2151 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2396 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][1]  ( .D(\unit_memory/DRAM/n2150 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2397 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][23]  ( .D(\unit_memory/DRAM/n2172 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2375 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][22]  ( .D(\unit_memory/DRAM/n2171 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2376 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][21]  ( .D(\unit_memory/DRAM/n2170 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2377 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][20]  ( .D(\unit_memory/DRAM/n2169 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2378 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][19]  ( .D(\unit_memory/DRAM/n2168 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2379 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][18]  ( .D(\unit_memory/DRAM/n2167 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2380 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][17]  ( .D(\unit_memory/DRAM/n2166 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2381 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][16]  ( .D(\unit_memory/DRAM/n2165 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2382 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][15]  ( .D(\unit_memory/DRAM/n2164 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2383 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][14]  ( .D(\unit_memory/DRAM/n2163 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2384 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][13]  ( .D(\unit_memory/DRAM/n2162 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2385 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][12]  ( .D(\unit_memory/DRAM/n2161 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2386 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][11]  ( .D(\unit_memory/DRAM/n2160 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2387 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][10]  ( .D(\unit_memory/DRAM/n2159 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2388 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][9]  ( .D(\unit_memory/DRAM/n2158 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2389 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][8]  ( .D(\unit_memory/DRAM/n2157 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2390 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[0][0]  ( .D(\unit_memory/DRAM/n2149 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2398 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][23]  ( .D(
        \unit_memory/DRAM/n1244 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n425 ), .QN(\unit_memory/DRAM/n3303 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][22]  ( .D(
        \unit_memory/DRAM/n1243 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n426 ), .QN(\unit_memory/DRAM/n3304 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][21]  ( .D(
        \unit_memory/DRAM/n1242 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n427 ), .QN(\unit_memory/DRAM/n3305 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][20]  ( .D(
        \unit_memory/DRAM/n1241 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n428 ), .QN(\unit_memory/DRAM/n3306 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][19]  ( .D(
        \unit_memory/DRAM/n1240 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n429 ), .QN(\unit_memory/DRAM/n3307 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][18]  ( .D(
        \unit_memory/DRAM/n1239 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n430 ), .QN(\unit_memory/DRAM/n3308 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][17]  ( .D(
        \unit_memory/DRAM/n1238 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n431 ), .QN(\unit_memory/DRAM/n3309 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][16]  ( .D(
        \unit_memory/DRAM/n1237 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n432 ), .QN(\unit_memory/DRAM/n3310 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][15]  ( .D(
        \unit_memory/DRAM/n1236 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n433 ), .QN(\unit_memory/DRAM/n3311 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][14]  ( .D(
        \unit_memory/DRAM/n1235 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n434 ), .QN(\unit_memory/DRAM/n3312 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][13]  ( .D(
        \unit_memory/DRAM/n1234 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n435 ), .QN(\unit_memory/DRAM/n3313 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][12]  ( .D(
        \unit_memory/DRAM/n1233 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n436 ), .QN(\unit_memory/DRAM/n3314 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][11]  ( .D(
        \unit_memory/DRAM/n1232 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n437 ), .QN(\unit_memory/DRAM/n3315 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][10]  ( .D(
        \unit_memory/DRAM/n1231 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n438 ), .QN(\unit_memory/DRAM/n3316 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][9]  ( .D(\unit_memory/DRAM/n1230 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n439 ), .QN(
        \unit_memory/DRAM/n3317 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][8]  ( .D(\unit_memory/DRAM/n1229 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n440 ), .QN(
        \unit_memory/DRAM/n3318 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][7]  ( .D(\unit_memory/DRAM/n1228 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n441 ), .QN(
        \unit_memory/DRAM/n3319 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][6]  ( .D(\unit_memory/DRAM/n1227 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n442 ), .QN(
        \unit_memory/DRAM/n3320 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][5]  ( .D(\unit_memory/DRAM/n1226 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n443 ), .QN(
        \unit_memory/DRAM/n3321 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][4]  ( .D(\unit_memory/DRAM/n1225 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n444 ), .QN(
        \unit_memory/DRAM/n3322 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][3]  ( .D(\unit_memory/DRAM/n1224 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n445 ), .QN(
        \unit_memory/DRAM/n3323 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][2]  ( .D(\unit_memory/DRAM/n1223 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n446 ), .QN(
        \unit_memory/DRAM/n3324 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][1]  ( .D(\unit_memory/DRAM/n1222 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n447 ), .QN(
        \unit_memory/DRAM/n3325 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[29][0]  ( .D(\unit_memory/DRAM/n1221 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n448 ), .QN(
        \unit_memory/DRAM/n3326 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][23]  ( .D(
        \unit_memory/DRAM/n1372 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n297 ), .QN(\unit_memory/DRAM/n3175 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][22]  ( .D(
        \unit_memory/DRAM/n1371 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n298 ), .QN(\unit_memory/DRAM/n3176 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][21]  ( .D(
        \unit_memory/DRAM/n1370 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n299 ), .QN(\unit_memory/DRAM/n3177 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][20]  ( .D(
        \unit_memory/DRAM/n1369 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n300 ), .QN(\unit_memory/DRAM/n3178 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][19]  ( .D(
        \unit_memory/DRAM/n1368 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n301 ), .QN(\unit_memory/DRAM/n3179 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][18]  ( .D(
        \unit_memory/DRAM/n1367 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n302 ), .QN(\unit_memory/DRAM/n3180 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][17]  ( .D(
        \unit_memory/DRAM/n1366 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n303 ), .QN(\unit_memory/DRAM/n3181 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][16]  ( .D(
        \unit_memory/DRAM/n1365 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n304 ), .QN(\unit_memory/DRAM/n3182 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][15]  ( .D(
        \unit_memory/DRAM/n1364 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n305 ), .QN(\unit_memory/DRAM/n3183 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][14]  ( .D(
        \unit_memory/DRAM/n1363 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n306 ), .QN(\unit_memory/DRAM/n3184 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][13]  ( .D(
        \unit_memory/DRAM/n1362 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n307 ), .QN(\unit_memory/DRAM/n3185 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][12]  ( .D(
        \unit_memory/DRAM/n1361 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n308 ), .QN(\unit_memory/DRAM/n3186 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][11]  ( .D(
        \unit_memory/DRAM/n1360 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n309 ), .QN(\unit_memory/DRAM/n3187 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][10]  ( .D(
        \unit_memory/DRAM/n1359 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n310 ), .QN(\unit_memory/DRAM/n3188 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][9]  ( .D(\unit_memory/DRAM/n1358 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n311 ), .QN(
        \unit_memory/DRAM/n3189 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][8]  ( .D(\unit_memory/DRAM/n1357 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n312 ), .QN(
        \unit_memory/DRAM/n3190 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][7]  ( .D(\unit_memory/DRAM/n1356 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n313 ), .QN(
        \unit_memory/DRAM/n3191 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][6]  ( .D(\unit_memory/DRAM/n1355 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n314 ), .QN(
        \unit_memory/DRAM/n3192 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][5]  ( .D(\unit_memory/DRAM/n1354 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n315 ), .QN(
        \unit_memory/DRAM/n3193 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][4]  ( .D(\unit_memory/DRAM/n1353 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n316 ), .QN(
        \unit_memory/DRAM/n3194 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][3]  ( .D(\unit_memory/DRAM/n1352 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n317 ), .QN(
        \unit_memory/DRAM/n3195 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][2]  ( .D(\unit_memory/DRAM/n1351 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n318 ), .QN(
        \unit_memory/DRAM/n3196 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][1]  ( .D(\unit_memory/DRAM/n1350 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n319 ), .QN(
        \unit_memory/DRAM/n3197 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[25][0]  ( .D(\unit_memory/DRAM/n1349 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n320 ), .QN(
        \unit_memory/DRAM/n3198 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][23]  ( .D(
        \unit_memory/DRAM/n1500 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n169 ), .QN(\unit_memory/DRAM/n3047 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][22]  ( .D(
        \unit_memory/DRAM/n1499 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n170 ), .QN(\unit_memory/DRAM/n3048 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][21]  ( .D(
        \unit_memory/DRAM/n1498 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n171 ), .QN(\unit_memory/DRAM/n3049 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][20]  ( .D(
        \unit_memory/DRAM/n1497 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n172 ), .QN(\unit_memory/DRAM/n3050 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][19]  ( .D(
        \unit_memory/DRAM/n1496 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n173 ), .QN(\unit_memory/DRAM/n3051 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][18]  ( .D(
        \unit_memory/DRAM/n1495 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n174 ), .QN(\unit_memory/DRAM/n3052 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][17]  ( .D(
        \unit_memory/DRAM/n1494 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n175 ), .QN(\unit_memory/DRAM/n3053 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][16]  ( .D(
        \unit_memory/DRAM/n1493 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n176 ), .QN(\unit_memory/DRAM/n3054 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][15]  ( .D(
        \unit_memory/DRAM/n1492 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n177 ), .QN(\unit_memory/DRAM/n3055 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][14]  ( .D(
        \unit_memory/DRAM/n1491 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n178 ), .QN(\unit_memory/DRAM/n3056 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][13]  ( .D(
        \unit_memory/DRAM/n1490 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n179 ), .QN(\unit_memory/DRAM/n3057 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][12]  ( .D(
        \unit_memory/DRAM/n1489 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n180 ), .QN(\unit_memory/DRAM/n3058 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][11]  ( .D(
        \unit_memory/DRAM/n1488 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n181 ), .QN(\unit_memory/DRAM/n3059 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][10]  ( .D(
        \unit_memory/DRAM/n1487 ), .CK(CLK), .RN(n1351), .Q(
        \unit_memory/DRAM/n182 ), .QN(\unit_memory/DRAM/n3060 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][9]  ( .D(\unit_memory/DRAM/n1486 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n183 ), .QN(
        \unit_memory/DRAM/n3061 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][8]  ( .D(\unit_memory/DRAM/n1485 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n184 ), .QN(
        \unit_memory/DRAM/n3062 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][7]  ( .D(\unit_memory/DRAM/n1484 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n185 ), .QN(
        \unit_memory/DRAM/n3063 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][6]  ( .D(\unit_memory/DRAM/n1483 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n186 ), .QN(
        \unit_memory/DRAM/n3064 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][5]  ( .D(\unit_memory/DRAM/n1482 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n187 ), .QN(
        \unit_memory/DRAM/n3065 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][4]  ( .D(\unit_memory/DRAM/n1481 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n188 ), .QN(
        \unit_memory/DRAM/n3066 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][3]  ( .D(\unit_memory/DRAM/n1480 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n189 ), .QN(
        \unit_memory/DRAM/n3067 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][2]  ( .D(\unit_memory/DRAM/n1479 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n190 ), .QN(
        \unit_memory/DRAM/n3068 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][1]  ( .D(\unit_memory/DRAM/n1478 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n191 ), .QN(
        \unit_memory/DRAM/n3069 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[21][0]  ( .D(\unit_memory/DRAM/n1477 ), .CK(CLK), .RN(n1351), .Q(\unit_memory/DRAM/n192 ), .QN(
        \unit_memory/DRAM/n3070 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][23]  ( .D(
        \unit_memory/DRAM/n1628 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n41 ), .QN(\unit_memory/DRAM/n2919 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][22]  ( .D(
        \unit_memory/DRAM/n1627 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n42 ), .QN(\unit_memory/DRAM/n2920 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][21]  ( .D(
        \unit_memory/DRAM/n1626 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n43 ), .QN(\unit_memory/DRAM/n2921 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][20]  ( .D(
        \unit_memory/DRAM/n1625 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n44 ), .QN(\unit_memory/DRAM/n2922 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][19]  ( .D(
        \unit_memory/DRAM/n1624 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n45 ), .QN(\unit_memory/DRAM/n2923 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][18]  ( .D(
        \unit_memory/DRAM/n1623 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n46 ), .QN(\unit_memory/DRAM/n2924 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][17]  ( .D(
        \unit_memory/DRAM/n1622 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n47 ), .QN(\unit_memory/DRAM/n2925 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][16]  ( .D(
        \unit_memory/DRAM/n1621 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n48 ), .QN(\unit_memory/DRAM/n2926 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][15]  ( .D(
        \unit_memory/DRAM/n1620 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n49 ), .QN(\unit_memory/DRAM/n2927 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][14]  ( .D(
        \unit_memory/DRAM/n1619 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n50 ), .QN(\unit_memory/DRAM/n2928 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][13]  ( .D(
        \unit_memory/DRAM/n1618 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n51 ), .QN(\unit_memory/DRAM/n2929 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][12]  ( .D(
        \unit_memory/DRAM/n1617 ), .CK(CLK), .RN(n55), .Q(
        \unit_memory/DRAM/n52 ), .QN(\unit_memory/DRAM/n2930 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][11]  ( .D(
        \unit_memory/DRAM/n1616 ), .CK(CLK), .RN(n54), .Q(
        \unit_memory/DRAM/n53 ), .QN(\unit_memory/DRAM/n2931 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][10]  ( .D(
        \unit_memory/DRAM/n1615 ), .CK(CLK), .RN(n53), .Q(
        \unit_memory/DRAM/n54 ), .QN(\unit_memory/DRAM/n2932 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][9]  ( .D(\unit_memory/DRAM/n1614 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n55 ), .QN(\unit_memory/DRAM/n2933 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][8]  ( .D(\unit_memory/DRAM/n1613 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n56 ), .QN(\unit_memory/DRAM/n2934 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][7]  ( .D(\unit_memory/DRAM/n1612 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n57 ), .QN(\unit_memory/DRAM/n2935 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][6]  ( .D(\unit_memory/DRAM/n1611 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n58 ), .QN(\unit_memory/DRAM/n2936 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][5]  ( .D(\unit_memory/DRAM/n1610 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n59 ), .QN(\unit_memory/DRAM/n2937 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][4]  ( .D(\unit_memory/DRAM/n1609 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n60 ), .QN(\unit_memory/DRAM/n2938 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][3]  ( .D(\unit_memory/DRAM/n1608 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n61 ), .QN(\unit_memory/DRAM/n2939 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][2]  ( .D(\unit_memory/DRAM/n1607 ), .CK(CLK), .RN(n54), .Q(\unit_memory/DRAM/n62 ), .QN(\unit_memory/DRAM/n2940 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][1]  ( .D(\unit_memory/DRAM/n1606 ), .CK(CLK), .RN(n53), .Q(\unit_memory/DRAM/n63 ), .QN(\unit_memory/DRAM/n2941 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[17][0]  ( .D(\unit_memory/DRAM/n1605 ), .CK(CLK), .RN(n55), .Q(\unit_memory/DRAM/n64 ), .QN(\unit_memory/DRAM/n2942 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][23]  ( .D(
        \unit_memory/DRAM/n1756 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2791 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][22]  ( .D(
        \unit_memory/DRAM/n1755 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2792 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][21]  ( .D(
        \unit_memory/DRAM/n1754 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2793 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][20]  ( .D(
        \unit_memory/DRAM/n1753 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2794 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][19]  ( .D(
        \unit_memory/DRAM/n1752 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2795 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][18]  ( .D(
        \unit_memory/DRAM/n1751 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2796 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][17]  ( .D(
        \unit_memory/DRAM/n1750 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2797 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][16]  ( .D(
        \unit_memory/DRAM/n1749 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2798 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][15]  ( .D(
        \unit_memory/DRAM/n1748 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2799 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][14]  ( .D(
        \unit_memory/DRAM/n1747 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2800 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][13]  ( .D(
        \unit_memory/DRAM/n1746 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2801 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][12]  ( .D(
        \unit_memory/DRAM/n1745 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2802 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][11]  ( .D(
        \unit_memory/DRAM/n1744 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2803 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][10]  ( .D(
        \unit_memory/DRAM/n1743 ), .CK(CLK), .RN(n1351), .QN(
        \unit_memory/DRAM/n2804 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][9]  ( .D(\unit_memory/DRAM/n1742 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2805 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][8]  ( .D(\unit_memory/DRAM/n1741 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2806 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][7]  ( .D(\unit_memory/DRAM/n1740 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2807 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][6]  ( .D(\unit_memory/DRAM/n1739 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2808 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][5]  ( .D(\unit_memory/DRAM/n1738 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2809 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][4]  ( .D(\unit_memory/DRAM/n1737 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2810 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][3]  ( .D(\unit_memory/DRAM/n1736 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2811 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][2]  ( .D(\unit_memory/DRAM/n1735 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2812 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][1]  ( .D(\unit_memory/DRAM/n1734 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2813 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[13][0]  ( .D(\unit_memory/DRAM/n1733 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2814 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][23]  ( .D(\unit_memory/DRAM/n1884 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2663 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][22]  ( .D(\unit_memory/DRAM/n1883 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2664 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][21]  ( .D(\unit_memory/DRAM/n1882 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2665 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][20]  ( .D(\unit_memory/DRAM/n1881 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2666 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][19]  ( .D(\unit_memory/DRAM/n1880 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2667 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][18]  ( .D(\unit_memory/DRAM/n1879 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2668 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][17]  ( .D(\unit_memory/DRAM/n1878 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2669 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][16]  ( .D(\unit_memory/DRAM/n1877 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2670 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][15]  ( .D(\unit_memory/DRAM/n1876 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2671 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][14]  ( .D(\unit_memory/DRAM/n1875 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2672 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][13]  ( .D(\unit_memory/DRAM/n1874 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2673 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][12]  ( .D(\unit_memory/DRAM/n1873 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2674 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][11]  ( .D(\unit_memory/DRAM/n1872 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2675 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][10]  ( .D(\unit_memory/DRAM/n1871 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2676 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][9]  ( .D(\unit_memory/DRAM/n1870 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2677 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][8]  ( .D(\unit_memory/DRAM/n1869 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2678 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][7]  ( .D(\unit_memory/DRAM/n1868 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2679 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][6]  ( .D(\unit_memory/DRAM/n1867 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2680 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][5]  ( .D(\unit_memory/DRAM/n1866 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2681 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][4]  ( .D(\unit_memory/DRAM/n1865 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2682 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][3]  ( .D(\unit_memory/DRAM/n1864 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2683 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][2]  ( .D(\unit_memory/DRAM/n1863 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2684 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][1]  ( .D(\unit_memory/DRAM/n1862 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2685 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[9][0]  ( .D(\unit_memory/DRAM/n1861 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2686 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][23]  ( .D(\unit_memory/DRAM/n2012 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2535 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][22]  ( .D(\unit_memory/DRAM/n2011 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2536 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][21]  ( .D(\unit_memory/DRAM/n2010 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2537 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][20]  ( .D(\unit_memory/DRAM/n2009 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2538 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][19]  ( .D(\unit_memory/DRAM/n2008 ), .CK(CLK), .RN(n53), .QN(\unit_memory/DRAM/n2539 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][18]  ( .D(\unit_memory/DRAM/n2007 ), .CK(CLK), .RN(n55), .QN(\unit_memory/DRAM/n2540 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][17]  ( .D(\unit_memory/DRAM/n2006 ), .CK(CLK), .RN(n54), .QN(\unit_memory/DRAM/n2541 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][16]  ( .D(\unit_memory/DRAM/n2005 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2542 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][15]  ( .D(\unit_memory/DRAM/n2004 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2543 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][14]  ( .D(\unit_memory/DRAM/n2003 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2544 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][13]  ( .D(\unit_memory/DRAM/n2002 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2545 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][12]  ( .D(\unit_memory/DRAM/n2001 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2546 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][11]  ( .D(\unit_memory/DRAM/n2000 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2547 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][10]  ( .D(\unit_memory/DRAM/n1999 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2548 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][9]  ( .D(\unit_memory/DRAM/n1998 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2549 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][8]  ( .D(\unit_memory/DRAM/n1997 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2550 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][7]  ( .D(\unit_memory/DRAM/n1996 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2551 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][6]  ( .D(\unit_memory/DRAM/n1995 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2552 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][5]  ( .D(\unit_memory/DRAM/n1994 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2553 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][4]  ( .D(\unit_memory/DRAM/n1993 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2554 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][3]  ( .D(\unit_memory/DRAM/n1992 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2555 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][2]  ( .D(\unit_memory/DRAM/n1991 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2556 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][1]  ( .D(\unit_memory/DRAM/n1990 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2557 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[5][0]  ( .D(\unit_memory/DRAM/n1989 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2558 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][23]  ( .D(\unit_memory/DRAM/n2140 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2407 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][22]  ( .D(\unit_memory/DRAM/n2139 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2408 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][21]  ( .D(\unit_memory/DRAM/n2138 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2409 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][20]  ( .D(\unit_memory/DRAM/n2137 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2410 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][19]  ( .D(\unit_memory/DRAM/n2136 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2411 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][18]  ( .D(\unit_memory/DRAM/n2135 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2412 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][17]  ( .D(\unit_memory/DRAM/n2134 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2413 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][16]  ( .D(\unit_memory/DRAM/n2133 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2414 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][15]  ( .D(\unit_memory/DRAM/n2132 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2415 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][14]  ( .D(\unit_memory/DRAM/n2131 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2416 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][13]  ( .D(\unit_memory/DRAM/n2130 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2417 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][12]  ( .D(\unit_memory/DRAM/n2129 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2418 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][11]  ( .D(\unit_memory/DRAM/n2128 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2419 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][10]  ( .D(\unit_memory/DRAM/n2127 ), .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2420 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][9]  ( .D(\unit_memory/DRAM/n2126 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2421 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][8]  ( .D(\unit_memory/DRAM/n2125 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2422 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][7]  ( .D(\unit_memory/DRAM/n2124 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2423 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][6]  ( .D(\unit_memory/DRAM/n2123 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2424 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][5]  ( .D(\unit_memory/DRAM/n2122 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2425 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][4]  ( .D(\unit_memory/DRAM/n2121 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2426 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][3]  ( .D(\unit_memory/DRAM/n2120 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2427 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][2]  ( .D(\unit_memory/DRAM/n2119 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2428 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][1]  ( .D(\unit_memory/DRAM/n2118 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2429 ) );
  DFFR_X1 \unit_memory/DRAM/DRAM_mem_reg[1][0]  ( .D(\unit_memory/DRAM/n2117 ), 
        .CK(CLK), .RN(n1351), .QN(\unit_memory/DRAM/n2430 ) );
  DFFR_X1 \unit_control/current_state_reg[1]  ( .D(
        \unit_control/next_state[1] ), .CK(CLK), .RN(n53), .Q(n1693), .QN(
        \unit_control/n266 ) );
  DFFR_X1 \unit_control/current_state_reg[0]  ( .D(
        \unit_control/next_state[0] ), .CK(CLK), .RN(n1351), .Q(
        \unit_control/n373 ), .QN(n1431) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[22]  ( .D(n100), .CK(
        CLK), .Q(IR_OUT[22]), .QN(\unit_decode/n2094 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_2/Q_reg  ( .D(\unit_decode/IMMreg/ffi_2/n5 ), 
        .CK(CLK), .Q(imm_out[2]), .QN(\unit_decode/n225 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_0/Q_reg  ( .D(\unit_decode/IMMreg/ffi_0/n5 ), 
        .CK(CLK), .Q(imm_out[0]), .QN(\unit_decode/n237 ) );
  DFF_X1 \unit_decode/Areg/ffi_2/Q_reg  ( .D(\unit_decode/Areg/ffi_2/n5 ), 
        .CK(CLK), .Q(rega_out[2]), .QN(\unit_decode/n193 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_2/Q_reg  ( .D(\unit_decode/NPC1reg/ffi_2/n5 ), .CK(CLK), .Q(npc1_out[2]), .QN(\unit_decode/n195 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_3/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_3/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[3] ), .QN(n1655) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_2/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_2/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[2] ), .QN(n81) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_4/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_4/n5 ), .CK(CLK), .QN(
        \unit_decode/n2144 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_6/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_6/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[6] ), .QN(n124) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_24/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_24/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[24] ), .QN(n87) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_20/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_20/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[20] ), .QN(n1567) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_10/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_10/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[10] ), .QN(n1545) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_22/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_22/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[22] ), .QN(n1573) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_23/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_23/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[23] ), .QN(n76) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_25/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_25/n5 ), .CK(CLK), .QN(n1581) );
  DFF_X1 \unit_control/uut_second_stage/ffi_24/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_24/n5 ), .CK(CLK), .Q(cw_dec[4]) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_4/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_4/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[4] ), .QN(n1539) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_31/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_31/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[31] ), .QN(n1597) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_15/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_15/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[15] ), .QN(n1651) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_16/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_16/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[16] ), .QN(n1555) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_12/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_12/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[12] ), .QN(n1551) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_29/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_29/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[29] ), .QN(n1593) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_19/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_19/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[19] ), .QN(n1565) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_17/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_17/n5 ), .CK(CLK), .QN(n1559) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[25]  ( .D(
        \unit_fetch/unit_instructionRegister/n74 ), .CK(CLK), .Q(IR_OUT[25]), 
        .QN(\unit_decode/n2091 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[26]  ( .D(
        \unit_fetch/unit_instructionRegister/n68 ), .CK(CLK), .Q(IR_OUT[26]), 
        .QN(n83) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[28]  ( .D(
        \unit_fetch/unit_instructionRegister/n69 ), .CK(CLK), .QN(
        \unit_decode/n2090 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[27]  ( .D(
        \unit_fetch/unit_instructionRegister/n73 ), .CK(CLK), .Q(IR_OUT[27]), 
        .QN(n82) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[29]  ( .D(
        \unit_fetch/unit_instructionRegister/n72 ), .CK(CLK), .Q(IR_OUT[29]), 
        .QN(n61) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[31]  ( .D(
        \unit_fetch/unit_instructionRegister/n71 ), .CK(CLK), .Q(IR_OUT[31]), 
        .QN(n62) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_7/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_7/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[7] ), .QN(n121) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_21/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_21/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[21] ), .QN(n1571) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_9/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_9/n5 ), .CK(CLK), .QN(n1543) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_8/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_8/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[8] ), .QN(n92) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_5/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_5/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[5] ), .QN(n1697) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_26/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_26/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[26] ), .QN(n1583) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_18/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_18/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[18] ), .QN(n1561) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_30/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_30/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[30] ), .QN(n1595) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_14/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_14/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[14] ), .QN(n1553) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_28/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_28/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[28] ), .QN(n1589) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_0/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_0/n5 ), .CK(CLK), .QN(n70) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_27/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_27/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[27] ), .QN(n1587) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_0/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_0/n5 ), .CK(CLK), .Q(n35), .QN(
        net130925) );
  DFF_X2 \unit_control/uut_second_stage/ffi_20/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_15/n5 ), .CK(CLK), .Q(cw_dec[0]) );
  DFF_X2 \unit_control/uut_second_stage/ffi_19/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_15/n5 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_19/n2 ) );
  DFF_X2 \unit_control/uut_second_stage/ffi_15/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_15/n5 ), .CK(CLK), .QN(
        \unit_control/n385 ) );
  DFF_X2 \unit_fetch/unit_npcregister/ffi_1/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_1/n5 ), .CK(CLK), .QN(
        \unit_decode/n2147 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_11/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_11/n5 ), .CK(CLK), .Q(
        \unit_fetch/pc_regout[11] ), .QN(n38) );
  DFF_X2 \unit_control/uut_third_stage/ffi_9/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_9/n6 ), .CK(CLK), .Q(cw_ex[0]) );
  INV_X2 U5 ( .A(bout_regn[0]), .ZN(\unit_memory/DRAM/n754 ) );
  INV_X2 U6 ( .A(bout_regn[1]), .ZN(\unit_memory/DRAM/n753 ) );
  INV_X2 U7 ( .A(bout_regn[2]), .ZN(\unit_memory/DRAM/n752 ) );
  INV_X2 U8 ( .A(bout_regn[3]), .ZN(\unit_memory/DRAM/n751 ) );
  INV_X2 U9 ( .A(bout_regn[4]), .ZN(\unit_memory/DRAM/n750 ) );
  INV_X2 U10 ( .A(bout_regn[5]), .ZN(\unit_memory/DRAM/n749 ) );
  INV_X2 U11 ( .A(bout_regn[6]), .ZN(\unit_memory/DRAM/n748 ) );
  INV_X2 U12 ( .A(bout_regn[7]), .ZN(\unit_memory/DRAM/n747 ) );
  INV_X2 U13 ( .A(\unit_memory/DRAM/n548 ), .ZN(\unit_memory/DRAM/n819 ) );
  INV_X2 U14 ( .A(\unit_memory/DRAM/n1135 ), .ZN(\unit_memory/DRAM/n1134 ) );
  INV_X2 U15 ( .A(\unit_memory/DRAM/n1114 ), .ZN(\unit_memory/DRAM/n1113 ) );
  INV_X2 U16 ( .A(\unit_memory/DRAM/n1093 ), .ZN(\unit_memory/DRAM/n1092 ) );
  INV_X2 U17 ( .A(\unit_memory/DRAM/n1072 ), .ZN(\unit_memory/DRAM/n1071 ) );
  INV_X2 U18 ( .A(\unit_memory/DRAM/n1051 ), .ZN(\unit_memory/DRAM/n1050 ) );
  INV_X2 U19 ( .A(\unit_memory/DRAM/n1030 ), .ZN(\unit_memory/DRAM/n1029 ) );
  INV_X2 U20 ( .A(\unit_memory/DRAM/n1009 ), .ZN(\unit_memory/DRAM/n1008 ) );
  INV_X2 U21 ( .A(\unit_memory/DRAM/n988 ), .ZN(\unit_memory/DRAM/n987 ) );
  INV_X2 U22 ( .A(\unit_memory/DRAM/n967 ), .ZN(\unit_memory/DRAM/n966 ) );
  INV_X2 U23 ( .A(\unit_memory/DRAM/n946 ), .ZN(\unit_memory/DRAM/n945 ) );
  INV_X2 U24 ( .A(\unit_memory/DRAM/n925 ), .ZN(\unit_memory/DRAM/n924 ) );
  INV_X2 U25 ( .A(\unit_memory/DRAM/n904 ), .ZN(\unit_memory/DRAM/n903 ) );
  INV_X2 U26 ( .A(\unit_memory/DRAM/n883 ), .ZN(\unit_memory/DRAM/n882 ) );
  INV_X2 U27 ( .A(\unit_memory/DRAM/n862 ), .ZN(\unit_memory/DRAM/n861 ) );
  INV_X2 U28 ( .A(\unit_memory/DRAM/n815 ), .ZN(\unit_memory/DRAM/n814 ) );
  INV_X2 U29 ( .A(\unit_memory/DRAM/n841 ), .ZN(\unit_memory/DRAM/n840 ) );
  INV_X2 U30 ( .A(bout_regn[15]), .ZN(\unit_memory/DRAM/n739 ) );
  INV_X2 U31 ( .A(bout_regn[16]), .ZN(\unit_memory/DRAM/n738 ) );
  INV_X2 U32 ( .A(bout_regn[17]), .ZN(\unit_memory/DRAM/n737 ) );
  INV_X2 U33 ( .A(bout_regn[18]), .ZN(\unit_memory/DRAM/n736 ) );
  INV_X2 U34 ( .A(bout_regn[19]), .ZN(\unit_memory/DRAM/n735 ) );
  INV_X2 U35 ( .A(bout_regn[20]), .ZN(\unit_memory/DRAM/n734 ) );
  INV_X2 U36 ( .A(bout_regn[21]), .ZN(\unit_memory/DRAM/n733 ) );
  INV_X2 U37 ( .A(bout_regn[22]), .ZN(\unit_memory/DRAM/n732 ) );
  INV_X2 U38 ( .A(bout_regn[23]), .ZN(\unit_memory/DRAM/n731 ) );
  INV_X2 U39 ( .A(bout_regn[24]), .ZN(\unit_memory/DRAM/n730 ) );
  INV_X2 U40 ( .A(bout_regn[25]), .ZN(\unit_memory/DRAM/n729 ) );
  INV_X2 U41 ( .A(bout_regn[26]), .ZN(\unit_memory/DRAM/n728 ) );
  INV_X2 U42 ( .A(bout_regn[27]), .ZN(\unit_memory/DRAM/n727 ) );
  INV_X2 U43 ( .A(bout_regn[28]), .ZN(\unit_memory/DRAM/n726 ) );
  INV_X2 U44 ( .A(bout_regn[29]), .ZN(\unit_memory/DRAM/n725 ) );
  INV_X2 U45 ( .A(bout_regn[30]), .ZN(\unit_memory/DRAM/n724 ) );
  INV_X2 U46 ( .A(bout_regn[31]), .ZN(\unit_memory/DRAM/n722 ) );
  INV_X2 U47 ( .A(\unit_memory/DRAM/n561 ), .ZN(\unit_memory/DRAM/n3391 ) );
  INV_X2 U48 ( .A(\unit_memory/DRAM/n699 ), .ZN(\unit_memory/DRAM/n3398 ) );
  INV_X2 U49 ( .A(\unit_memory/DRAM/n678 ), .ZN(\unit_memory/DRAM/n3397 ) );
  INV_X2 U50 ( .A(\unit_memory/DRAM/n657 ), .ZN(\unit_memory/DRAM/n3396 ) );
  INV_X2 U51 ( .A(\unit_memory/DRAM/n636 ), .ZN(\unit_memory/DRAM/n3395 ) );
  INV_X2 U52 ( .A(\unit_memory/DRAM/n615 ), .ZN(\unit_memory/DRAM/n3394 ) );
  INV_X2 U53 ( .A(\unit_memory/DRAM/n594 ), .ZN(\unit_memory/DRAM/n3393 ) );
  INV_X2 U54 ( .A(\unit_memory/DRAM/n563 ), .ZN(\unit_memory/DRAM/n3392 ) );
  INV_X2 U55 ( .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n824 ) );
  INV_X2 U56 ( .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n829 ) );
  INV_X2 U57 ( .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n834 ) );
  INV_X2 U58 ( .A(bout_regn[8]), .ZN(\unit_memory/DRAM/n746 ) );
  INV_X2 U59 ( .A(bout_regn[9]), .ZN(\unit_memory/DRAM/n745 ) );
  INV_X2 U60 ( .A(bout_regn[10]), .ZN(\unit_memory/DRAM/n744 ) );
  INV_X2 U61 ( .A(bout_regn[11]), .ZN(\unit_memory/DRAM/n743 ) );
  INV_X2 U62 ( .A(bout_regn[12]), .ZN(\unit_memory/DRAM/n742 ) );
  INV_X2 U63 ( .A(bout_regn[13]), .ZN(\unit_memory/DRAM/n741 ) );
  INV_X2 U64 ( .A(bout_regn[14]), .ZN(\unit_memory/DRAM/n740 ) );
  INV_X2 U65 ( .A(\unit_memory/DRAM/n2346 ), .ZN(\unit_memory/DRAM/N566 ) );
  INV_X2 U66 ( .A(\unit_memory/DRAM/n2325 ), .ZN(\unit_memory/DRAM/N567 ) );
  INV_X2 U67 ( .A(\unit_memory/DRAM/n2304 ), .ZN(\unit_memory/DRAM/N568 ) );
  INV_X2 U68 ( .A(\unit_memory/DRAM/n2283 ), .ZN(\unit_memory/DRAM/N569 ) );
  INV_X2 U69 ( .A(\unit_memory/DRAM/n2262 ), .ZN(\unit_memory/DRAM/N570 ) );
  INV_X2 U70 ( .A(\unit_memory/DRAM/n2241 ), .ZN(\unit_memory/DRAM/N571 ) );
  INV_X2 U71 ( .A(\unit_memory/DRAM/n2220 ), .ZN(\unit_memory/DRAM/N572 ) );
  CLKBUF_X3 U72 ( .A(net130903), .Z(n50) );
  CLKBUF_X3 U73 ( .A(net130903), .Z(net130326) );
  CLKBUF_X3 U74 ( .A(net130903), .Z(net130324) );
  XNOR2_X1 U75 ( .A(n1486), .B(n1415), .ZN(n1427) );
  NOR2_X1 U76 ( .A1(\unit_decode/n2099 ), .A2(IR_OUT[16]), .ZN(
        \unit_decode/n2873 ) );
  NOR2_X1 U77 ( .A1(\unit_decode/n2094 ), .A2(IR_OUT[21]), .ZN(
        \unit_decode/n3493 ) );
  AND3_X1 U78 ( .A1(n1432), .A2(n1352), .A3(n1431), .ZN(n90) );
  OR2_X1 U79 ( .A1(net130925), .A2(n113), .ZN(n1446) );
  AND2_X1 U80 ( .A1(\unit_memory/DRAM/n758 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n3) );
  AND2_X1 U81 ( .A1(\unit_memory/DRAM/n766 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n4) );
  AND2_X1 U82 ( .A1(\unit_memory/DRAM/n760 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n5) );
  AND2_X1 U83 ( .A1(\unit_memory/DRAM/n764 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n6) );
  AND2_X1 U84 ( .A1(\unit_memory/DRAM/n768 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n7) );
  AND2_X1 U85 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n758 ), 
        .ZN(n8) );
  AND2_X1 U86 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n766 ), 
        .ZN(n9) );
  AND2_X1 U87 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n758 ), 
        .ZN(n10) );
  AND2_X1 U88 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n766 ), 
        .ZN(n11) );
  AND2_X1 U89 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n755 ), 
        .ZN(n12) );
  AND2_X1 U90 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n760 ), 
        .ZN(n13) );
  AND2_X1 U91 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n762 ), 
        .ZN(n14) );
  AND2_X1 U92 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n764 ), 
        .ZN(n15) );
  AND2_X1 U93 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n768 ), 
        .ZN(n16) );
  AND2_X1 U94 ( .A1(\unit_memory/DRAM/n784 ), .A2(\unit_memory/DRAM/n770 ), 
        .ZN(n17) );
  AND2_X1 U95 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n755 ), 
        .ZN(n18) );
  AND2_X1 U96 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n760 ), 
        .ZN(n19) );
  AND2_X1 U97 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n762 ), 
        .ZN(n20) );
  AND2_X1 U98 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n764 ), 
        .ZN(n21) );
  AND2_X1 U99 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n768 ), 
        .ZN(n22) );
  AND2_X1 U100 ( .A1(\unit_memory/DRAM/n762 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n23) );
  AND2_X1 U101 ( .A1(\unit_memory/DRAM/n770 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(n24) );
  AND2_X1 U102 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n762 ), 
        .ZN(n25) );
  AND2_X1 U103 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n770 ), 
        .ZN(n26) );
  AND2_X1 U104 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n758 ), 
        .ZN(n27) );
  AND2_X1 U105 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n766 ), 
        .ZN(n28) );
  AND2_X1 U106 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n755 ), 
        .ZN(n29) );
  AND2_X1 U107 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n760 ), 
        .ZN(n30) );
  AND2_X1 U108 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n764 ), 
        .ZN(n31) );
  AND2_X1 U109 ( .A1(\unit_memory/DRAM/n774 ), .A2(\unit_memory/DRAM/n768 ), 
        .ZN(n32) );
  AND2_X1 U110 ( .A1(\unit_decode/n2191 ), .A2(\unit_decode/n2190 ), .ZN(n37)
         );
  AND2_X1 U111 ( .A1(n1691), .A2(n1690), .ZN(n39) );
  INV_X1 U112 ( .A(n90), .ZN(n1695) );
  NAND4_X1 U113 ( .A1(n82), .A2(\unit_decode/n2090 ), .A3(n83), .A4(n84), .ZN(
        n40) );
  NAND2_X1 U114 ( .A1(\unit_decode/n3514 ), .A2(\unit_decode/n3516 ), .ZN(n41)
         );
  NAND4_X1 U115 ( .A1(n82), .A2(\unit_decode/n2090 ), .A3(n83), .A4(n84), .ZN(
        \unit_decode/n3514 ) );
  AND3_X2 U116 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n84) );
  CLKBUF_X1 U117 ( .A(n110), .Z(n42) );
  INV_X2 U118 ( .A(n69), .ZN(net130306) );
  AND3_X1 U119 ( .A1(\unit_decode/n2192 ), .A2(\unit_decode/n2194 ), .A3(
        \unit_decode/n2193 ), .ZN(n1372) );
  INV_X1 U120 ( .A(n1425), .ZN(n43) );
  NAND2_X1 U121 ( .A1(n73), .A2(n90), .ZN(n44) );
  OR2_X2 U122 ( .A1(n93), .A2(n94), .ZN(n45) );
  OR2_X2 U123 ( .A1(n93), .A2(n94), .ZN(n46) );
  OR2_X1 U124 ( .A1(n93), .A2(n94), .ZN(n47) );
  CLKBUF_X1 U125 ( .A(n141), .Z(n48) );
  AND2_X1 U126 ( .A1(\unit_control/uut_second_stage/ffi_15/n5 ), .A2(n1669), 
        .ZN(n49) );
  NOR2_X2 U127 ( .A1(n1497), .A2(n89), .ZN(net130903) );
  NOR2_X1 U128 ( .A1(n75), .A2(n1645), .ZN(n51) );
  AOI21_X1 U129 ( .B1(alu_out[27]), .B2(n50), .A(n1586), .ZN(n52) );
  INV_X8 U130 ( .A(n1340), .ZN(n53) );
  INV_X8 U131 ( .A(n1325), .ZN(n54) );
  INV_X8 U132 ( .A(n1340), .ZN(n55) );
  INV_X32 U133 ( .A(n1343), .ZN(n1351) );
  INV_X2 U134 ( .A(net141230), .ZN(net141231) );
  AND2_X2 U135 ( .A1(n1388), .A2(n81), .ZN(n103) );
  AND4_X1 U136 ( .A1(n56), .A2(n1567), .A3(n1571), .A4(n1573), .ZN(n1358) );
  AND3_X1 U137 ( .A1(n1565), .A2(n1561), .A3(n1559), .ZN(n56) );
  OR2_X1 U138 ( .A1(n1480), .A2(n1416), .ZN(n1599) );
  INV_X1 U139 ( .A(n59), .ZN(n57) );
  INV_X1 U140 ( .A(n1406), .ZN(n58) );
  BUF_X1 U141 ( .A(n1404), .Z(n59) );
  AOI21_X1 U142 ( .B1(alu_out[17]), .B2(net130328), .A(n1558), .ZN(n60) );
  XNOR2_X1 U143 ( .A(n1417), .B(n1422), .ZN(n96) );
  INV_X1 U144 ( .A(net130326), .ZN(n64) );
  NOR2_X1 U145 ( .A1(net130302), .A2(n70), .ZN(n65) );
  NOR2_X1 U146 ( .A1(n45), .A2(net130925), .ZN(n66) );
  NOR2_X1 U147 ( .A1(n65), .A2(n66), .ZN(n67) );
  OAI21_X1 U148 ( .B1(n64), .B2(n68), .A(n67), .ZN(
        \unit_fetch/unit_npcregister/ffi_0/n5 ) );
  INV_X1 U149 ( .A(alu_out[0]), .ZN(n68) );
  OAI22_X1 U150 ( .A1(n68), .A2(n64), .B1(net126984), .B2(net130925), .ZN(
        \unit_fetch/unit_programCounter/ffi_0/n5 ) );
  INV_X1 U151 ( .A(net126982), .ZN(n69) );
  OR2_X1 U152 ( .A1(\unit_control/n266 ), .A2(\unit_control/n373 ), .ZN(n71)
         );
  NAND2_X1 U153 ( .A1(n71), .A2(n1433), .ZN(n1491) );
  CLKBUF_X1 U154 ( .A(n110), .Z(n72) );
  OR2_X1 U155 ( .A1(n123), .A2(n1692), .ZN(n73) );
  NAND2_X1 U156 ( .A1(n73), .A2(n90), .ZN(n1433) );
  CLKBUF_X1 U157 ( .A(n1417), .Z(n74) );
  NAND2_X1 U158 ( .A1(\unit_decode/n3514 ), .A2(\unit_decode/n3516 ), .ZN(
        \unit_decode/n3515 ) );
  BUF_X2 U159 ( .A(net130903), .Z(net130328) );
  AND2_X1 U160 ( .A1(alu_out[7]), .A2(net130328), .ZN(n75) );
  NOR2_X1 U161 ( .A1(n75), .A2(n1645), .ZN(n1662) );
  NOR2_X1 U162 ( .A1(n1459), .A2(n1416), .ZN(n102) );
  AND2_X1 U163 ( .A1(n110), .A2(n86), .ZN(n77) );
  AND2_X1 U164 ( .A1(n110), .A2(n86), .ZN(n127) );
  AND4_X2 U165 ( .A1(n1357), .A2(n1359), .A3(n1360), .A4(n1358), .ZN(n110) );
  NOR2_X1 U166 ( .A1(n79), .A2(n1666), .ZN(n78) );
  XNOR2_X1 U167 ( .A(n1488), .B(n1413), .ZN(n79) );
  CLKBUF_X1 U168 ( .A(\unit_fetch/pc_regout[2] ), .Z(n80) );
  BUF_X1 U169 ( .A(\unit_fetch/n329 ), .Z(n113) );
  OR2_X1 U170 ( .A1(net130304), .A2(n1581), .ZN(n85) );
  NAND2_X1 U171 ( .A1(n1629), .A2(n85), .ZN(
        \unit_fetch/unit_programCounter/ffi_25/n5 ) );
  BUF_X2 U172 ( .A(net126982), .Z(net130304) );
  AND2_X1 U173 ( .A1(n1392), .A2(n1697), .ZN(n86) );
  NAND2_X1 U174 ( .A1(n1672), .A2(n39), .ZN(
        \unit_control/uut_second_stage/ffi_4/n5 ) );
  INV_X1 U175 ( .A(n1493), .ZN(n88) );
  BUF_X1 U176 ( .A(net126982), .Z(net141181) );
  BUF_X1 U177 ( .A(n93), .Z(n115) );
  OR2_X2 U178 ( .A1(n1491), .A2(n1322), .ZN(n89) );
  XNOR2_X1 U179 ( .A(n1599), .B(n1424), .ZN(n97) );
  OR2_X1 U180 ( .A1(\unit_control/n266 ), .A2(\unit_control/n373 ), .ZN(n91)
         );
  NAND2_X1 U181 ( .A1(n91), .A2(n44), .ZN(n93) );
  BUF_X2 U182 ( .A(net130302), .Z(net141182) );
  OR2_X1 U183 ( .A1(n1322), .A2(jump), .ZN(n94) );
  AND3_X1 U184 ( .A1(n95), .A2(n96), .A3(n97), .ZN(n1426) );
  XOR2_X1 U185 ( .A(n1423), .B(n102), .Z(n95) );
  NAND2_X1 U186 ( .A1(n37), .A2(n1372), .ZN(n1694) );
  BUF_X1 U187 ( .A(n1694), .Z(n118) );
  BUF_X1 U188 ( .A(n1694), .Z(n98) );
  INV_X1 U189 ( .A(n413), .ZN(n404) );
  INV_X1 U190 ( .A(n413), .ZN(n403) );
  INV_X1 U191 ( .A(n501), .ZN(n492) );
  INV_X1 U192 ( .A(n501), .ZN(n491) );
  INV_X1 U193 ( .A(n589), .ZN(n580) );
  INV_X1 U194 ( .A(n589), .ZN(n579) );
  INV_X1 U195 ( .A(n677), .ZN(n668) );
  INV_X1 U196 ( .A(n677), .ZN(n667) );
  INV_X1 U197 ( .A(n402), .ZN(n393) );
  INV_X1 U198 ( .A(n402), .ZN(n392) );
  INV_X1 U199 ( .A(n424), .ZN(n415) );
  INV_X1 U200 ( .A(n424), .ZN(n414) );
  INV_X1 U201 ( .A(n435), .ZN(n426) );
  INV_X1 U202 ( .A(n435), .ZN(n425) );
  INV_X1 U203 ( .A(n490), .ZN(n481) );
  INV_X1 U204 ( .A(n490), .ZN(n480) );
  INV_X1 U205 ( .A(n512), .ZN(n503) );
  INV_X1 U206 ( .A(n512), .ZN(n502) );
  INV_X1 U207 ( .A(n523), .ZN(n514) );
  INV_X1 U208 ( .A(n523), .ZN(n513) );
  INV_X1 U209 ( .A(n578), .ZN(n569) );
  INV_X1 U210 ( .A(n578), .ZN(n568) );
  INV_X1 U211 ( .A(n600), .ZN(n591) );
  INV_X1 U212 ( .A(n600), .ZN(n590) );
  INV_X1 U213 ( .A(n611), .ZN(n602) );
  INV_X1 U214 ( .A(n611), .ZN(n601) );
  INV_X1 U215 ( .A(n666), .ZN(n657) );
  INV_X1 U216 ( .A(n666), .ZN(n656) );
  INV_X1 U217 ( .A(n688), .ZN(n679) );
  INV_X1 U218 ( .A(n688), .ZN(n678) );
  INV_X1 U219 ( .A(n702), .ZN(n692) );
  INV_X1 U220 ( .A(n702), .ZN(n693) );
  INV_X1 U221 ( .A(n719), .ZN(n712) );
  INV_X1 U222 ( .A(n369), .ZN(n360) );
  INV_X1 U223 ( .A(n369), .ZN(n359) );
  INV_X1 U224 ( .A(n457), .ZN(n448) );
  INV_X1 U225 ( .A(n457), .ZN(n447) );
  INV_X1 U226 ( .A(n545), .ZN(n536) );
  INV_X1 U227 ( .A(n545), .ZN(n535) );
  INV_X1 U228 ( .A(n633), .ZN(n624) );
  INV_X1 U229 ( .A(n633), .ZN(n623) );
  INV_X1 U230 ( .A(n380), .ZN(n371) );
  INV_X1 U231 ( .A(n380), .ZN(n370) );
  INV_X1 U232 ( .A(n391), .ZN(n382) );
  INV_X1 U233 ( .A(n391), .ZN(n381) );
  INV_X1 U234 ( .A(n446), .ZN(n437) );
  INV_X1 U235 ( .A(n446), .ZN(n436) );
  INV_X1 U236 ( .A(n468), .ZN(n459) );
  INV_X1 U237 ( .A(n468), .ZN(n458) );
  INV_X1 U238 ( .A(n479), .ZN(n470) );
  INV_X1 U239 ( .A(n479), .ZN(n469) );
  INV_X1 U240 ( .A(n534), .ZN(n525) );
  INV_X1 U241 ( .A(n534), .ZN(n524) );
  INV_X1 U242 ( .A(n556), .ZN(n547) );
  INV_X1 U243 ( .A(n556), .ZN(n546) );
  INV_X1 U244 ( .A(n567), .ZN(n558) );
  INV_X1 U245 ( .A(n567), .ZN(n557) );
  INV_X1 U246 ( .A(n622), .ZN(n613) );
  INV_X1 U247 ( .A(n622), .ZN(n612) );
  INV_X1 U248 ( .A(n644), .ZN(n635) );
  INV_X1 U249 ( .A(n644), .ZN(n634) );
  INV_X1 U250 ( .A(n655), .ZN(n646) );
  INV_X1 U251 ( .A(n655), .ZN(n645) );
  INV_X1 U252 ( .A(n265), .ZN(n256) );
  INV_X1 U253 ( .A(n265), .ZN(n255) );
  BUF_X1 U254 ( .A(n4), .Z(n413) );
  BUF_X1 U255 ( .A(n6), .Z(n402) );
  BUF_X1 U256 ( .A(n7), .Z(n424) );
  BUF_X1 U257 ( .A(n24), .Z(n435) );
  BUF_X1 U258 ( .A(n28), .Z(n501) );
  BUF_X1 U259 ( .A(n9), .Z(n589) );
  BUF_X1 U260 ( .A(n11), .Z(n677) );
  BUF_X1 U261 ( .A(n31), .Z(n490) );
  BUF_X1 U262 ( .A(n15), .Z(n578) );
  BUF_X1 U263 ( .A(n21), .Z(n666) );
  BUF_X1 U264 ( .A(n32), .Z(n512) );
  BUF_X1 U265 ( .A(n26), .Z(n523) );
  BUF_X1 U266 ( .A(n16), .Z(n600) );
  BUF_X1 U267 ( .A(n17), .Z(n611) );
  BUF_X1 U268 ( .A(n22), .Z(n688) );
  BUF_X1 U269 ( .A(n691), .Z(n702) );
  BUF_X1 U270 ( .A(n689), .Z(n694) );
  BUF_X1 U271 ( .A(n6), .Z(n394) );
  BUF_X1 U272 ( .A(n6), .Z(n395) );
  BUF_X1 U273 ( .A(n6), .Z(n396) );
  BUF_X1 U274 ( .A(n6), .Z(n397) );
  BUF_X1 U275 ( .A(n6), .Z(n398) );
  BUF_X1 U276 ( .A(n6), .Z(n399) );
  BUF_X1 U277 ( .A(n397), .Z(n400) );
  BUF_X1 U278 ( .A(n398), .Z(n401) );
  BUF_X1 U279 ( .A(n4), .Z(n405) );
  BUF_X1 U280 ( .A(n4), .Z(n406) );
  BUF_X1 U281 ( .A(n4), .Z(n407) );
  BUF_X1 U282 ( .A(n4), .Z(n408) );
  BUF_X1 U283 ( .A(n4), .Z(n409) );
  BUF_X1 U284 ( .A(n4), .Z(n410) );
  BUF_X1 U285 ( .A(n408), .Z(n411) );
  BUF_X1 U286 ( .A(n409), .Z(n412) );
  BUF_X1 U287 ( .A(n7), .Z(n416) );
  BUF_X1 U288 ( .A(n7), .Z(n417) );
  BUF_X1 U289 ( .A(n7), .Z(n418) );
  BUF_X1 U290 ( .A(n7), .Z(n419) );
  BUF_X1 U291 ( .A(n7), .Z(n420) );
  BUF_X1 U292 ( .A(n7), .Z(n421) );
  BUF_X1 U293 ( .A(n419), .Z(n422) );
  BUF_X1 U294 ( .A(n420), .Z(n423) );
  BUF_X1 U295 ( .A(n24), .Z(n427) );
  BUF_X1 U296 ( .A(n24), .Z(n428) );
  BUF_X1 U297 ( .A(n24), .Z(n429) );
  BUF_X1 U298 ( .A(n24), .Z(n430) );
  BUF_X1 U299 ( .A(n24), .Z(n431) );
  BUF_X1 U300 ( .A(n24), .Z(n432) );
  BUF_X1 U301 ( .A(n430), .Z(n433) );
  BUF_X1 U302 ( .A(n431), .Z(n434) );
  BUF_X1 U303 ( .A(n31), .Z(n482) );
  BUF_X1 U304 ( .A(n31), .Z(n483) );
  BUF_X1 U305 ( .A(n31), .Z(n484) );
  BUF_X1 U306 ( .A(n31), .Z(n485) );
  BUF_X1 U307 ( .A(n31), .Z(n486) );
  BUF_X1 U308 ( .A(n31), .Z(n487) );
  BUF_X1 U309 ( .A(n485), .Z(n488) );
  BUF_X1 U310 ( .A(n486), .Z(n489) );
  BUF_X1 U311 ( .A(n28), .Z(n493) );
  BUF_X1 U312 ( .A(n28), .Z(n494) );
  BUF_X1 U313 ( .A(n28), .Z(n495) );
  BUF_X1 U314 ( .A(n28), .Z(n496) );
  BUF_X1 U315 ( .A(n28), .Z(n497) );
  BUF_X1 U316 ( .A(n28), .Z(n498) );
  BUF_X1 U317 ( .A(n496), .Z(n499) );
  BUF_X1 U318 ( .A(n497), .Z(n500) );
  BUF_X1 U319 ( .A(n32), .Z(n504) );
  BUF_X1 U320 ( .A(n32), .Z(n505) );
  BUF_X1 U321 ( .A(n32), .Z(n506) );
  BUF_X1 U322 ( .A(n32), .Z(n507) );
  BUF_X1 U323 ( .A(n32), .Z(n508) );
  BUF_X1 U324 ( .A(n32), .Z(n509) );
  BUF_X1 U325 ( .A(n507), .Z(n510) );
  BUF_X1 U326 ( .A(n508), .Z(n511) );
  BUF_X1 U327 ( .A(n26), .Z(n515) );
  BUF_X1 U328 ( .A(n26), .Z(n516) );
  BUF_X1 U329 ( .A(n26), .Z(n517) );
  BUF_X1 U330 ( .A(n26), .Z(n518) );
  BUF_X1 U331 ( .A(n26), .Z(n519) );
  BUF_X1 U332 ( .A(n26), .Z(n520) );
  BUF_X1 U333 ( .A(n518), .Z(n521) );
  BUF_X1 U334 ( .A(n519), .Z(n522) );
  BUF_X1 U335 ( .A(n15), .Z(n570) );
  BUF_X1 U336 ( .A(n15), .Z(n571) );
  BUF_X1 U337 ( .A(n15), .Z(n572) );
  BUF_X1 U338 ( .A(n15), .Z(n573) );
  BUF_X1 U339 ( .A(n15), .Z(n574) );
  BUF_X1 U340 ( .A(n15), .Z(n575) );
  BUF_X1 U341 ( .A(n573), .Z(n576) );
  BUF_X1 U342 ( .A(n574), .Z(n577) );
  BUF_X1 U343 ( .A(n9), .Z(n581) );
  BUF_X1 U344 ( .A(n9), .Z(n582) );
  BUF_X1 U345 ( .A(n9), .Z(n583) );
  BUF_X1 U346 ( .A(n9), .Z(n584) );
  BUF_X1 U347 ( .A(n9), .Z(n585) );
  BUF_X1 U348 ( .A(n9), .Z(n586) );
  BUF_X1 U349 ( .A(n584), .Z(n587) );
  BUF_X1 U350 ( .A(n585), .Z(n588) );
  BUF_X1 U351 ( .A(n16), .Z(n592) );
  BUF_X1 U352 ( .A(n16), .Z(n593) );
  BUF_X1 U353 ( .A(n16), .Z(n594) );
  BUF_X1 U354 ( .A(n16), .Z(n595) );
  BUF_X1 U355 ( .A(n16), .Z(n596) );
  BUF_X1 U356 ( .A(n16), .Z(n597) );
  BUF_X1 U357 ( .A(n595), .Z(n598) );
  BUF_X1 U358 ( .A(n596), .Z(n599) );
  BUF_X1 U359 ( .A(n17), .Z(n603) );
  BUF_X1 U360 ( .A(n17), .Z(n604) );
  BUF_X1 U361 ( .A(n17), .Z(n605) );
  BUF_X1 U362 ( .A(n17), .Z(n606) );
  BUF_X1 U363 ( .A(n17), .Z(n607) );
  BUF_X1 U364 ( .A(n17), .Z(n608) );
  BUF_X1 U365 ( .A(n606), .Z(n609) );
  BUF_X1 U366 ( .A(n607), .Z(n610) );
  BUF_X1 U367 ( .A(n21), .Z(n658) );
  BUF_X1 U368 ( .A(n21), .Z(n659) );
  BUF_X1 U369 ( .A(n21), .Z(n660) );
  BUF_X1 U370 ( .A(n21), .Z(n661) );
  BUF_X1 U371 ( .A(n21), .Z(n662) );
  BUF_X1 U372 ( .A(n21), .Z(n663) );
  BUF_X1 U373 ( .A(n661), .Z(n664) );
  BUF_X1 U374 ( .A(n662), .Z(n665) );
  BUF_X1 U375 ( .A(n11), .Z(n669) );
  BUF_X1 U376 ( .A(n11), .Z(n670) );
  BUF_X1 U377 ( .A(n11), .Z(n671) );
  BUF_X1 U378 ( .A(n11), .Z(n672) );
  BUF_X1 U379 ( .A(n11), .Z(n673) );
  BUF_X1 U380 ( .A(n11), .Z(n674) );
  BUF_X1 U381 ( .A(n672), .Z(n675) );
  BUF_X1 U382 ( .A(n673), .Z(n676) );
  BUF_X1 U383 ( .A(n22), .Z(n680) );
  BUF_X1 U384 ( .A(n22), .Z(n681) );
  BUF_X1 U385 ( .A(n22), .Z(n682) );
  BUF_X1 U386 ( .A(n22), .Z(n683) );
  BUF_X1 U387 ( .A(n22), .Z(n684) );
  BUF_X1 U388 ( .A(n22), .Z(n685) );
  BUF_X1 U389 ( .A(n683), .Z(n686) );
  BUF_X1 U390 ( .A(n684), .Z(n687) );
  BUF_X1 U391 ( .A(n689), .Z(n695) );
  BUF_X1 U392 ( .A(n689), .Z(n696) );
  BUF_X1 U393 ( .A(n690), .Z(n697) );
  BUF_X1 U394 ( .A(n690), .Z(n698) );
  BUF_X1 U395 ( .A(n690), .Z(n699) );
  BUF_X1 U396 ( .A(n691), .Z(n700) );
  BUF_X1 U397 ( .A(n691), .Z(n701) );
  INV_X1 U398 ( .A(n1064), .ZN(n1057) );
  INV_X1 U399 ( .A(n1055), .ZN(n1048) );
  INV_X1 U400 ( .A(n1046), .ZN(n1039) );
  INV_X1 U401 ( .A(n1037), .ZN(n1030) );
  INV_X1 U402 ( .A(n1028), .ZN(n1021) );
  INV_X1 U403 ( .A(n965), .ZN(n958) );
  INV_X1 U404 ( .A(n1019), .ZN(n1012) );
  INV_X1 U405 ( .A(n1010), .ZN(n1003) );
  INV_X1 U406 ( .A(n1001), .ZN(n994) );
  INV_X1 U407 ( .A(n992), .ZN(n985) );
  INV_X1 U408 ( .A(n983), .ZN(n976) );
  INV_X1 U409 ( .A(n956), .ZN(n949) );
  INV_X1 U410 ( .A(n1082), .ZN(n1075) );
  INV_X1 U411 ( .A(n1073), .ZN(n1066) );
  INV_X1 U412 ( .A(n947), .ZN(n940) );
  INV_X1 U413 ( .A(n938), .ZN(n931) );
  INV_X1 U414 ( .A(n929), .ZN(n922) );
  INV_X1 U415 ( .A(n920), .ZN(n913) );
  INV_X1 U416 ( .A(n911), .ZN(n904) );
  INV_X1 U417 ( .A(n902), .ZN(n895) );
  INV_X1 U418 ( .A(n893), .ZN(n886) );
  INV_X1 U419 ( .A(n884), .ZN(n877) );
  INV_X1 U420 ( .A(n875), .ZN(n868) );
  INV_X1 U421 ( .A(n866), .ZN(n859) );
  INV_X1 U422 ( .A(n857), .ZN(n850) );
  INV_X1 U423 ( .A(n848), .ZN(n841) );
  INV_X1 U424 ( .A(n839), .ZN(n832) );
  INV_X1 U425 ( .A(n830), .ZN(n823) );
  INV_X1 U426 ( .A(n821), .ZN(n814) );
  INV_X1 U427 ( .A(n974), .ZN(n967) );
  INV_X1 U428 ( .A(n1092), .ZN(n1085) );
  INV_X1 U429 ( .A(n1092), .ZN(n1084) );
  INV_X1 U430 ( .A(n1293), .ZN(n1289) );
  INV_X1 U431 ( .A(n1293), .ZN(n1290) );
  INV_X1 U432 ( .A(n1293), .ZN(n1292) );
  INV_X1 U433 ( .A(n1293), .ZN(n1291) );
  INV_X1 U434 ( .A(n1293), .ZN(n1288) );
  INV_X1 U435 ( .A(n1293), .ZN(n1287) );
  INV_X1 U436 ( .A(n1293), .ZN(n1286) );
  INV_X1 U437 ( .A(n1293), .ZN(n1285) );
  BUF_X1 U438 ( .A(n1294), .Z(n1301) );
  BUF_X1 U439 ( .A(n1295), .Z(n1302) );
  BUF_X1 U440 ( .A(n1295), .Z(n1304) );
  BUF_X1 U441 ( .A(n1295), .Z(n1303) );
  BUF_X1 U442 ( .A(n1294), .Z(n1298) );
  BUF_X1 U443 ( .A(n1294), .Z(n1297) );
  BUF_X1 U444 ( .A(n1294), .Z(n1299) );
  BUF_X1 U445 ( .A(n1294), .Z(n1300) );
  BUF_X1 U446 ( .A(n1294), .Z(n1296) );
  BUF_X1 U447 ( .A(n720), .Z(n718) );
  BUF_X1 U448 ( .A(n720), .Z(n717) );
  BUF_X1 U449 ( .A(n720), .Z(n716) );
  BUF_X1 U450 ( .A(n720), .Z(n715) );
  BUF_X1 U451 ( .A(n720), .Z(n713) );
  BUF_X1 U452 ( .A(n720), .Z(n714) );
  BUF_X1 U453 ( .A(n720), .Z(n719) );
  BUF_X1 U454 ( .A(n3), .Z(n369) );
  BUF_X1 U455 ( .A(n5), .Z(n380) );
  BUF_X1 U456 ( .A(n23), .Z(n391) );
  BUF_X1 U457 ( .A(n27), .Z(n457) );
  BUF_X1 U458 ( .A(n8), .Z(n545) );
  BUF_X1 U459 ( .A(n10), .Z(n633) );
  BUF_X1 U460 ( .A(n29), .Z(n446) );
  BUF_X1 U461 ( .A(n12), .Z(n534) );
  BUF_X1 U462 ( .A(n18), .Z(n622) );
  BUF_X1 U463 ( .A(n30), .Z(n468) );
  BUF_X1 U464 ( .A(n25), .Z(n479) );
  BUF_X1 U465 ( .A(n13), .Z(n556) );
  BUF_X1 U466 ( .A(n14), .Z(n567) );
  BUF_X1 U467 ( .A(n19), .Z(n644) );
  BUF_X1 U468 ( .A(n20), .Z(n655) );
  BUF_X1 U469 ( .A(n254), .Z(n265) );
  BUF_X1 U470 ( .A(n3), .Z(n361) );
  BUF_X1 U471 ( .A(n3), .Z(n362) );
  BUF_X1 U472 ( .A(n3), .Z(n363) );
  BUF_X1 U473 ( .A(n3), .Z(n364) );
  BUF_X1 U474 ( .A(n3), .Z(n365) );
  BUF_X1 U475 ( .A(n3), .Z(n366) );
  BUF_X1 U476 ( .A(n364), .Z(n367) );
  BUF_X1 U477 ( .A(n365), .Z(n368) );
  BUF_X1 U478 ( .A(n5), .Z(n372) );
  BUF_X1 U479 ( .A(n5), .Z(n373) );
  BUF_X1 U480 ( .A(n5), .Z(n374) );
  BUF_X1 U481 ( .A(n5), .Z(n375) );
  BUF_X1 U482 ( .A(n5), .Z(n376) );
  BUF_X1 U483 ( .A(n5), .Z(n377) );
  BUF_X1 U484 ( .A(n375), .Z(n378) );
  BUF_X1 U485 ( .A(n376), .Z(n379) );
  BUF_X1 U486 ( .A(n23), .Z(n383) );
  BUF_X1 U487 ( .A(n23), .Z(n384) );
  BUF_X1 U488 ( .A(n23), .Z(n385) );
  BUF_X1 U489 ( .A(n23), .Z(n386) );
  BUF_X1 U490 ( .A(n23), .Z(n387) );
  BUF_X1 U491 ( .A(n23), .Z(n388) );
  BUF_X1 U492 ( .A(n386), .Z(n389) );
  BUF_X1 U493 ( .A(n387), .Z(n390) );
  BUF_X1 U494 ( .A(n29), .Z(n438) );
  BUF_X1 U495 ( .A(n29), .Z(n439) );
  BUF_X1 U496 ( .A(n29), .Z(n440) );
  BUF_X1 U497 ( .A(n29), .Z(n441) );
  BUF_X1 U498 ( .A(n29), .Z(n442) );
  BUF_X1 U499 ( .A(n29), .Z(n443) );
  BUF_X1 U500 ( .A(n441), .Z(n444) );
  BUF_X1 U501 ( .A(n442), .Z(n445) );
  BUF_X1 U502 ( .A(n27), .Z(n449) );
  BUF_X1 U503 ( .A(n27), .Z(n450) );
  BUF_X1 U504 ( .A(n27), .Z(n451) );
  BUF_X1 U505 ( .A(n27), .Z(n452) );
  BUF_X1 U506 ( .A(n27), .Z(n453) );
  BUF_X1 U507 ( .A(n27), .Z(n454) );
  BUF_X1 U508 ( .A(n452), .Z(n455) );
  BUF_X1 U509 ( .A(n453), .Z(n456) );
  BUF_X1 U510 ( .A(n30), .Z(n460) );
  BUF_X1 U511 ( .A(n30), .Z(n461) );
  BUF_X1 U512 ( .A(n30), .Z(n462) );
  BUF_X1 U513 ( .A(n30), .Z(n463) );
  BUF_X1 U514 ( .A(n30), .Z(n464) );
  BUF_X1 U515 ( .A(n30), .Z(n465) );
  BUF_X1 U516 ( .A(n463), .Z(n466) );
  BUF_X1 U517 ( .A(n464), .Z(n467) );
  BUF_X1 U518 ( .A(n25), .Z(n471) );
  BUF_X1 U519 ( .A(n25), .Z(n472) );
  BUF_X1 U520 ( .A(n25), .Z(n473) );
  BUF_X1 U521 ( .A(n25), .Z(n474) );
  BUF_X1 U522 ( .A(n25), .Z(n475) );
  BUF_X1 U523 ( .A(n25), .Z(n476) );
  BUF_X1 U524 ( .A(n474), .Z(n477) );
  BUF_X1 U525 ( .A(n475), .Z(n478) );
  BUF_X1 U526 ( .A(n12), .Z(n526) );
  BUF_X1 U527 ( .A(n12), .Z(n527) );
  BUF_X1 U528 ( .A(n12), .Z(n528) );
  BUF_X1 U529 ( .A(n12), .Z(n529) );
  BUF_X1 U530 ( .A(n12), .Z(n530) );
  BUF_X1 U531 ( .A(n12), .Z(n531) );
  BUF_X1 U532 ( .A(n529), .Z(n532) );
  BUF_X1 U533 ( .A(n530), .Z(n533) );
  BUF_X1 U534 ( .A(n8), .Z(n537) );
  BUF_X1 U535 ( .A(n8), .Z(n538) );
  BUF_X1 U536 ( .A(n8), .Z(n539) );
  BUF_X1 U537 ( .A(n8), .Z(n540) );
  BUF_X1 U538 ( .A(n8), .Z(n541) );
  BUF_X1 U539 ( .A(n8), .Z(n542) );
  BUF_X1 U540 ( .A(n540), .Z(n543) );
  BUF_X1 U541 ( .A(n541), .Z(n544) );
  BUF_X1 U542 ( .A(n13), .Z(n548) );
  BUF_X1 U543 ( .A(n13), .Z(n549) );
  BUF_X1 U544 ( .A(n13), .Z(n550) );
  BUF_X1 U545 ( .A(n13), .Z(n551) );
  BUF_X1 U546 ( .A(n13), .Z(n552) );
  BUF_X1 U547 ( .A(n13), .Z(n553) );
  BUF_X1 U548 ( .A(n551), .Z(n554) );
  BUF_X1 U549 ( .A(n552), .Z(n555) );
  BUF_X1 U550 ( .A(n14), .Z(n559) );
  BUF_X1 U551 ( .A(n14), .Z(n560) );
  BUF_X1 U552 ( .A(n14), .Z(n561) );
  BUF_X1 U553 ( .A(n14), .Z(n562) );
  BUF_X1 U554 ( .A(n14), .Z(n563) );
  BUF_X1 U555 ( .A(n14), .Z(n564) );
  BUF_X1 U556 ( .A(n562), .Z(n565) );
  BUF_X1 U557 ( .A(n563), .Z(n566) );
  BUF_X1 U558 ( .A(n18), .Z(n614) );
  BUF_X1 U559 ( .A(n18), .Z(n615) );
  BUF_X1 U560 ( .A(n18), .Z(n616) );
  BUF_X1 U561 ( .A(n18), .Z(n617) );
  BUF_X1 U562 ( .A(n18), .Z(n618) );
  BUF_X1 U563 ( .A(n18), .Z(n619) );
  BUF_X1 U564 ( .A(n617), .Z(n620) );
  BUF_X1 U565 ( .A(n618), .Z(n621) );
  BUF_X1 U566 ( .A(n10), .Z(n625) );
  BUF_X1 U567 ( .A(n10), .Z(n626) );
  BUF_X1 U568 ( .A(n10), .Z(n627) );
  BUF_X1 U569 ( .A(n10), .Z(n628) );
  BUF_X1 U570 ( .A(n10), .Z(n629) );
  BUF_X1 U571 ( .A(n10), .Z(n630) );
  BUF_X1 U572 ( .A(n628), .Z(n631) );
  BUF_X1 U573 ( .A(n629), .Z(n632) );
  BUF_X1 U574 ( .A(n19), .Z(n636) );
  BUF_X1 U575 ( .A(n19), .Z(n637) );
  BUF_X1 U576 ( .A(n19), .Z(n638) );
  BUF_X1 U577 ( .A(n19), .Z(n639) );
  BUF_X1 U578 ( .A(n19), .Z(n640) );
  BUF_X1 U579 ( .A(n19), .Z(n641) );
  BUF_X1 U580 ( .A(n639), .Z(n642) );
  BUF_X1 U581 ( .A(n640), .Z(n643) );
  BUF_X1 U582 ( .A(n20), .Z(n647) );
  BUF_X1 U583 ( .A(n20), .Z(n648) );
  BUF_X1 U584 ( .A(n20), .Z(n649) );
  BUF_X1 U585 ( .A(n20), .Z(n650) );
  BUF_X1 U586 ( .A(n20), .Z(n651) );
  BUF_X1 U587 ( .A(n20), .Z(n652) );
  BUF_X1 U588 ( .A(n650), .Z(n653) );
  BUF_X1 U589 ( .A(n651), .Z(n654) );
  BUF_X1 U590 ( .A(n252), .Z(n257) );
  BUF_X1 U591 ( .A(n252), .Z(n258) );
  BUF_X1 U592 ( .A(n252), .Z(n259) );
  BUF_X1 U593 ( .A(n253), .Z(n260) );
  BUF_X1 U594 ( .A(n253), .Z(n261) );
  BUF_X1 U595 ( .A(n253), .Z(n262) );
  BUF_X1 U596 ( .A(n254), .Z(n263) );
  BUF_X1 U597 ( .A(n254), .Z(n264) );
  AND2_X1 U598 ( .A1(n141), .A2(n1688), .ZN(n99) );
  AND2_X1 U599 ( .A1(n48), .A2(n43), .ZN(n100) );
  BUF_X1 U600 ( .A(\unit_memory/DRAM/n801 ), .Z(n691) );
  BUF_X1 U601 ( .A(\unit_memory/DRAM/n801 ), .Z(n690) );
  BUF_X1 U602 ( .A(\unit_memory/DRAM/n801 ), .Z(n689) );
  INV_X1 U603 ( .A(n1335), .ZN(n1348) );
  INV_X1 U604 ( .A(n1335), .ZN(n1349) );
  INV_X1 U605 ( .A(n1335), .ZN(n1345) );
  INV_X1 U606 ( .A(n1335), .ZN(n1346) );
  INV_X1 U607 ( .A(n1335), .ZN(n1347) );
  INV_X1 U608 ( .A(n1335), .ZN(n1350) );
  BUF_X1 U609 ( .A(n185), .Z(n192) );
  BUF_X1 U610 ( .A(n185), .Z(n193) );
  BUF_X1 U611 ( .A(n185), .Z(n195) );
  BUF_X1 U612 ( .A(n185), .Z(n194) );
  BUF_X1 U613 ( .A(n171), .Z(n174) );
  BUF_X1 U614 ( .A(n171), .Z(n175) );
  BUF_X1 U615 ( .A(n171), .Z(n177) );
  BUF_X1 U616 ( .A(n171), .Z(n178) );
  BUF_X1 U617 ( .A(n171), .Z(n176) );
  BUF_X1 U618 ( .A(n171), .Z(n173) );
  BUF_X1 U619 ( .A(n184), .Z(n187) );
  BUF_X1 U620 ( .A(n184), .Z(n188) );
  BUF_X1 U621 ( .A(n184), .Z(n190) );
  BUF_X1 U622 ( .A(n184), .Z(n191) );
  BUF_X1 U623 ( .A(n184), .Z(n189) );
  BUF_X1 U624 ( .A(n184), .Z(n186) );
  BUF_X1 U625 ( .A(n172), .Z(n179) );
  BUF_X1 U626 ( .A(n172), .Z(n180) );
  BUF_X1 U627 ( .A(n172), .Z(n182) );
  BUF_X1 U628 ( .A(n172), .Z(n181) );
  BUF_X1 U629 ( .A(\unit_decode/n2914 ), .Z(n1228) );
  BUF_X1 U630 ( .A(\unit_decode/n2914 ), .Z(n1229) );
  BUF_X1 U631 ( .A(n145), .Z(n148) );
  BUF_X1 U632 ( .A(n145), .Z(n149) );
  BUF_X1 U633 ( .A(n145), .Z(n151) );
  BUF_X1 U634 ( .A(n145), .Z(n152) );
  BUF_X1 U635 ( .A(n145), .Z(n150) );
  BUF_X1 U636 ( .A(n145), .Z(n147) );
  BUF_X1 U637 ( .A(n158), .Z(n161) );
  BUF_X1 U638 ( .A(n158), .Z(n162) );
  BUF_X1 U639 ( .A(n158), .Z(n164) );
  BUF_X1 U640 ( .A(n158), .Z(n165) );
  BUF_X1 U641 ( .A(n158), .Z(n163) );
  BUF_X1 U642 ( .A(n158), .Z(n160) );
  BUF_X1 U643 ( .A(n146), .Z(n153) );
  BUF_X1 U644 ( .A(n146), .Z(n154) );
  BUF_X1 U645 ( .A(n146), .Z(n156) );
  BUF_X1 U646 ( .A(n146), .Z(n155) );
  BUF_X1 U647 ( .A(n159), .Z(n166) );
  BUF_X1 U648 ( .A(n159), .Z(n167) );
  BUF_X1 U649 ( .A(n159), .Z(n169) );
  BUF_X1 U650 ( .A(n159), .Z(n168) );
  BUF_X1 U651 ( .A(\unit_decode/n2297 ), .Z(n1139) );
  BUF_X1 U652 ( .A(\unit_decode/n2297 ), .Z(n1138) );
  BUF_X1 U653 ( .A(\unit_decode/n2917 ), .Z(n1235) );
  BUF_X1 U654 ( .A(\unit_decode/n2917 ), .Z(n1234) );
  BUF_X1 U655 ( .A(\unit_decode/n2914 ), .Z(n1230) );
  BUF_X1 U656 ( .A(\unit_decode/n2297 ), .Z(n1140) );
  BUF_X1 U657 ( .A(\unit_decode/n2917 ), .Z(n1236) );
  BUF_X1 U658 ( .A(net126982), .Z(net130302) );
  BUF_X1 U659 ( .A(net126982), .Z(net130310) );
  BUF_X1 U660 ( .A(net126982), .Z(net130308) );
  BUF_X1 U661 ( .A(\unit_decode/n3513 ), .Z(n1294) );
  BUF_X1 U662 ( .A(\unit_decode/n2271 ), .Z(n1089) );
  BUF_X1 U663 ( .A(\unit_decode/n2271 ), .Z(n1088) );
  BUF_X1 U664 ( .A(\unit_decode/n2271 ), .Z(n1087) );
  BUF_X1 U665 ( .A(\unit_decode/n2271 ), .Z(n1086) );
  BUF_X1 U666 ( .A(\unit_decode/n2271 ), .Z(n1090) );
  BUF_X1 U667 ( .A(\unit_decode/n2271 ), .Z(n1091) );
  BUF_X1 U668 ( .A(n1083), .Z(n1081) );
  BUF_X1 U669 ( .A(n1083), .Z(n1080) );
  BUF_X1 U670 ( .A(n1083), .Z(n1079) );
  BUF_X1 U671 ( .A(n1083), .Z(n1078) );
  BUF_X1 U672 ( .A(n1074), .Z(n1072) );
  BUF_X1 U673 ( .A(n1074), .Z(n1071) );
  BUF_X1 U674 ( .A(n1074), .Z(n1070) );
  BUF_X1 U675 ( .A(n1074), .Z(n1069) );
  BUF_X1 U676 ( .A(n1065), .Z(n1063) );
  BUF_X1 U677 ( .A(n1065), .Z(n1062) );
  BUF_X1 U678 ( .A(n1065), .Z(n1061) );
  BUF_X1 U679 ( .A(n1065), .Z(n1060) );
  BUF_X1 U680 ( .A(n1056), .Z(n1054) );
  BUF_X1 U681 ( .A(n1056), .Z(n1053) );
  BUF_X1 U682 ( .A(n1056), .Z(n1052) );
  BUF_X1 U683 ( .A(n1056), .Z(n1051) );
  BUF_X1 U684 ( .A(n1047), .Z(n1045) );
  BUF_X1 U685 ( .A(n1047), .Z(n1044) );
  BUF_X1 U686 ( .A(n1047), .Z(n1043) );
  BUF_X1 U687 ( .A(n1047), .Z(n1042) );
  BUF_X1 U688 ( .A(n1038), .Z(n1036) );
  BUF_X1 U689 ( .A(n1038), .Z(n1035) );
  BUF_X1 U690 ( .A(n1038), .Z(n1034) );
  BUF_X1 U691 ( .A(n1038), .Z(n1033) );
  BUF_X1 U692 ( .A(n1029), .Z(n1027) );
  BUF_X1 U693 ( .A(n1029), .Z(n1026) );
  BUF_X1 U694 ( .A(n1029), .Z(n1025) );
  BUF_X1 U695 ( .A(n1029), .Z(n1024) );
  BUF_X1 U696 ( .A(n948), .Z(n946) );
  BUF_X1 U697 ( .A(n948), .Z(n945) );
  BUF_X1 U698 ( .A(n948), .Z(n944) );
  BUF_X1 U699 ( .A(n948), .Z(n943) );
  BUF_X1 U700 ( .A(n939), .Z(n937) );
  BUF_X1 U701 ( .A(n939), .Z(n936) );
  BUF_X1 U702 ( .A(n939), .Z(n935) );
  BUF_X1 U703 ( .A(n939), .Z(n934) );
  BUF_X1 U704 ( .A(n930), .Z(n928) );
  BUF_X1 U705 ( .A(n930), .Z(n927) );
  BUF_X1 U706 ( .A(n930), .Z(n926) );
  BUF_X1 U707 ( .A(n930), .Z(n925) );
  BUF_X1 U708 ( .A(n921), .Z(n919) );
  BUF_X1 U709 ( .A(n921), .Z(n918) );
  BUF_X1 U710 ( .A(n921), .Z(n917) );
  BUF_X1 U711 ( .A(n921), .Z(n916) );
  BUF_X1 U712 ( .A(n912), .Z(n910) );
  BUF_X1 U713 ( .A(n912), .Z(n909) );
  BUF_X1 U714 ( .A(n912), .Z(n908) );
  BUF_X1 U715 ( .A(n912), .Z(n907) );
  BUF_X1 U716 ( .A(n903), .Z(n901) );
  BUF_X1 U717 ( .A(n903), .Z(n900) );
  BUF_X1 U718 ( .A(n903), .Z(n899) );
  BUF_X1 U719 ( .A(n903), .Z(n898) );
  BUF_X1 U720 ( .A(n894), .Z(n892) );
  BUF_X1 U721 ( .A(n894), .Z(n891) );
  BUF_X1 U722 ( .A(n894), .Z(n890) );
  BUF_X1 U723 ( .A(n894), .Z(n889) );
  BUF_X1 U724 ( .A(n885), .Z(n883) );
  BUF_X1 U725 ( .A(n885), .Z(n882) );
  BUF_X1 U726 ( .A(n885), .Z(n881) );
  BUF_X1 U727 ( .A(n885), .Z(n880) );
  BUF_X1 U728 ( .A(n1020), .Z(n1013) );
  BUF_X1 U729 ( .A(n1011), .Z(n1004) );
  BUF_X1 U730 ( .A(n1002), .Z(n995) );
  BUF_X1 U731 ( .A(n993), .Z(n986) );
  BUF_X1 U732 ( .A(n984), .Z(n977) );
  BUF_X1 U733 ( .A(n975), .Z(n968) );
  BUF_X1 U734 ( .A(n966), .Z(n959) );
  BUF_X1 U735 ( .A(n957), .Z(n950) );
  BUF_X1 U736 ( .A(n948), .Z(n941) );
  BUF_X1 U737 ( .A(n939), .Z(n932) );
  BUF_X1 U738 ( .A(n939), .Z(n933) );
  BUF_X1 U739 ( .A(n930), .Z(n923) );
  BUF_X1 U740 ( .A(n930), .Z(n924) );
  BUF_X1 U741 ( .A(n921), .Z(n914) );
  BUF_X1 U742 ( .A(n921), .Z(n915) );
  BUF_X1 U743 ( .A(n912), .Z(n905) );
  BUF_X1 U744 ( .A(n912), .Z(n906) );
  BUF_X1 U745 ( .A(n903), .Z(n896) );
  BUF_X1 U746 ( .A(n903), .Z(n897) );
  BUF_X1 U747 ( .A(n894), .Z(n887) );
  BUF_X1 U748 ( .A(n894), .Z(n888) );
  BUF_X1 U749 ( .A(n885), .Z(n878) );
  BUF_X1 U750 ( .A(n885), .Z(n879) );
  BUF_X1 U751 ( .A(n1083), .Z(n1076) );
  BUF_X1 U752 ( .A(n1083), .Z(n1077) );
  BUF_X1 U753 ( .A(n1074), .Z(n1067) );
  BUF_X1 U754 ( .A(n1074), .Z(n1068) );
  BUF_X1 U755 ( .A(n1065), .Z(n1058) );
  BUF_X1 U756 ( .A(n1065), .Z(n1059) );
  BUF_X1 U757 ( .A(n1056), .Z(n1049) );
  BUF_X1 U758 ( .A(n1056), .Z(n1050) );
  BUF_X1 U759 ( .A(n1047), .Z(n1040) );
  BUF_X1 U760 ( .A(n1047), .Z(n1041) );
  BUF_X1 U761 ( .A(n1038), .Z(n1031) );
  BUF_X1 U762 ( .A(n1038), .Z(n1032) );
  BUF_X1 U763 ( .A(n1029), .Z(n1022) );
  BUF_X1 U764 ( .A(n1029), .Z(n1023) );
  BUF_X1 U765 ( .A(n1020), .Z(n1014) );
  BUF_X1 U766 ( .A(n1020), .Z(n1015) );
  BUF_X1 U767 ( .A(n1020), .Z(n1016) );
  BUF_X1 U768 ( .A(n1020), .Z(n1017) );
  BUF_X1 U769 ( .A(n1020), .Z(n1018) );
  BUF_X1 U770 ( .A(n1011), .Z(n1005) );
  BUF_X1 U771 ( .A(n1011), .Z(n1006) );
  BUF_X1 U772 ( .A(n1011), .Z(n1007) );
  BUF_X1 U773 ( .A(n1011), .Z(n1008) );
  BUF_X1 U774 ( .A(n1011), .Z(n1009) );
  BUF_X1 U775 ( .A(n1002), .Z(n996) );
  BUF_X1 U776 ( .A(n1002), .Z(n997) );
  BUF_X1 U777 ( .A(n1002), .Z(n998) );
  BUF_X1 U778 ( .A(n1002), .Z(n999) );
  BUF_X1 U779 ( .A(n1002), .Z(n1000) );
  BUF_X1 U780 ( .A(n993), .Z(n987) );
  BUF_X1 U781 ( .A(n993), .Z(n988) );
  BUF_X1 U782 ( .A(n993), .Z(n989) );
  BUF_X1 U783 ( .A(n993), .Z(n990) );
  BUF_X1 U784 ( .A(n993), .Z(n991) );
  BUF_X1 U785 ( .A(n984), .Z(n978) );
  BUF_X1 U786 ( .A(n984), .Z(n979) );
  BUF_X1 U787 ( .A(n984), .Z(n980) );
  BUF_X1 U788 ( .A(n984), .Z(n981) );
  BUF_X1 U789 ( .A(n984), .Z(n982) );
  BUF_X1 U790 ( .A(n975), .Z(n969) );
  BUF_X1 U791 ( .A(n975), .Z(n970) );
  BUF_X1 U792 ( .A(n975), .Z(n971) );
  BUF_X1 U793 ( .A(n975), .Z(n972) );
  BUF_X1 U794 ( .A(n975), .Z(n973) );
  BUF_X1 U795 ( .A(n966), .Z(n960) );
  BUF_X1 U796 ( .A(n966), .Z(n961) );
  BUF_X1 U797 ( .A(n966), .Z(n962) );
  BUF_X1 U798 ( .A(n966), .Z(n963) );
  BUF_X1 U799 ( .A(n966), .Z(n964) );
  BUF_X1 U800 ( .A(n957), .Z(n951) );
  BUF_X1 U801 ( .A(n957), .Z(n952) );
  BUF_X1 U802 ( .A(n957), .Z(n953) );
  BUF_X1 U803 ( .A(n957), .Z(n954) );
  BUF_X1 U804 ( .A(n957), .Z(n955) );
  BUF_X1 U805 ( .A(n948), .Z(n942) );
  BUF_X1 U806 ( .A(n876), .Z(n874) );
  BUF_X1 U807 ( .A(n876), .Z(n873) );
  BUF_X1 U808 ( .A(n876), .Z(n872) );
  BUF_X1 U809 ( .A(n876), .Z(n871) );
  BUF_X1 U810 ( .A(n867), .Z(n865) );
  BUF_X1 U811 ( .A(n867), .Z(n864) );
  BUF_X1 U812 ( .A(n867), .Z(n863) );
  BUF_X1 U813 ( .A(n867), .Z(n862) );
  BUF_X1 U814 ( .A(n858), .Z(n856) );
  BUF_X1 U815 ( .A(n858), .Z(n855) );
  BUF_X1 U816 ( .A(n858), .Z(n854) );
  BUF_X1 U817 ( .A(n858), .Z(n853) );
  BUF_X1 U818 ( .A(n849), .Z(n847) );
  BUF_X1 U819 ( .A(n849), .Z(n846) );
  BUF_X1 U820 ( .A(n849), .Z(n845) );
  BUF_X1 U821 ( .A(n849), .Z(n844) );
  BUF_X1 U822 ( .A(n840), .Z(n838) );
  BUF_X1 U823 ( .A(n840), .Z(n837) );
  BUF_X1 U824 ( .A(n840), .Z(n836) );
  BUF_X1 U825 ( .A(n840), .Z(n835) );
  BUF_X1 U826 ( .A(n831), .Z(n829) );
  BUF_X1 U827 ( .A(n831), .Z(n828) );
  BUF_X1 U828 ( .A(n831), .Z(n827) );
  BUF_X1 U829 ( .A(n831), .Z(n826) );
  BUF_X1 U830 ( .A(n822), .Z(n820) );
  BUF_X1 U831 ( .A(n822), .Z(n819) );
  BUF_X1 U832 ( .A(n822), .Z(n818) );
  BUF_X1 U833 ( .A(n822), .Z(n817) );
  BUF_X1 U834 ( .A(n876), .Z(n869) );
  BUF_X1 U835 ( .A(n876), .Z(n870) );
  BUF_X1 U836 ( .A(n867), .Z(n860) );
  BUF_X1 U837 ( .A(n867), .Z(n861) );
  BUF_X1 U838 ( .A(n858), .Z(n851) );
  BUF_X1 U839 ( .A(n858), .Z(n852) );
  BUF_X1 U840 ( .A(n849), .Z(n842) );
  BUF_X1 U841 ( .A(n849), .Z(n843) );
  BUF_X1 U842 ( .A(n840), .Z(n833) );
  BUF_X1 U843 ( .A(n840), .Z(n834) );
  BUF_X1 U844 ( .A(n831), .Z(n824) );
  BUF_X1 U845 ( .A(n831), .Z(n825) );
  BUF_X1 U846 ( .A(n822), .Z(n815) );
  BUF_X1 U847 ( .A(n822), .Z(n816) );
  BUF_X1 U848 ( .A(\unit_decode/n2271 ), .Z(n1092) );
  BUF_X1 U849 ( .A(n939), .Z(n938) );
  BUF_X1 U850 ( .A(n930), .Z(n929) );
  BUF_X1 U851 ( .A(n921), .Z(n920) );
  BUF_X1 U852 ( .A(n912), .Z(n911) );
  BUF_X1 U853 ( .A(n903), .Z(n902) );
  BUF_X1 U854 ( .A(n894), .Z(n893) );
  BUF_X1 U855 ( .A(n885), .Z(n884) );
  BUF_X1 U856 ( .A(n1083), .Z(n1082) );
  BUF_X1 U857 ( .A(n1074), .Z(n1073) );
  BUF_X1 U858 ( .A(n1065), .Z(n1064) );
  BUF_X1 U859 ( .A(n1056), .Z(n1055) );
  BUF_X1 U860 ( .A(n1047), .Z(n1046) );
  BUF_X1 U861 ( .A(n1038), .Z(n1037) );
  BUF_X1 U862 ( .A(n1029), .Z(n1028) );
  BUF_X1 U863 ( .A(n1020), .Z(n1019) );
  BUF_X1 U864 ( .A(n1011), .Z(n1010) );
  BUF_X1 U865 ( .A(n1002), .Z(n1001) );
  BUF_X1 U866 ( .A(n993), .Z(n992) );
  BUF_X1 U867 ( .A(n984), .Z(n983) );
  BUF_X1 U868 ( .A(n975), .Z(n974) );
  BUF_X1 U869 ( .A(n966), .Z(n965) );
  BUF_X1 U870 ( .A(n957), .Z(n956) );
  BUF_X1 U871 ( .A(n948), .Z(n947) );
  BUF_X1 U872 ( .A(n876), .Z(n875) );
  BUF_X1 U873 ( .A(n867), .Z(n866) );
  BUF_X1 U874 ( .A(n858), .Z(n857) );
  BUF_X1 U875 ( .A(n849), .Z(n848) );
  BUF_X1 U876 ( .A(n840), .Z(n839) );
  BUF_X1 U877 ( .A(n831), .Z(n830) );
  BUF_X1 U878 ( .A(n822), .Z(n821) );
  NAND2_X1 U879 ( .A1(\unit_memory/DRAM/n794 ), .A2(\unit_memory/DRAM/n770 ), 
        .ZN(\unit_memory/DRAM/n801 ) );
  BUF_X1 U880 ( .A(\unit_decode/n3513 ), .Z(n1295) );
  AND2_X1 U881 ( .A1(n1598), .A2(n1679), .ZN(n101) );
  INV_X1 U882 ( .A(\unit_decode/n2196 ), .ZN(n720) );
  OAI21_X1 U883 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2229 ), .A(n1348), .ZN(\unit_decode/n2196 ) );
  BUF_X1 U884 ( .A(\unit_memory/DRAM/n723 ), .Z(n254) );
  BUF_X1 U885 ( .A(\unit_memory/DRAM/n723 ), .Z(n252) );
  BUF_X1 U886 ( .A(\unit_memory/DRAM/n723 ), .Z(n253) );
  BUF_X1 U887 ( .A(n237), .Z(n244) );
  BUF_X1 U888 ( .A(n237), .Z(n245) );
  BUF_X1 U889 ( .A(n237), .Z(n247) );
  BUF_X1 U890 ( .A(n237), .Z(n246) );
  BUF_X1 U891 ( .A(n223), .Z(n226) );
  BUF_X1 U892 ( .A(n223), .Z(n227) );
  BUF_X1 U893 ( .A(n223), .Z(n229) );
  BUF_X1 U894 ( .A(n223), .Z(n230) );
  BUF_X1 U895 ( .A(n223), .Z(n228) );
  BUF_X1 U896 ( .A(n223), .Z(n225) );
  BUF_X1 U897 ( .A(n236), .Z(n239) );
  BUF_X1 U898 ( .A(n236), .Z(n240) );
  BUF_X1 U899 ( .A(n236), .Z(n242) );
  BUF_X1 U900 ( .A(n236), .Z(n243) );
  BUF_X1 U901 ( .A(n236), .Z(n241) );
  BUF_X1 U902 ( .A(n236), .Z(n238) );
  BUF_X1 U903 ( .A(n224), .Z(n231) );
  BUF_X1 U904 ( .A(n224), .Z(n232) );
  BUF_X1 U905 ( .A(n224), .Z(n234) );
  BUF_X1 U906 ( .A(n224), .Z(n233) );
  BUF_X1 U907 ( .A(\unit_decode/n2279 ), .Z(n1096) );
  BUF_X1 U908 ( .A(\unit_decode/n2284 ), .Z(n1108) );
  BUF_X1 U909 ( .A(\unit_decode/n2289 ), .Z(n1120) );
  BUF_X1 U910 ( .A(\unit_decode/n2294 ), .Z(n1132) );
  BUF_X1 U911 ( .A(\unit_decode/n2303 ), .Z(n1144) );
  BUF_X1 U912 ( .A(\unit_decode/n2308 ), .Z(n1156) );
  BUF_X1 U913 ( .A(\unit_decode/n2313 ), .Z(n1168) );
  BUF_X1 U914 ( .A(\unit_decode/n2318 ), .Z(n1180) );
  BUF_X1 U915 ( .A(\unit_decode/n2279 ), .Z(n1097) );
  BUF_X1 U916 ( .A(\unit_decode/n2284 ), .Z(n1109) );
  BUF_X1 U917 ( .A(\unit_decode/n2289 ), .Z(n1121) );
  BUF_X1 U918 ( .A(\unit_decode/n2294 ), .Z(n1133) );
  BUF_X1 U919 ( .A(\unit_decode/n2303 ), .Z(n1145) );
  BUF_X1 U920 ( .A(\unit_decode/n2308 ), .Z(n1157) );
  BUF_X1 U921 ( .A(\unit_decode/n2313 ), .Z(n1169) );
  BUF_X1 U922 ( .A(\unit_decode/n2318 ), .Z(n1181) );
  BUF_X1 U923 ( .A(\unit_decode/n2899 ), .Z(n1192) );
  BUF_X1 U924 ( .A(\unit_decode/n2904 ), .Z(n1204) );
  BUF_X1 U925 ( .A(\unit_decode/n2909 ), .Z(n1216) );
  BUF_X1 U926 ( .A(\unit_decode/n2923 ), .Z(n1240) );
  BUF_X1 U927 ( .A(\unit_decode/n2928 ), .Z(n1252) );
  BUF_X1 U928 ( .A(\unit_decode/n2933 ), .Z(n1264) );
  BUF_X1 U929 ( .A(\unit_decode/n2938 ), .Z(n1276) );
  BUF_X1 U930 ( .A(\unit_decode/n2899 ), .Z(n1193) );
  BUF_X1 U931 ( .A(\unit_decode/n2904 ), .Z(n1205) );
  BUF_X1 U932 ( .A(\unit_decode/n2909 ), .Z(n1217) );
  BUF_X1 U933 ( .A(\unit_decode/n2923 ), .Z(n1241) );
  BUF_X1 U934 ( .A(\unit_decode/n2928 ), .Z(n1253) );
  BUF_X1 U935 ( .A(\unit_decode/n2933 ), .Z(n1265) );
  BUF_X1 U936 ( .A(\unit_decode/n2938 ), .Z(n1277) );
  BUF_X1 U937 ( .A(n197), .Z(n200) );
  BUF_X1 U938 ( .A(n197), .Z(n201) );
  BUF_X1 U939 ( .A(n197), .Z(n203) );
  BUF_X1 U940 ( .A(n197), .Z(n204) );
  BUF_X1 U941 ( .A(n197), .Z(n202) );
  BUF_X1 U942 ( .A(n197), .Z(n199) );
  BUF_X1 U943 ( .A(n210), .Z(n213) );
  BUF_X1 U944 ( .A(n210), .Z(n214) );
  BUF_X1 U945 ( .A(n210), .Z(n216) );
  BUF_X1 U946 ( .A(n210), .Z(n217) );
  BUF_X1 U947 ( .A(n210), .Z(n215) );
  BUF_X1 U948 ( .A(n210), .Z(n212) );
  BUF_X1 U949 ( .A(n198), .Z(n205) );
  BUF_X1 U950 ( .A(n198), .Z(n206) );
  BUF_X1 U951 ( .A(n198), .Z(n208) );
  BUF_X1 U952 ( .A(n198), .Z(n207) );
  BUF_X1 U953 ( .A(\unit_decode/n2281 ), .Z(n1099) );
  BUF_X1 U954 ( .A(\unit_decode/n2286 ), .Z(n1111) );
  BUF_X1 U955 ( .A(\unit_decode/n2291 ), .Z(n1123) );
  BUF_X1 U956 ( .A(\unit_decode/n2296 ), .Z(n1135) );
  BUF_X1 U957 ( .A(\unit_decode/n2305 ), .Z(n1147) );
  BUF_X1 U958 ( .A(\unit_decode/n2310 ), .Z(n1159) );
  BUF_X1 U959 ( .A(\unit_decode/n2315 ), .Z(n1171) );
  BUF_X1 U960 ( .A(\unit_decode/n2320 ), .Z(n1183) );
  BUF_X1 U961 ( .A(\unit_decode/n2281 ), .Z(n1100) );
  BUF_X1 U962 ( .A(\unit_decode/n2286 ), .Z(n1112) );
  BUF_X1 U963 ( .A(\unit_decode/n2291 ), .Z(n1124) );
  BUF_X1 U964 ( .A(\unit_decode/n2296 ), .Z(n1136) );
  BUF_X1 U965 ( .A(\unit_decode/n2305 ), .Z(n1148) );
  BUF_X1 U966 ( .A(\unit_decode/n2310 ), .Z(n1160) );
  BUF_X1 U967 ( .A(\unit_decode/n2315 ), .Z(n1172) );
  BUF_X1 U968 ( .A(\unit_decode/n2320 ), .Z(n1184) );
  BUF_X1 U969 ( .A(\unit_decode/n2901 ), .Z(n1195) );
  BUF_X1 U970 ( .A(\unit_decode/n2906 ), .Z(n1207) );
  BUF_X1 U971 ( .A(\unit_decode/n2911 ), .Z(n1219) );
  BUF_X1 U972 ( .A(\unit_decode/n2916 ), .Z(n1231) );
  BUF_X1 U973 ( .A(\unit_decode/n2925 ), .Z(n1243) );
  BUF_X1 U974 ( .A(\unit_decode/n2930 ), .Z(n1255) );
  BUF_X1 U975 ( .A(\unit_decode/n2935 ), .Z(n1267) );
  BUF_X1 U976 ( .A(\unit_decode/n2940 ), .Z(n1279) );
  BUF_X1 U977 ( .A(\unit_decode/n2901 ), .Z(n1196) );
  BUF_X1 U978 ( .A(\unit_decode/n2906 ), .Z(n1208) );
  BUF_X1 U979 ( .A(\unit_decode/n2911 ), .Z(n1220) );
  BUF_X1 U980 ( .A(\unit_decode/n2916 ), .Z(n1232) );
  BUF_X1 U981 ( .A(\unit_decode/n2925 ), .Z(n1244) );
  BUF_X1 U982 ( .A(\unit_decode/n2930 ), .Z(n1256) );
  BUF_X1 U983 ( .A(\unit_decode/n2935 ), .Z(n1268) );
  BUF_X1 U984 ( .A(\unit_decode/n2940 ), .Z(n1280) );
  BUF_X1 U985 ( .A(\unit_decode/n2278 ), .Z(n1093) );
  BUF_X1 U986 ( .A(\unit_decode/n2283 ), .Z(n1105) );
  BUF_X1 U987 ( .A(\unit_decode/n2288 ), .Z(n1117) );
  BUF_X1 U988 ( .A(\unit_decode/n2293 ), .Z(n1129) );
  BUF_X1 U989 ( .A(\unit_decode/n2302 ), .Z(n1141) );
  BUF_X1 U990 ( .A(\unit_decode/n2307 ), .Z(n1153) );
  BUF_X1 U991 ( .A(\unit_decode/n2312 ), .Z(n1165) );
  BUF_X1 U992 ( .A(\unit_decode/n2317 ), .Z(n1177) );
  BUF_X1 U993 ( .A(\unit_decode/n2278 ), .Z(n1094) );
  BUF_X1 U994 ( .A(\unit_decode/n2283 ), .Z(n1106) );
  BUF_X1 U995 ( .A(\unit_decode/n2288 ), .Z(n1118) );
  BUF_X1 U996 ( .A(\unit_decode/n2293 ), .Z(n1130) );
  BUF_X1 U997 ( .A(\unit_decode/n2302 ), .Z(n1142) );
  BUF_X1 U998 ( .A(\unit_decode/n2307 ), .Z(n1154) );
  BUF_X1 U999 ( .A(\unit_decode/n2312 ), .Z(n1166) );
  BUF_X1 U1000 ( .A(\unit_decode/n2317 ), .Z(n1178) );
  BUF_X1 U1001 ( .A(\unit_decode/n2898 ), .Z(n1189) );
  BUF_X1 U1002 ( .A(\unit_decode/n2903 ), .Z(n1201) );
  BUF_X1 U1003 ( .A(\unit_decode/n2908 ), .Z(n1213) );
  BUF_X1 U1004 ( .A(\unit_decode/n2913 ), .Z(n1225) );
  BUF_X1 U1005 ( .A(\unit_decode/n2922 ), .Z(n1237) );
  BUF_X1 U1006 ( .A(\unit_decode/n2927 ), .Z(n1249) );
  BUF_X1 U1007 ( .A(\unit_decode/n2932 ), .Z(n1261) );
  BUF_X1 U1008 ( .A(\unit_decode/n2937 ), .Z(n1273) );
  BUF_X1 U1009 ( .A(\unit_decode/n2898 ), .Z(n1190) );
  BUF_X1 U1010 ( .A(\unit_decode/n2903 ), .Z(n1202) );
  BUF_X1 U1011 ( .A(\unit_decode/n2908 ), .Z(n1214) );
  BUF_X1 U1012 ( .A(\unit_decode/n2913 ), .Z(n1226) );
  BUF_X1 U1013 ( .A(\unit_decode/n2922 ), .Z(n1238) );
  BUF_X1 U1014 ( .A(\unit_decode/n2927 ), .Z(n1250) );
  BUF_X1 U1015 ( .A(\unit_decode/n2932 ), .Z(n1262) );
  BUF_X1 U1016 ( .A(\unit_decode/n2937 ), .Z(n1274) );
  BUF_X1 U1017 ( .A(n211), .Z(n218) );
  BUF_X1 U1018 ( .A(n211), .Z(n219) );
  BUF_X1 U1019 ( .A(n211), .Z(n221) );
  BUF_X1 U1020 ( .A(n211), .Z(n220) );
  BUF_X1 U1021 ( .A(\unit_decode/n2282 ), .Z(n1103) );
  BUF_X1 U1022 ( .A(\unit_decode/n2287 ), .Z(n1115) );
  BUF_X1 U1023 ( .A(\unit_decode/n2292 ), .Z(n1127) );
  BUF_X1 U1024 ( .A(\unit_decode/n2306 ), .Z(n1151) );
  BUF_X1 U1025 ( .A(\unit_decode/n2311 ), .Z(n1163) );
  BUF_X1 U1026 ( .A(\unit_decode/n2316 ), .Z(n1175) );
  BUF_X1 U1027 ( .A(\unit_decode/n2321 ), .Z(n1187) );
  BUF_X1 U1028 ( .A(\unit_decode/n2282 ), .Z(n1102) );
  BUF_X1 U1029 ( .A(\unit_decode/n2287 ), .Z(n1114) );
  BUF_X1 U1030 ( .A(\unit_decode/n2292 ), .Z(n1126) );
  BUF_X1 U1031 ( .A(\unit_decode/n2306 ), .Z(n1150) );
  BUF_X1 U1032 ( .A(\unit_decode/n2311 ), .Z(n1162) );
  BUF_X1 U1033 ( .A(\unit_decode/n2316 ), .Z(n1174) );
  BUF_X1 U1034 ( .A(\unit_decode/n2321 ), .Z(n1186) );
  BUF_X1 U1035 ( .A(\unit_decode/n2902 ), .Z(n1199) );
  BUF_X1 U1036 ( .A(\unit_decode/n2907 ), .Z(n1211) );
  BUF_X1 U1037 ( .A(\unit_decode/n2912 ), .Z(n1223) );
  BUF_X1 U1038 ( .A(\unit_decode/n2926 ), .Z(n1247) );
  BUF_X1 U1039 ( .A(\unit_decode/n2931 ), .Z(n1259) );
  BUF_X1 U1040 ( .A(\unit_decode/n2936 ), .Z(n1271) );
  BUF_X1 U1041 ( .A(\unit_decode/n2941 ), .Z(n1283) );
  BUF_X1 U1042 ( .A(\unit_decode/n2902 ), .Z(n1198) );
  BUF_X1 U1043 ( .A(\unit_decode/n2907 ), .Z(n1210) );
  BUF_X1 U1044 ( .A(\unit_decode/n2912 ), .Z(n1222) );
  BUF_X1 U1045 ( .A(\unit_decode/n2926 ), .Z(n1246) );
  BUF_X1 U1046 ( .A(\unit_decode/n2931 ), .Z(n1258) );
  BUF_X1 U1047 ( .A(\unit_decode/n2936 ), .Z(n1270) );
  BUF_X1 U1048 ( .A(\unit_decode/n2941 ), .Z(n1282) );
  BUF_X1 U1049 ( .A(\unit_decode/n2279 ), .Z(n1098) );
  BUF_X1 U1050 ( .A(\unit_decode/n2284 ), .Z(n1110) );
  BUF_X1 U1051 ( .A(\unit_decode/n2289 ), .Z(n1122) );
  BUF_X1 U1052 ( .A(\unit_decode/n2294 ), .Z(n1134) );
  BUF_X1 U1053 ( .A(\unit_decode/n2303 ), .Z(n1146) );
  BUF_X1 U1054 ( .A(\unit_decode/n2308 ), .Z(n1158) );
  BUF_X1 U1055 ( .A(\unit_decode/n2313 ), .Z(n1170) );
  BUF_X1 U1056 ( .A(\unit_decode/n2318 ), .Z(n1182) );
  BUF_X1 U1057 ( .A(\unit_decode/n2899 ), .Z(n1194) );
  BUF_X1 U1058 ( .A(\unit_decode/n2904 ), .Z(n1206) );
  BUF_X1 U1059 ( .A(\unit_decode/n2909 ), .Z(n1218) );
  BUF_X1 U1060 ( .A(\unit_decode/n2923 ), .Z(n1242) );
  BUF_X1 U1061 ( .A(\unit_decode/n2928 ), .Z(n1254) );
  BUF_X1 U1062 ( .A(\unit_decode/n2933 ), .Z(n1266) );
  BUF_X1 U1063 ( .A(\unit_decode/n2938 ), .Z(n1278) );
  BUF_X1 U1064 ( .A(\unit_decode/n2281 ), .Z(n1101) );
  BUF_X1 U1065 ( .A(\unit_decode/n2286 ), .Z(n1113) );
  BUF_X1 U1066 ( .A(\unit_decode/n2291 ), .Z(n1125) );
  BUF_X1 U1067 ( .A(\unit_decode/n2296 ), .Z(n1137) );
  BUF_X1 U1068 ( .A(\unit_decode/n2305 ), .Z(n1149) );
  BUF_X1 U1069 ( .A(\unit_decode/n2310 ), .Z(n1161) );
  BUF_X1 U1070 ( .A(\unit_decode/n2315 ), .Z(n1173) );
  BUF_X1 U1071 ( .A(\unit_decode/n2320 ), .Z(n1185) );
  BUF_X1 U1072 ( .A(\unit_decode/n2901 ), .Z(n1197) );
  BUF_X1 U1073 ( .A(\unit_decode/n2906 ), .Z(n1209) );
  BUF_X1 U1074 ( .A(\unit_decode/n2911 ), .Z(n1221) );
  BUF_X1 U1075 ( .A(\unit_decode/n2916 ), .Z(n1233) );
  BUF_X1 U1076 ( .A(\unit_decode/n2925 ), .Z(n1245) );
  BUF_X1 U1077 ( .A(\unit_decode/n2930 ), .Z(n1257) );
  BUF_X1 U1078 ( .A(\unit_decode/n2935 ), .Z(n1269) );
  BUF_X1 U1079 ( .A(\unit_decode/n2940 ), .Z(n1281) );
  BUF_X1 U1080 ( .A(\unit_decode/n2278 ), .Z(n1095) );
  BUF_X1 U1081 ( .A(\unit_decode/n2283 ), .Z(n1107) );
  BUF_X1 U1082 ( .A(\unit_decode/n2288 ), .Z(n1119) );
  BUF_X1 U1083 ( .A(\unit_decode/n2302 ), .Z(n1143) );
  BUF_X1 U1084 ( .A(\unit_decode/n2307 ), .Z(n1155) );
  BUF_X1 U1085 ( .A(\unit_decode/n2312 ), .Z(n1167) );
  BUF_X1 U1086 ( .A(\unit_decode/n2317 ), .Z(n1179) );
  BUF_X1 U1087 ( .A(\unit_decode/n2293 ), .Z(n1131) );
  BUF_X1 U1088 ( .A(\unit_decode/n2898 ), .Z(n1191) );
  BUF_X1 U1089 ( .A(\unit_decode/n2903 ), .Z(n1203) );
  BUF_X1 U1090 ( .A(\unit_decode/n2908 ), .Z(n1215) );
  BUF_X1 U1091 ( .A(\unit_decode/n2913 ), .Z(n1227) );
  BUF_X1 U1092 ( .A(\unit_decode/n2922 ), .Z(n1239) );
  BUF_X1 U1093 ( .A(\unit_decode/n2927 ), .Z(n1251) );
  BUF_X1 U1094 ( .A(\unit_decode/n2932 ), .Z(n1263) );
  BUF_X1 U1095 ( .A(\unit_decode/n2937 ), .Z(n1275) );
  BUF_X1 U1096 ( .A(\unit_decode/n2282 ), .Z(n1104) );
  BUF_X1 U1097 ( .A(\unit_decode/n2287 ), .Z(n1116) );
  BUF_X1 U1098 ( .A(\unit_decode/n2292 ), .Z(n1128) );
  BUF_X1 U1099 ( .A(\unit_decode/n2306 ), .Z(n1152) );
  BUF_X1 U1100 ( .A(\unit_decode/n2311 ), .Z(n1164) );
  BUF_X1 U1101 ( .A(\unit_decode/n2316 ), .Z(n1176) );
  BUF_X1 U1102 ( .A(\unit_decode/n2321 ), .Z(n1188) );
  BUF_X1 U1103 ( .A(\unit_decode/n2902 ), .Z(n1200) );
  BUF_X1 U1104 ( .A(\unit_decode/n2907 ), .Z(n1212) );
  BUF_X1 U1105 ( .A(\unit_decode/n2912 ), .Z(n1224) );
  BUF_X1 U1106 ( .A(\unit_decode/n2926 ), .Z(n1248) );
  BUF_X1 U1107 ( .A(\unit_decode/n2931 ), .Z(n1260) );
  BUF_X1 U1108 ( .A(\unit_decode/n2936 ), .Z(n1272) );
  BUF_X1 U1109 ( .A(\unit_decode/n2941 ), .Z(n1284) );
  BUF_X1 U1110 ( .A(\unit_memory/DRAM/n574 ), .Z(n171) );
  BUF_X1 U1111 ( .A(\unit_memory/DRAM/n575 ), .Z(n184) );
  BUF_X1 U1112 ( .A(\unit_memory/DRAM/n571 ), .Z(n145) );
  BUF_X1 U1113 ( .A(\unit_memory/DRAM/n572 ), .Z(n158) );
  BUF_X1 U1114 ( .A(n1336), .Z(n1335) );
  NAND2_X1 U1115 ( .A1(\unit_decode/n3490 ), .A2(\unit_decode/n3499 ), .ZN(
        \unit_decode/n2914 ) );
  BUF_X1 U1116 ( .A(\unit_memory/DRAM/n575 ), .Z(n185) );
  BUF_X1 U1117 ( .A(\unit_memory/DRAM/n574 ), .Z(n172) );
  BUF_X1 U1118 ( .A(\unit_memory/DRAM/n571 ), .Z(n146) );
  BUF_X1 U1119 ( .A(\unit_memory/DRAM/n572 ), .Z(n159) );
  BUF_X1 U1120 ( .A(n1341), .Z(n1322) );
  AND2_X1 U1121 ( .A1(\unit_decode/n2872 ), .A2(\unit_decode/n2879 ), .ZN(
        \unit_decode/n2297 ) );
  AND2_X1 U1122 ( .A1(\unit_decode/n3492 ), .A2(\unit_decode/n3499 ), .ZN(
        \unit_decode/n2917 ) );
  BUF_X1 U1123 ( .A(n1337), .Z(n1333) );
  BUF_X1 U1124 ( .A(n1340), .Z(n1325) );
  BUF_X1 U1125 ( .A(n1340), .Z(n1326) );
  BUF_X1 U1126 ( .A(n1340), .Z(n1324) );
  BUF_X1 U1127 ( .A(n1341), .Z(n1323) );
  BUF_X1 U1128 ( .A(n1339), .Z(n1327) );
  BUF_X1 U1129 ( .A(n1339), .Z(n1329) );
  BUF_X1 U1130 ( .A(n1339), .Z(n1328) );
  BUF_X1 U1131 ( .A(n1337), .Z(n1334) );
  BUF_X1 U1132 ( .A(n1338), .Z(n1331) );
  BUF_X1 U1133 ( .A(n1338), .Z(n1332) );
  BUF_X1 U1134 ( .A(n1338), .Z(n1330) );
  INV_X1 U1135 ( .A(\unit_memory/DRAM/n1148 ), .ZN(\unit_memory/DRAM/n550 ) );
  INV_X1 U1136 ( .A(\unit_memory/DRAM/n1143 ), .ZN(\unit_memory/DRAM/n551 ) );
  INV_X1 U1137 ( .A(n1321), .ZN(n1314) );
  INV_X1 U1138 ( .A(n1313), .ZN(n1306) );
  OAI21_X1 U1139 ( .B1(\unit_decode/n2243 ), .B2(\unit_decode/n2264 ), .A(
        n1350), .ZN(\unit_decode/n2271 ) );
  INV_X1 U1140 ( .A(\unit_decode/n2252 ), .ZN(n939) );
  OAI21_X1 U1141 ( .B1(\unit_decode/n2241 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2252 ) );
  INV_X1 U1142 ( .A(\unit_decode/n2251 ), .ZN(n930) );
  OAI21_X1 U1143 ( .B1(\unit_decode/n2239 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2251 ) );
  INV_X1 U1144 ( .A(\unit_decode/n2250 ), .ZN(n921) );
  OAI21_X1 U1145 ( .B1(\unit_decode/n2237 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2250 ) );
  INV_X1 U1146 ( .A(\unit_decode/n2249 ), .ZN(n912) );
  OAI21_X1 U1147 ( .B1(\unit_decode/n2235 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2249 ) );
  INV_X1 U1148 ( .A(\unit_decode/n2248 ), .ZN(n903) );
  OAI21_X1 U1149 ( .B1(\unit_decode/n2233 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2248 ) );
  INV_X1 U1150 ( .A(\unit_decode/n2247 ), .ZN(n894) );
  OAI21_X1 U1151 ( .B1(\unit_decode/n2231 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2247 ) );
  INV_X1 U1152 ( .A(\unit_decode/n2245 ), .ZN(n885) );
  OAI21_X1 U1153 ( .B1(\unit_decode/n2229 ), .B2(\unit_decode/n2246 ), .A(
        n1348), .ZN(\unit_decode/n2245 ) );
  INV_X1 U1154 ( .A(\unit_decode/n2262 ), .ZN(n1020) );
  OAI21_X1 U1155 ( .B1(\unit_decode/n2243 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2262 ) );
  INV_X1 U1156 ( .A(\unit_decode/n2261 ), .ZN(n1011) );
  OAI21_X1 U1157 ( .B1(\unit_decode/n2241 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2261 ) );
  INV_X1 U1158 ( .A(\unit_decode/n2260 ), .ZN(n1002) );
  OAI21_X1 U1159 ( .B1(\unit_decode/n2239 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2260 ) );
  INV_X1 U1160 ( .A(\unit_decode/n2259 ), .ZN(n993) );
  OAI21_X1 U1161 ( .B1(\unit_decode/n2237 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2259 ) );
  INV_X1 U1162 ( .A(\unit_decode/n2258 ), .ZN(n984) );
  OAI21_X1 U1163 ( .B1(\unit_decode/n2235 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2258 ) );
  INV_X1 U1164 ( .A(\unit_decode/n2257 ), .ZN(n975) );
  OAI21_X1 U1165 ( .B1(\unit_decode/n2233 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2257 ) );
  INV_X1 U1166 ( .A(\unit_decode/n2256 ), .ZN(n966) );
  OAI21_X1 U1167 ( .B1(\unit_decode/n2231 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2256 ) );
  INV_X1 U1168 ( .A(\unit_decode/n2254 ), .ZN(n957) );
  OAI21_X1 U1169 ( .B1(\unit_decode/n2229 ), .B2(\unit_decode/n2255 ), .A(
        n1349), .ZN(\unit_decode/n2254 ) );
  INV_X1 U1170 ( .A(\unit_decode/n2253 ), .ZN(n948) );
  OAI21_X1 U1171 ( .B1(\unit_decode/n2243 ), .B2(\unit_decode/n2246 ), .A(
        n1349), .ZN(\unit_decode/n2253 ) );
  NOR2_X1 U1172 ( .A1(\unit_memory/DRAM/n550 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n766 ) );
  NOR2_X1 U1173 ( .A1(\unit_memory/DRAM/n551 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n764 ) );
  NOR2_X1 U1174 ( .A1(\unit_memory/DRAM/n583 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n768 ) );
  NOR2_X1 U1175 ( .A1(\unit_memory/DRAM/n570 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n770 ) );
  AND2_X1 U1176 ( .A1(\unit_memory/DRAM/n771 ), .A2(\unit_memory/DRAM/n772 ), 
        .ZN(\unit_memory/DRAM/n756 ) );
  AND2_X1 U1177 ( .A1(\unit_memory/DRAM/n771 ), .A2(\unit_memory/DRAM/n782 ), 
        .ZN(\unit_memory/DRAM/n774 ) );
  AND2_X1 U1178 ( .A1(\unit_memory/DRAM/n771 ), .A2(\unit_memory/DRAM/n809 ), 
        .ZN(\unit_memory/DRAM/n794 ) );
  AND2_X1 U1179 ( .A1(\unit_memory/DRAM/n771 ), .A2(\unit_memory/DRAM/n792 ), 
        .ZN(\unit_memory/DRAM/n784 ) );
  BUF_X1 U1180 ( .A(\unit_memory/DRAM/n724 ), .Z(n266) );
  BUF_X1 U1181 ( .A(\unit_memory/DRAM/n725 ), .Z(n269) );
  BUF_X1 U1182 ( .A(\unit_memory/DRAM/n726 ), .Z(n272) );
  BUF_X1 U1183 ( .A(\unit_memory/DRAM/n727 ), .Z(n275) );
  BUF_X1 U1184 ( .A(\unit_memory/DRAM/n728 ), .Z(n278) );
  BUF_X1 U1185 ( .A(\unit_memory/DRAM/n729 ), .Z(n281) );
  BUF_X1 U1186 ( .A(\unit_memory/DRAM/n730 ), .Z(n284) );
  BUF_X1 U1187 ( .A(\unit_memory/DRAM/n731 ), .Z(n287) );
  BUF_X1 U1188 ( .A(\unit_memory/DRAM/n732 ), .Z(n290) );
  BUF_X1 U1189 ( .A(\unit_memory/DRAM/n733 ), .Z(n293) );
  BUF_X1 U1190 ( .A(\unit_memory/DRAM/n734 ), .Z(n296) );
  BUF_X1 U1191 ( .A(\unit_memory/DRAM/n735 ), .Z(n299) );
  BUF_X1 U1192 ( .A(\unit_memory/DRAM/n736 ), .Z(n302) );
  BUF_X1 U1193 ( .A(\unit_memory/DRAM/n737 ), .Z(n305) );
  BUF_X1 U1194 ( .A(\unit_memory/DRAM/n738 ), .Z(n308) );
  BUF_X1 U1195 ( .A(\unit_memory/DRAM/n739 ), .Z(n311) );
  BUF_X1 U1196 ( .A(\unit_memory/DRAM/n740 ), .Z(n314) );
  BUF_X1 U1197 ( .A(\unit_memory/DRAM/n741 ), .Z(n317) );
  BUF_X1 U1198 ( .A(\unit_memory/DRAM/n742 ), .Z(n320) );
  BUF_X1 U1199 ( .A(\unit_memory/DRAM/n743 ), .Z(n323) );
  BUF_X1 U1200 ( .A(\unit_memory/DRAM/n744 ), .Z(n326) );
  BUF_X1 U1201 ( .A(\unit_memory/DRAM/n745 ), .Z(n329) );
  BUF_X1 U1202 ( .A(\unit_memory/DRAM/n746 ), .Z(n332) );
  BUF_X1 U1203 ( .A(\unit_memory/DRAM/n747 ), .Z(n335) );
  BUF_X1 U1204 ( .A(\unit_memory/DRAM/n748 ), .Z(n338) );
  BUF_X1 U1205 ( .A(\unit_memory/DRAM/n749 ), .Z(n341) );
  BUF_X1 U1206 ( .A(\unit_memory/DRAM/n750 ), .Z(n344) );
  BUF_X1 U1207 ( .A(\unit_memory/DRAM/n751 ), .Z(n347) );
  BUF_X1 U1208 ( .A(\unit_memory/DRAM/n752 ), .Z(n350) );
  BUF_X1 U1209 ( .A(\unit_memory/DRAM/n753 ), .Z(n353) );
  BUF_X1 U1210 ( .A(\unit_memory/DRAM/n754 ), .Z(n356) );
  BUF_X1 U1211 ( .A(\unit_memory/DRAM/n724 ), .Z(n267) );
  BUF_X1 U1212 ( .A(\unit_memory/DRAM/n725 ), .Z(n270) );
  BUF_X1 U1213 ( .A(\unit_memory/DRAM/n726 ), .Z(n273) );
  BUF_X1 U1214 ( .A(\unit_memory/DRAM/n727 ), .Z(n276) );
  BUF_X1 U1215 ( .A(\unit_memory/DRAM/n728 ), .Z(n279) );
  BUF_X1 U1216 ( .A(\unit_memory/DRAM/n729 ), .Z(n282) );
  BUF_X1 U1217 ( .A(\unit_memory/DRAM/n730 ), .Z(n285) );
  BUF_X1 U1218 ( .A(\unit_memory/DRAM/n731 ), .Z(n288) );
  BUF_X1 U1219 ( .A(\unit_memory/DRAM/n732 ), .Z(n291) );
  BUF_X1 U1220 ( .A(\unit_memory/DRAM/n733 ), .Z(n294) );
  BUF_X1 U1221 ( .A(\unit_memory/DRAM/n734 ), .Z(n297) );
  BUF_X1 U1222 ( .A(\unit_memory/DRAM/n735 ), .Z(n300) );
  BUF_X1 U1223 ( .A(\unit_memory/DRAM/n736 ), .Z(n303) );
  BUF_X1 U1224 ( .A(\unit_memory/DRAM/n737 ), .Z(n306) );
  BUF_X1 U1225 ( .A(\unit_memory/DRAM/n738 ), .Z(n309) );
  BUF_X1 U1226 ( .A(\unit_memory/DRAM/n739 ), .Z(n312) );
  BUF_X1 U1227 ( .A(\unit_memory/DRAM/n740 ), .Z(n315) );
  BUF_X1 U1228 ( .A(\unit_memory/DRAM/n741 ), .Z(n318) );
  BUF_X1 U1229 ( .A(\unit_memory/DRAM/n742 ), .Z(n321) );
  BUF_X1 U1230 ( .A(\unit_memory/DRAM/n743 ), .Z(n324) );
  BUF_X1 U1231 ( .A(\unit_memory/DRAM/n744 ), .Z(n327) );
  BUF_X1 U1232 ( .A(\unit_memory/DRAM/n745 ), .Z(n330) );
  BUF_X1 U1233 ( .A(\unit_memory/DRAM/n746 ), .Z(n333) );
  BUF_X1 U1234 ( .A(\unit_memory/DRAM/n747 ), .Z(n336) );
  BUF_X1 U1235 ( .A(\unit_memory/DRAM/n748 ), .Z(n339) );
  BUF_X1 U1236 ( .A(\unit_memory/DRAM/n749 ), .Z(n342) );
  BUF_X1 U1237 ( .A(\unit_memory/DRAM/n750 ), .Z(n345) );
  BUF_X1 U1238 ( .A(\unit_memory/DRAM/n751 ), .Z(n348) );
  BUF_X1 U1239 ( .A(\unit_memory/DRAM/n752 ), .Z(n351) );
  BUF_X1 U1240 ( .A(\unit_memory/DRAM/n753 ), .Z(n354) );
  BUF_X1 U1241 ( .A(\unit_memory/DRAM/n754 ), .Z(n357) );
  BUF_X1 U1242 ( .A(\unit_decode/n2227 ), .Z(n811) );
  BUF_X1 U1243 ( .A(\unit_decode/n2226 ), .Z(n808) );
  BUF_X1 U1244 ( .A(\unit_decode/n2225 ), .Z(n805) );
  BUF_X1 U1245 ( .A(\unit_decode/n2224 ), .Z(n802) );
  BUF_X1 U1246 ( .A(\unit_decode/n2223 ), .Z(n799) );
  BUF_X1 U1247 ( .A(\unit_decode/n2222 ), .Z(n796) );
  BUF_X1 U1248 ( .A(\unit_decode/n2221 ), .Z(n793) );
  BUF_X1 U1249 ( .A(\unit_decode/n2220 ), .Z(n790) );
  BUF_X1 U1250 ( .A(\unit_decode/n2219 ), .Z(n787) );
  BUF_X1 U1251 ( .A(\unit_decode/n2218 ), .Z(n784) );
  BUF_X1 U1252 ( .A(\unit_decode/n2217 ), .Z(n781) );
  BUF_X1 U1253 ( .A(\unit_decode/n2216 ), .Z(n778) );
  BUF_X1 U1254 ( .A(\unit_decode/n2215 ), .Z(n775) );
  BUF_X1 U1255 ( .A(\unit_decode/n2214 ), .Z(n772) );
  BUF_X1 U1256 ( .A(\unit_decode/n2213 ), .Z(n769) );
  BUF_X1 U1257 ( .A(\unit_decode/n2212 ), .Z(n766) );
  BUF_X1 U1258 ( .A(\unit_decode/n2211 ), .Z(n763) );
  BUF_X1 U1259 ( .A(\unit_decode/n2210 ), .Z(n760) );
  BUF_X1 U1260 ( .A(\unit_decode/n2209 ), .Z(n757) );
  BUF_X1 U1261 ( .A(\unit_decode/n2208 ), .Z(n754) );
  BUF_X1 U1262 ( .A(\unit_decode/n2207 ), .Z(n751) );
  BUF_X1 U1263 ( .A(\unit_decode/n2206 ), .Z(n748) );
  BUF_X1 U1264 ( .A(\unit_decode/n2205 ), .Z(n745) );
  BUF_X1 U1265 ( .A(\unit_decode/n2204 ), .Z(n742) );
  BUF_X1 U1266 ( .A(\unit_decode/n2195 ), .Z(n710) );
  BUF_X1 U1267 ( .A(\unit_decode/n2197 ), .Z(n722) );
  BUF_X1 U1268 ( .A(\unit_decode/n2198 ), .Z(n725) );
  BUF_X1 U1269 ( .A(\unit_decode/n2199 ), .Z(n728) );
  BUF_X1 U1270 ( .A(\unit_decode/n2200 ), .Z(n731) );
  BUF_X1 U1271 ( .A(\unit_decode/n2201 ), .Z(n734) );
  BUF_X1 U1272 ( .A(\unit_decode/n2202 ), .Z(n737) );
  BUF_X1 U1273 ( .A(\unit_decode/n2203 ), .Z(n740) );
  BUF_X1 U1274 ( .A(\unit_decode/n2195 ), .Z(n709) );
  BUF_X1 U1275 ( .A(\unit_decode/n2197 ), .Z(n721) );
  BUF_X1 U1276 ( .A(\unit_decode/n2198 ), .Z(n724) );
  BUF_X1 U1277 ( .A(\unit_decode/n2199 ), .Z(n727) );
  BUF_X1 U1278 ( .A(\unit_decode/n2200 ), .Z(n730) );
  BUF_X1 U1279 ( .A(\unit_decode/n2201 ), .Z(n733) );
  BUF_X1 U1280 ( .A(\unit_decode/n2202 ), .Z(n736) );
  BUF_X1 U1281 ( .A(\unit_decode/n2203 ), .Z(n739) );
  BUF_X1 U1282 ( .A(\unit_decode/n2205 ), .Z(n746) );
  BUF_X1 U1283 ( .A(\unit_decode/n2206 ), .Z(n749) );
  BUF_X1 U1284 ( .A(\unit_decode/n2207 ), .Z(n752) );
  BUF_X1 U1285 ( .A(\unit_decode/n2208 ), .Z(n755) );
  BUF_X1 U1286 ( .A(\unit_decode/n2209 ), .Z(n758) );
  BUF_X1 U1287 ( .A(\unit_decode/n2210 ), .Z(n761) );
  BUF_X1 U1288 ( .A(\unit_decode/n2211 ), .Z(n764) );
  BUF_X1 U1289 ( .A(\unit_decode/n2212 ), .Z(n767) );
  BUF_X1 U1290 ( .A(\unit_decode/n2213 ), .Z(n770) );
  BUF_X1 U1291 ( .A(\unit_decode/n2214 ), .Z(n773) );
  BUF_X1 U1292 ( .A(\unit_decode/n2215 ), .Z(n776) );
  BUF_X1 U1293 ( .A(\unit_decode/n2216 ), .Z(n779) );
  BUF_X1 U1294 ( .A(\unit_decode/n2217 ), .Z(n782) );
  BUF_X1 U1295 ( .A(\unit_decode/n2218 ), .Z(n785) );
  BUF_X1 U1296 ( .A(\unit_decode/n2219 ), .Z(n788) );
  BUF_X1 U1297 ( .A(\unit_decode/n2220 ), .Z(n791) );
  BUF_X1 U1298 ( .A(\unit_decode/n2221 ), .Z(n794) );
  BUF_X1 U1299 ( .A(\unit_decode/n2222 ), .Z(n797) );
  BUF_X1 U1300 ( .A(\unit_decode/n2223 ), .Z(n800) );
  BUF_X1 U1301 ( .A(\unit_decode/n2224 ), .Z(n803) );
  BUF_X1 U1302 ( .A(\unit_decode/n2225 ), .Z(n806) );
  BUF_X1 U1303 ( .A(\unit_decode/n2226 ), .Z(n809) );
  BUF_X1 U1304 ( .A(\unit_decode/n2227 ), .Z(n812) );
  BUF_X1 U1305 ( .A(\unit_decode/n2204 ), .Z(n743) );
  BUF_X1 U1306 ( .A(\unit_memory/DRAM/n722 ), .Z(n249) );
  BUF_X1 U1307 ( .A(\unit_memory/DRAM/n722 ), .Z(n250) );
  BUF_X1 U1308 ( .A(\unit_decode/n2219 ), .Z(n789) );
  BUF_X1 U1309 ( .A(\unit_decode/n2218 ), .Z(n786) );
  BUF_X1 U1310 ( .A(\unit_decode/n2217 ), .Z(n783) );
  BUF_X1 U1311 ( .A(\unit_decode/n2216 ), .Z(n780) );
  BUF_X1 U1312 ( .A(\unit_decode/n2215 ), .Z(n777) );
  BUF_X1 U1313 ( .A(\unit_decode/n2214 ), .Z(n774) );
  BUF_X1 U1314 ( .A(\unit_decode/n2213 ), .Z(n771) );
  BUF_X1 U1315 ( .A(\unit_decode/n2212 ), .Z(n768) );
  BUF_X1 U1316 ( .A(\unit_decode/n2211 ), .Z(n765) );
  BUF_X1 U1317 ( .A(\unit_decode/n2210 ), .Z(n762) );
  BUF_X1 U1318 ( .A(\unit_decode/n2209 ), .Z(n759) );
  BUF_X1 U1319 ( .A(\unit_decode/n2208 ), .Z(n756) );
  BUF_X1 U1320 ( .A(\unit_decode/n2207 ), .Z(n753) );
  BUF_X1 U1321 ( .A(\unit_decode/n2206 ), .Z(n750) );
  BUF_X1 U1322 ( .A(\unit_decode/n2205 ), .Z(n747) );
  BUF_X1 U1323 ( .A(\unit_decode/n2204 ), .Z(n744) );
  BUF_X1 U1324 ( .A(\unit_decode/n2195 ), .Z(n711) );
  BUF_X1 U1325 ( .A(\unit_decode/n2197 ), .Z(n723) );
  BUF_X1 U1326 ( .A(\unit_decode/n2198 ), .Z(n726) );
  BUF_X1 U1327 ( .A(\unit_decode/n2199 ), .Z(n729) );
  BUF_X1 U1328 ( .A(\unit_decode/n2200 ), .Z(n732) );
  BUF_X1 U1329 ( .A(\unit_decode/n2201 ), .Z(n735) );
  BUF_X1 U1330 ( .A(\unit_decode/n2202 ), .Z(n738) );
  BUF_X1 U1331 ( .A(\unit_decode/n2203 ), .Z(n741) );
  BUF_X1 U1332 ( .A(\unit_decode/n2220 ), .Z(n792) );
  BUF_X1 U1333 ( .A(\unit_decode/n2221 ), .Z(n795) );
  BUF_X1 U1334 ( .A(\unit_decode/n2222 ), .Z(n798) );
  BUF_X1 U1335 ( .A(\unit_decode/n2223 ), .Z(n801) );
  BUF_X1 U1336 ( .A(\unit_decode/n2224 ), .Z(n804) );
  BUF_X1 U1337 ( .A(\unit_decode/n2225 ), .Z(n807) );
  BUF_X1 U1338 ( .A(\unit_decode/n2226 ), .Z(n810) );
  BUF_X1 U1339 ( .A(\unit_decode/n2227 ), .Z(n813) );
  OAI22_X1 U1340 ( .A1(n977), .A2(n710), .B1(\unit_decode/n2258 ), .B2(
        \unit_decode/n1764 ), .ZN(\unit_decode/RegisterFile/n1555 ) );
  OAI22_X1 U1341 ( .A1(n977), .A2(n722), .B1(\unit_decode/n2258 ), .B2(
        \unit_decode/n1765 ), .ZN(\unit_decode/RegisterFile/n1554 ) );
  OAI22_X1 U1342 ( .A1(n977), .A2(n725), .B1(\unit_decode/n2258 ), .B2(
        \unit_decode/n1766 ), .ZN(\unit_decode/RegisterFile/n1553 ) );
  OAI22_X1 U1343 ( .A1(n968), .A2(n710), .B1(n967), .B2(\unit_decode/n1767 ), 
        .ZN(\unit_decode/RegisterFile/n1587 ) );
  OAI22_X1 U1344 ( .A1(n968), .A2(n722), .B1(n967), .B2(\unit_decode/n1768 ), 
        .ZN(\unit_decode/RegisterFile/n1586 ) );
  OAI22_X1 U1345 ( .A1(n968), .A2(n725), .B1(n967), .B2(\unit_decode/n1769 ), 
        .ZN(\unit_decode/RegisterFile/n1585 ) );
  OAI22_X1 U1346 ( .A1(n968), .A2(n728), .B1(n967), .B2(\unit_decode/n1770 ), 
        .ZN(\unit_decode/RegisterFile/n1584 ) );
  OAI22_X1 U1347 ( .A1(n968), .A2(n731), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n1771 ), .ZN(\unit_decode/RegisterFile/n1583 ) );
  OAI22_X1 U1348 ( .A1(n969), .A2(n734), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n1772 ), .ZN(\unit_decode/RegisterFile/n1582 ) );
  OAI22_X1 U1349 ( .A1(n969), .A2(n737), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n1773 ), .ZN(\unit_decode/RegisterFile/n1581 ) );
  OAI22_X1 U1350 ( .A1(n969), .A2(n740), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n1774 ), .ZN(\unit_decode/RegisterFile/n1580 ) );
  OAI22_X1 U1351 ( .A1(n941), .A2(n710), .B1(n940), .B2(\unit_decode/n1791 ), 
        .ZN(\unit_decode/RegisterFile/n1683 ) );
  OAI22_X1 U1352 ( .A1(n941), .A2(n722), .B1(n940), .B2(\unit_decode/n1792 ), 
        .ZN(\unit_decode/RegisterFile/n1682 ) );
  OAI22_X1 U1353 ( .A1(n941), .A2(n725), .B1(n940), .B2(\unit_decode/n1793 ), 
        .ZN(\unit_decode/RegisterFile/n1681 ) );
  OAI22_X1 U1354 ( .A1(n941), .A2(n728), .B1(n940), .B2(\unit_decode/n1794 ), 
        .ZN(\unit_decode/RegisterFile/n1680 ) );
  OAI22_X1 U1355 ( .A1(n941), .A2(n731), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1795 ), .ZN(\unit_decode/RegisterFile/n1679 ) );
  OAI22_X1 U1356 ( .A1(n942), .A2(n734), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1796 ), .ZN(\unit_decode/RegisterFile/n1678 ) );
  OAI22_X1 U1357 ( .A1(n942), .A2(n737), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1797 ), .ZN(\unit_decode/RegisterFile/n1677 ) );
  OAI22_X1 U1358 ( .A1(n942), .A2(n740), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1798 ), .ZN(\unit_decode/RegisterFile/n1676 ) );
  OAI22_X1 U1359 ( .A1(n932), .A2(n710), .B1(n931), .B2(\unit_decode/n1799 ), 
        .ZN(\unit_decode/RegisterFile/n1715 ) );
  OAI22_X1 U1360 ( .A1(n932), .A2(n722), .B1(n931), .B2(\unit_decode/n1800 ), 
        .ZN(\unit_decode/RegisterFile/n1714 ) );
  OAI22_X1 U1361 ( .A1(n932), .A2(n725), .B1(n931), .B2(\unit_decode/n1801 ), 
        .ZN(\unit_decode/RegisterFile/n1713 ) );
  OAI22_X1 U1362 ( .A1(n932), .A2(n728), .B1(n931), .B2(\unit_decode/n1802 ), 
        .ZN(\unit_decode/RegisterFile/n1712 ) );
  OAI22_X1 U1363 ( .A1(n932), .A2(n731), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1803 ), .ZN(\unit_decode/RegisterFile/n1711 ) );
  OAI22_X1 U1364 ( .A1(n933), .A2(n734), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1804 ), .ZN(\unit_decode/RegisterFile/n1710 ) );
  OAI22_X1 U1365 ( .A1(n933), .A2(n737), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1805 ), .ZN(\unit_decode/RegisterFile/n1709 ) );
  OAI22_X1 U1366 ( .A1(n933), .A2(n740), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1806 ), .ZN(\unit_decode/RegisterFile/n1708 ) );
  OAI22_X1 U1367 ( .A1(n905), .A2(n709), .B1(n904), .B2(\unit_decode/n1823 ), 
        .ZN(\unit_decode/RegisterFile/n1811 ) );
  OAI22_X1 U1368 ( .A1(n905), .A2(n721), .B1(n904), .B2(\unit_decode/n1824 ), 
        .ZN(\unit_decode/RegisterFile/n1810 ) );
  OAI22_X1 U1369 ( .A1(n905), .A2(n724), .B1(n904), .B2(\unit_decode/n1825 ), 
        .ZN(\unit_decode/RegisterFile/n1809 ) );
  OAI22_X1 U1370 ( .A1(n905), .A2(n727), .B1(n904), .B2(\unit_decode/n1826 ), 
        .ZN(\unit_decode/RegisterFile/n1808 ) );
  OAI22_X1 U1371 ( .A1(n905), .A2(n730), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1827 ), .ZN(\unit_decode/RegisterFile/n1807 ) );
  OAI22_X1 U1372 ( .A1(n906), .A2(n733), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1828 ), .ZN(\unit_decode/RegisterFile/n1806 ) );
  OAI22_X1 U1373 ( .A1(n906), .A2(n736), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1829 ), .ZN(\unit_decode/RegisterFile/n1805 ) );
  OAI22_X1 U1374 ( .A1(n906), .A2(n739), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1830 ), .ZN(\unit_decode/RegisterFile/n1804 ) );
  OAI22_X1 U1375 ( .A1(n896), .A2(n709), .B1(n895), .B2(\unit_decode/n1831 ), 
        .ZN(\unit_decode/RegisterFile/n1843 ) );
  OAI22_X1 U1376 ( .A1(n896), .A2(n721), .B1(n895), .B2(\unit_decode/n1832 ), 
        .ZN(\unit_decode/RegisterFile/n1842 ) );
  OAI22_X1 U1377 ( .A1(n896), .A2(n724), .B1(n895), .B2(\unit_decode/n1833 ), 
        .ZN(\unit_decode/RegisterFile/n1841 ) );
  OAI22_X1 U1378 ( .A1(n896), .A2(n727), .B1(n895), .B2(\unit_decode/n1834 ), 
        .ZN(\unit_decode/RegisterFile/n1840 ) );
  OAI22_X1 U1379 ( .A1(n896), .A2(n730), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1835 ), .ZN(\unit_decode/RegisterFile/n1839 ) );
  OAI22_X1 U1380 ( .A1(n897), .A2(n733), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1836 ), .ZN(\unit_decode/RegisterFile/n1838 ) );
  OAI22_X1 U1381 ( .A1(n897), .A2(n736), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1837 ), .ZN(\unit_decode/RegisterFile/n1837 ) );
  OAI22_X1 U1382 ( .A1(n897), .A2(n739), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1838 ), .ZN(\unit_decode/RegisterFile/n1836 ) );
  OAI22_X1 U1383 ( .A1(n1067), .A2(n711), .B1(n1066), .B2(\unit_decode/n1863 ), 
        .ZN(\unit_decode/RegisterFile/n1235 ) );
  OAI22_X1 U1384 ( .A1(n1067), .A2(n723), .B1(n1066), .B2(\unit_decode/n1864 ), 
        .ZN(\unit_decode/RegisterFile/n1234 ) );
  OAI22_X1 U1385 ( .A1(n1067), .A2(n726), .B1(n1066), .B2(\unit_decode/n1865 ), 
        .ZN(\unit_decode/RegisterFile/n1233 ) );
  OAI22_X1 U1386 ( .A1(n1067), .A2(n729), .B1(n1066), .B2(\unit_decode/n1866 ), 
        .ZN(\unit_decode/RegisterFile/n1232 ) );
  OAI22_X1 U1387 ( .A1(n1067), .A2(n732), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1867 ), .ZN(\unit_decode/RegisterFile/n1231 ) );
  OAI22_X1 U1388 ( .A1(n1068), .A2(n735), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1868 ), .ZN(\unit_decode/RegisterFile/n1230 ) );
  OAI22_X1 U1389 ( .A1(n1068), .A2(n738), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1869 ), .ZN(\unit_decode/RegisterFile/n1229 ) );
  OAI22_X1 U1390 ( .A1(n1068), .A2(n741), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1870 ), .ZN(\unit_decode/RegisterFile/n1228 ) );
  OAI22_X1 U1391 ( .A1(n869), .A2(n709), .B1(n868), .B2(\unit_decode/n1892 ), 
        .ZN(\unit_decode/RegisterFile/n1939 ) );
  OAI22_X1 U1392 ( .A1(n869), .A2(n721), .B1(n868), .B2(\unit_decode/n1893 ), 
        .ZN(\unit_decode/RegisterFile/n1938 ) );
  OAI22_X1 U1393 ( .A1(n869), .A2(n724), .B1(n868), .B2(\unit_decode/n1894 ), 
        .ZN(\unit_decode/RegisterFile/n1937 ) );
  OAI22_X1 U1394 ( .A1(n869), .A2(n727), .B1(n868), .B2(\unit_decode/n1895 ), 
        .ZN(\unit_decode/RegisterFile/n1936 ) );
  OAI22_X1 U1395 ( .A1(n869), .A2(n730), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1896 ), .ZN(\unit_decode/RegisterFile/n1935 ) );
  OAI22_X1 U1396 ( .A1(n870), .A2(n733), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1897 ), .ZN(\unit_decode/RegisterFile/n1934 ) );
  OAI22_X1 U1397 ( .A1(n870), .A2(n736), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1898 ), .ZN(\unit_decode/RegisterFile/n1933 ) );
  OAI22_X1 U1398 ( .A1(n870), .A2(n739), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1899 ), .ZN(\unit_decode/RegisterFile/n1932 ) );
  OAI22_X1 U1399 ( .A1(n860), .A2(n709), .B1(n859), .B2(\unit_decode/n1900 ), 
        .ZN(\unit_decode/RegisterFile/n1971 ) );
  OAI22_X1 U1400 ( .A1(n860), .A2(n721), .B1(n859), .B2(\unit_decode/n1901 ), 
        .ZN(\unit_decode/RegisterFile/n1970 ) );
  OAI22_X1 U1401 ( .A1(n860), .A2(n724), .B1(n859), .B2(\unit_decode/n1902 ), 
        .ZN(\unit_decode/RegisterFile/n1969 ) );
  OAI22_X1 U1402 ( .A1(n860), .A2(n727), .B1(n859), .B2(\unit_decode/n1903 ), 
        .ZN(\unit_decode/RegisterFile/n1968 ) );
  OAI22_X1 U1403 ( .A1(n860), .A2(n730), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1904 ), .ZN(\unit_decode/RegisterFile/n1967 ) );
  OAI22_X1 U1404 ( .A1(n861), .A2(n733), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1905 ), .ZN(\unit_decode/RegisterFile/n1966 ) );
  OAI22_X1 U1405 ( .A1(n861), .A2(n736), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1906 ), .ZN(\unit_decode/RegisterFile/n1965 ) );
  OAI22_X1 U1406 ( .A1(n861), .A2(n739), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1907 ), .ZN(\unit_decode/RegisterFile/n1964 ) );
  OAI22_X1 U1407 ( .A1(n833), .A2(n709), .B1(n832), .B2(\unit_decode/n1924 ), 
        .ZN(\unit_decode/RegisterFile/n2067 ) );
  OAI22_X1 U1408 ( .A1(n833), .A2(n721), .B1(n832), .B2(\unit_decode/n1925 ), 
        .ZN(\unit_decode/RegisterFile/n2066 ) );
  OAI22_X1 U1409 ( .A1(n833), .A2(n724), .B1(n832), .B2(\unit_decode/n1926 ), 
        .ZN(\unit_decode/RegisterFile/n2065 ) );
  OAI22_X1 U1410 ( .A1(n833), .A2(n727), .B1(n832), .B2(\unit_decode/n1927 ), 
        .ZN(\unit_decode/RegisterFile/n2064 ) );
  OAI22_X1 U1411 ( .A1(n833), .A2(n730), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1928 ), .ZN(\unit_decode/RegisterFile/n2063 ) );
  OAI22_X1 U1412 ( .A1(n834), .A2(n733), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1929 ), .ZN(\unit_decode/RegisterFile/n2062 ) );
  OAI22_X1 U1413 ( .A1(n834), .A2(n736), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1930 ), .ZN(\unit_decode/RegisterFile/n2061 ) );
  OAI22_X1 U1414 ( .A1(n834), .A2(n739), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1931 ), .ZN(\unit_decode/RegisterFile/n2060 ) );
  OAI22_X1 U1415 ( .A1(n824), .A2(n709), .B1(n823), .B2(\unit_decode/n1932 ), 
        .ZN(\unit_decode/RegisterFile/n2099 ) );
  OAI22_X1 U1416 ( .A1(n824), .A2(n721), .B1(n823), .B2(\unit_decode/n1933 ), 
        .ZN(\unit_decode/RegisterFile/n2098 ) );
  OAI22_X1 U1417 ( .A1(n824), .A2(n724), .B1(n823), .B2(\unit_decode/n1934 ), 
        .ZN(\unit_decode/RegisterFile/n2097 ) );
  OAI22_X1 U1418 ( .A1(n824), .A2(n727), .B1(n823), .B2(\unit_decode/n1935 ), 
        .ZN(\unit_decode/RegisterFile/n2096 ) );
  OAI22_X1 U1419 ( .A1(n824), .A2(n730), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1936 ), .ZN(\unit_decode/RegisterFile/n2095 ) );
  OAI22_X1 U1420 ( .A1(n825), .A2(n733), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1937 ), .ZN(\unit_decode/RegisterFile/n2094 ) );
  OAI22_X1 U1421 ( .A1(n825), .A2(n736), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1938 ), .ZN(\unit_decode/RegisterFile/n2093 ) );
  OAI22_X1 U1422 ( .A1(n825), .A2(n739), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1939 ), .ZN(\unit_decode/RegisterFile/n2092 ) );
  OAI22_X1 U1423 ( .A1(n1064), .A2(n813), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1245 ), .ZN(\unit_decode/RegisterFile/n1236 ) );
  OAI22_X1 U1424 ( .A1(n1064), .A2(n810), .B1(n1057), .B2(\unit_decode/n1246 ), 
        .ZN(\unit_decode/RegisterFile/n1237 ) );
  OAI22_X1 U1425 ( .A1(n1063), .A2(n807), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1247 ), .ZN(\unit_decode/RegisterFile/n1238 ) );
  OAI22_X1 U1426 ( .A1(n1063), .A2(n804), .B1(n1057), .B2(\unit_decode/n1248 ), 
        .ZN(\unit_decode/RegisterFile/n1239 ) );
  OAI22_X1 U1427 ( .A1(n1063), .A2(n801), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1249 ), .ZN(\unit_decode/RegisterFile/n1240 ) );
  OAI22_X1 U1428 ( .A1(n1063), .A2(n798), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1250 ), .ZN(\unit_decode/RegisterFile/n1241 ) );
  OAI22_X1 U1429 ( .A1(n1063), .A2(n795), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1251 ), .ZN(\unit_decode/RegisterFile/n1242 ) );
  OAI22_X1 U1430 ( .A1(n1055), .A2(n813), .B1(\unit_decode/n2267 ), .B2(
        \unit_decode/n1269 ), .ZN(\unit_decode/RegisterFile/n1268 ) );
  OAI22_X1 U1431 ( .A1(n1055), .A2(n810), .B1(n1048), .B2(\unit_decode/n1270 ), 
        .ZN(\unit_decode/RegisterFile/n1269 ) );
  OAI22_X1 U1432 ( .A1(n1054), .A2(n807), .B1(\unit_decode/n2267 ), .B2(
        \unit_decode/n1271 ), .ZN(\unit_decode/RegisterFile/n1270 ) );
  OAI22_X1 U1433 ( .A1(n1054), .A2(n804), .B1(n1048), .B2(\unit_decode/n1272 ), 
        .ZN(\unit_decode/RegisterFile/n1271 ) );
  OAI22_X1 U1434 ( .A1(n1054), .A2(n801), .B1(\unit_decode/n2267 ), .B2(
        \unit_decode/n1273 ), .ZN(\unit_decode/RegisterFile/n1272 ) );
  OAI22_X1 U1435 ( .A1(n1054), .A2(n798), .B1(\unit_decode/n2267 ), .B2(
        \unit_decode/n1274 ), .ZN(\unit_decode/RegisterFile/n1273 ) );
  OAI22_X1 U1436 ( .A1(n1054), .A2(n795), .B1(\unit_decode/n2267 ), .B2(
        \unit_decode/n1275 ), .ZN(\unit_decode/RegisterFile/n1274 ) );
  OAI22_X1 U1437 ( .A1(n1046), .A2(n813), .B1(\unit_decode/n2266 ), .B2(
        \unit_decode/n1293 ), .ZN(\unit_decode/RegisterFile/n1300 ) );
  OAI22_X1 U1438 ( .A1(n1046), .A2(n810), .B1(n1039), .B2(\unit_decode/n1294 ), 
        .ZN(\unit_decode/RegisterFile/n1301 ) );
  OAI22_X1 U1439 ( .A1(n1045), .A2(n807), .B1(\unit_decode/n2266 ), .B2(
        \unit_decode/n1295 ), .ZN(\unit_decode/RegisterFile/n1302 ) );
  OAI22_X1 U1440 ( .A1(n1045), .A2(n804), .B1(n1039), .B2(\unit_decode/n1296 ), 
        .ZN(\unit_decode/RegisterFile/n1303 ) );
  OAI22_X1 U1441 ( .A1(n1045), .A2(n801), .B1(\unit_decode/n2266 ), .B2(
        \unit_decode/n1297 ), .ZN(\unit_decode/RegisterFile/n1304 ) );
  OAI22_X1 U1442 ( .A1(n1045), .A2(n798), .B1(\unit_decode/n2266 ), .B2(
        \unit_decode/n1298 ), .ZN(\unit_decode/RegisterFile/n1305 ) );
  OAI22_X1 U1443 ( .A1(n1045), .A2(n795), .B1(\unit_decode/n2266 ), .B2(
        \unit_decode/n1299 ), .ZN(\unit_decode/RegisterFile/n1306 ) );
  OAI22_X1 U1444 ( .A1(n1062), .A2(n792), .B1(n1057), .B2(\unit_decode/n1252 ), 
        .ZN(\unit_decode/RegisterFile/n1243 ) );
  OAI22_X1 U1445 ( .A1(n1062), .A2(n789), .B1(n1057), .B2(\unit_decode/n1253 ), 
        .ZN(\unit_decode/RegisterFile/n1244 ) );
  OAI22_X1 U1446 ( .A1(n1062), .A2(n786), .B1(n1057), .B2(\unit_decode/n1254 ), 
        .ZN(\unit_decode/RegisterFile/n1245 ) );
  OAI22_X1 U1447 ( .A1(n1062), .A2(n783), .B1(n1057), .B2(\unit_decode/n1255 ), 
        .ZN(\unit_decode/RegisterFile/n1246 ) );
  OAI22_X1 U1448 ( .A1(n1062), .A2(n780), .B1(n1057), .B2(\unit_decode/n1256 ), 
        .ZN(\unit_decode/RegisterFile/n1247 ) );
  OAI22_X1 U1449 ( .A1(n1061), .A2(n777), .B1(n1057), .B2(\unit_decode/n1257 ), 
        .ZN(\unit_decode/RegisterFile/n1248 ) );
  OAI22_X1 U1450 ( .A1(n1061), .A2(n774), .B1(n1057), .B2(\unit_decode/n1258 ), 
        .ZN(\unit_decode/RegisterFile/n1249 ) );
  OAI22_X1 U1451 ( .A1(n1061), .A2(n771), .B1(n1057), .B2(\unit_decode/n1259 ), 
        .ZN(\unit_decode/RegisterFile/n1250 ) );
  OAI22_X1 U1452 ( .A1(n1061), .A2(n768), .B1(n1057), .B2(\unit_decode/n1260 ), 
        .ZN(\unit_decode/RegisterFile/n1251 ) );
  OAI22_X1 U1453 ( .A1(n1061), .A2(n765), .B1(n1057), .B2(\unit_decode/n1261 ), 
        .ZN(\unit_decode/RegisterFile/n1252 ) );
  OAI22_X1 U1454 ( .A1(n1060), .A2(n762), .B1(n1057), .B2(\unit_decode/n1262 ), 
        .ZN(\unit_decode/RegisterFile/n1253 ) );
  OAI22_X1 U1455 ( .A1(n1060), .A2(n759), .B1(n1057), .B2(\unit_decode/n1263 ), 
        .ZN(\unit_decode/RegisterFile/n1254 ) );
  OAI22_X1 U1456 ( .A1(n1060), .A2(n756), .B1(n1057), .B2(\unit_decode/n1264 ), 
        .ZN(\unit_decode/RegisterFile/n1255 ) );
  OAI22_X1 U1457 ( .A1(n1053), .A2(n792), .B1(n1048), .B2(\unit_decode/n1276 ), 
        .ZN(\unit_decode/RegisterFile/n1275 ) );
  OAI22_X1 U1458 ( .A1(n1053), .A2(n789), .B1(n1048), .B2(\unit_decode/n1277 ), 
        .ZN(\unit_decode/RegisterFile/n1276 ) );
  OAI22_X1 U1459 ( .A1(n1053), .A2(n786), .B1(n1048), .B2(\unit_decode/n1278 ), 
        .ZN(\unit_decode/RegisterFile/n1277 ) );
  OAI22_X1 U1460 ( .A1(n1053), .A2(n783), .B1(n1048), .B2(\unit_decode/n1279 ), 
        .ZN(\unit_decode/RegisterFile/n1278 ) );
  OAI22_X1 U1461 ( .A1(n1053), .A2(n780), .B1(n1048), .B2(\unit_decode/n1280 ), 
        .ZN(\unit_decode/RegisterFile/n1279 ) );
  OAI22_X1 U1462 ( .A1(n1052), .A2(n777), .B1(n1048), .B2(\unit_decode/n1281 ), 
        .ZN(\unit_decode/RegisterFile/n1280 ) );
  OAI22_X1 U1463 ( .A1(n1052), .A2(n774), .B1(n1048), .B2(\unit_decode/n1282 ), 
        .ZN(\unit_decode/RegisterFile/n1281 ) );
  OAI22_X1 U1464 ( .A1(n1052), .A2(n771), .B1(n1048), .B2(\unit_decode/n1283 ), 
        .ZN(\unit_decode/RegisterFile/n1282 ) );
  OAI22_X1 U1465 ( .A1(n1052), .A2(n768), .B1(n1048), .B2(\unit_decode/n1284 ), 
        .ZN(\unit_decode/RegisterFile/n1283 ) );
  OAI22_X1 U1466 ( .A1(n1052), .A2(n765), .B1(n1048), .B2(\unit_decode/n1285 ), 
        .ZN(\unit_decode/RegisterFile/n1284 ) );
  OAI22_X1 U1467 ( .A1(n1051), .A2(n762), .B1(n1048), .B2(\unit_decode/n1286 ), 
        .ZN(\unit_decode/RegisterFile/n1285 ) );
  OAI22_X1 U1468 ( .A1(n1051), .A2(n759), .B1(n1048), .B2(\unit_decode/n1287 ), 
        .ZN(\unit_decode/RegisterFile/n1286 ) );
  OAI22_X1 U1469 ( .A1(n1051), .A2(n756), .B1(n1048), .B2(\unit_decode/n1288 ), 
        .ZN(\unit_decode/RegisterFile/n1287 ) );
  OAI22_X1 U1470 ( .A1(n1044), .A2(n792), .B1(n1039), .B2(\unit_decode/n1300 ), 
        .ZN(\unit_decode/RegisterFile/n1307 ) );
  OAI22_X1 U1471 ( .A1(n1044), .A2(n789), .B1(n1039), .B2(\unit_decode/n1301 ), 
        .ZN(\unit_decode/RegisterFile/n1308 ) );
  OAI22_X1 U1472 ( .A1(n1044), .A2(n786), .B1(n1039), .B2(\unit_decode/n1302 ), 
        .ZN(\unit_decode/RegisterFile/n1309 ) );
  OAI22_X1 U1473 ( .A1(n1044), .A2(n783), .B1(n1039), .B2(\unit_decode/n1303 ), 
        .ZN(\unit_decode/RegisterFile/n1310 ) );
  OAI22_X1 U1474 ( .A1(n1044), .A2(n780), .B1(n1039), .B2(\unit_decode/n1304 ), 
        .ZN(\unit_decode/RegisterFile/n1311 ) );
  OAI22_X1 U1475 ( .A1(n1043), .A2(n777), .B1(n1039), .B2(\unit_decode/n1305 ), 
        .ZN(\unit_decode/RegisterFile/n1312 ) );
  OAI22_X1 U1476 ( .A1(n1043), .A2(n774), .B1(n1039), .B2(\unit_decode/n1306 ), 
        .ZN(\unit_decode/RegisterFile/n1313 ) );
  OAI22_X1 U1477 ( .A1(n1043), .A2(n771), .B1(n1039), .B2(\unit_decode/n1307 ), 
        .ZN(\unit_decode/RegisterFile/n1314 ) );
  OAI22_X1 U1478 ( .A1(n1043), .A2(n768), .B1(n1039), .B2(\unit_decode/n1308 ), 
        .ZN(\unit_decode/RegisterFile/n1315 ) );
  OAI22_X1 U1479 ( .A1(n1043), .A2(n765), .B1(n1039), .B2(\unit_decode/n1309 ), 
        .ZN(\unit_decode/RegisterFile/n1316 ) );
  OAI22_X1 U1480 ( .A1(n1042), .A2(n762), .B1(n1039), .B2(\unit_decode/n1310 ), 
        .ZN(\unit_decode/RegisterFile/n1317 ) );
  OAI22_X1 U1481 ( .A1(n1042), .A2(n759), .B1(n1039), .B2(\unit_decode/n1311 ), 
        .ZN(\unit_decode/RegisterFile/n1318 ) );
  OAI22_X1 U1482 ( .A1(n1042), .A2(n756), .B1(n1039), .B2(\unit_decode/n1312 ), 
        .ZN(\unit_decode/RegisterFile/n1319 ) );
  OAI22_X1 U1483 ( .A1(n1051), .A2(n753), .B1(n1048), .B2(\unit_decode/n1289 ), 
        .ZN(\unit_decode/RegisterFile/n1288 ) );
  OAI22_X1 U1484 ( .A1(n1051), .A2(n750), .B1(n1048), .B2(\unit_decode/n1290 ), 
        .ZN(\unit_decode/RegisterFile/n1289 ) );
  OAI22_X1 U1485 ( .A1(n1050), .A2(n747), .B1(n1048), .B2(\unit_decode/n1291 ), 
        .ZN(\unit_decode/RegisterFile/n1290 ) );
  OAI22_X1 U1486 ( .A1(n1050), .A2(n744), .B1(n1048), .B2(\unit_decode/n1292 ), 
        .ZN(\unit_decode/RegisterFile/n1291 ) );
  OAI22_X1 U1487 ( .A1(n1042), .A2(n753), .B1(n1039), .B2(\unit_decode/n1313 ), 
        .ZN(\unit_decode/RegisterFile/n1320 ) );
  OAI22_X1 U1488 ( .A1(n1042), .A2(n750), .B1(n1039), .B2(\unit_decode/n1314 ), 
        .ZN(\unit_decode/RegisterFile/n1321 ) );
  OAI22_X1 U1489 ( .A1(n1041), .A2(n747), .B1(n1039), .B2(\unit_decode/n1315 ), 
        .ZN(\unit_decode/RegisterFile/n1322 ) );
  OAI22_X1 U1490 ( .A1(n1041), .A2(n744), .B1(n1039), .B2(\unit_decode/n1316 ), 
        .ZN(\unit_decode/RegisterFile/n1323 ) );
  OAI22_X1 U1491 ( .A1(n1060), .A2(n753), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1265 ), .ZN(\unit_decode/RegisterFile/n1256 ) );
  OAI22_X1 U1492 ( .A1(n1060), .A2(n750), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1266 ), .ZN(\unit_decode/RegisterFile/n1257 ) );
  OAI22_X1 U1493 ( .A1(n1059), .A2(n747), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1267 ), .ZN(\unit_decode/RegisterFile/n1258 ) );
  OAI22_X1 U1494 ( .A1(n1059), .A2(n744), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1268 ), .ZN(\unit_decode/RegisterFile/n1259 ) );
  OAI22_X1 U1495 ( .A1(n1058), .A2(n729), .B1(\unit_decode/n2268 ), .B2(
        \unit_decode/n1871 ), .ZN(\unit_decode/RegisterFile/n1264 ) );
  OAI22_X1 U1496 ( .A1(n1058), .A2(n732), .B1(n1057), .B2(\unit_decode/n1872 ), 
        .ZN(\unit_decode/RegisterFile/n1263 ) );
  OAI22_X1 U1497 ( .A1(n1059), .A2(n735), .B1(n1057), .B2(\unit_decode/n1873 ), 
        .ZN(\unit_decode/RegisterFile/n1262 ) );
  OAI22_X1 U1498 ( .A1(n1059), .A2(n738), .B1(n1057), .B2(\unit_decode/n1874 ), 
        .ZN(\unit_decode/RegisterFile/n1261 ) );
  OAI22_X1 U1499 ( .A1(n1059), .A2(n741), .B1(n1057), .B2(\unit_decode/n1875 ), 
        .ZN(\unit_decode/RegisterFile/n1260 ) );
  OAI22_X1 U1500 ( .A1(n1073), .A2(n813), .B1(n1066), .B2(\unit_decode/n1221 ), 
        .ZN(\unit_decode/RegisterFile/n1204 ) );
  OAI22_X1 U1501 ( .A1(n1073), .A2(n810), .B1(n1066), .B2(\unit_decode/n1222 ), 
        .ZN(\unit_decode/RegisterFile/n1205 ) );
  OAI22_X1 U1502 ( .A1(n1072), .A2(n807), .B1(n1066), .B2(\unit_decode/n1223 ), 
        .ZN(\unit_decode/RegisterFile/n1206 ) );
  OAI22_X1 U1503 ( .A1(n1072), .A2(n804), .B1(n1066), .B2(\unit_decode/n1224 ), 
        .ZN(\unit_decode/RegisterFile/n1207 ) );
  OAI22_X1 U1504 ( .A1(n1072), .A2(n801), .B1(n1066), .B2(\unit_decode/n1225 ), 
        .ZN(\unit_decode/RegisterFile/n1208 ) );
  OAI22_X1 U1505 ( .A1(n1072), .A2(n798), .B1(n1066), .B2(\unit_decode/n1226 ), 
        .ZN(\unit_decode/RegisterFile/n1209 ) );
  OAI22_X1 U1506 ( .A1(n1072), .A2(n795), .B1(n1066), .B2(\unit_decode/n1227 ), 
        .ZN(\unit_decode/RegisterFile/n1210 ) );
  OAI22_X1 U1507 ( .A1(n1071), .A2(n792), .B1(n1066), .B2(\unit_decode/n1228 ), 
        .ZN(\unit_decode/RegisterFile/n1211 ) );
  OAI22_X1 U1508 ( .A1(n1071), .A2(n789), .B1(n1066), .B2(\unit_decode/n1229 ), 
        .ZN(\unit_decode/RegisterFile/n1212 ) );
  OAI22_X1 U1509 ( .A1(n1071), .A2(n786), .B1(n1066), .B2(\unit_decode/n1230 ), 
        .ZN(\unit_decode/RegisterFile/n1213 ) );
  OAI22_X1 U1510 ( .A1(n1071), .A2(n783), .B1(n1066), .B2(\unit_decode/n1231 ), 
        .ZN(\unit_decode/RegisterFile/n1214 ) );
  OAI22_X1 U1511 ( .A1(n1071), .A2(n780), .B1(n1066), .B2(\unit_decode/n1232 ), 
        .ZN(\unit_decode/RegisterFile/n1215 ) );
  OAI22_X1 U1512 ( .A1(n1070), .A2(n777), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1233 ), .ZN(\unit_decode/RegisterFile/n1216 ) );
  OAI22_X1 U1513 ( .A1(n1070), .A2(n774), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1234 ), .ZN(\unit_decode/RegisterFile/n1217 ) );
  OAI22_X1 U1514 ( .A1(n1070), .A2(n771), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1235 ), .ZN(\unit_decode/RegisterFile/n1218 ) );
  OAI22_X1 U1515 ( .A1(n1070), .A2(n768), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1236 ), .ZN(\unit_decode/RegisterFile/n1219 ) );
  OAI22_X1 U1516 ( .A1(n1070), .A2(n765), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1237 ), .ZN(\unit_decode/RegisterFile/n1220 ) );
  OAI22_X1 U1517 ( .A1(n1069), .A2(n762), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1238 ), .ZN(\unit_decode/RegisterFile/n1221 ) );
  OAI22_X1 U1518 ( .A1(n1069), .A2(n759), .B1(\unit_decode/n2269 ), .B2(
        \unit_decode/n1239 ), .ZN(\unit_decode/RegisterFile/n1222 ) );
  OAI22_X1 U1519 ( .A1(n1069), .A2(n756), .B1(n1066), .B2(\unit_decode/n1240 ), 
        .ZN(\unit_decode/RegisterFile/n1223 ) );
  OAI22_X1 U1520 ( .A1(n1069), .A2(n753), .B1(n1066), .B2(\unit_decode/n1241 ), 
        .ZN(\unit_decode/RegisterFile/n1224 ) );
  OAI22_X1 U1521 ( .A1(n1069), .A2(n750), .B1(n1066), .B2(\unit_decode/n1242 ), 
        .ZN(\unit_decode/RegisterFile/n1225 ) );
  OAI22_X1 U1522 ( .A1(n1068), .A2(n747), .B1(n1066), .B2(\unit_decode/n1243 ), 
        .ZN(\unit_decode/RegisterFile/n1226 ) );
  OAI22_X1 U1523 ( .A1(n1068), .A2(n744), .B1(n1066), .B2(\unit_decode/n1244 ), 
        .ZN(\unit_decode/RegisterFile/n1227 ) );
  OAI22_X1 U1524 ( .A1(n947), .A2(n812), .B1(n940), .B2(\unit_decode/n1365 ), 
        .ZN(\unit_decode/RegisterFile/n1652 ) );
  OAI22_X1 U1525 ( .A1(n947), .A2(n809), .B1(n940), .B2(\unit_decode/n1366 ), 
        .ZN(\unit_decode/RegisterFile/n1653 ) );
  OAI22_X1 U1526 ( .A1(n946), .A2(n806), .B1(n940), .B2(\unit_decode/n1367 ), 
        .ZN(\unit_decode/RegisterFile/n1654 ) );
  OAI22_X1 U1527 ( .A1(n946), .A2(n803), .B1(n940), .B2(\unit_decode/n1368 ), 
        .ZN(\unit_decode/RegisterFile/n1655 ) );
  OAI22_X1 U1528 ( .A1(n946), .A2(n800), .B1(n940), .B2(\unit_decode/n1369 ), 
        .ZN(\unit_decode/RegisterFile/n1656 ) );
  OAI22_X1 U1529 ( .A1(n946), .A2(n797), .B1(n940), .B2(\unit_decode/n1370 ), 
        .ZN(\unit_decode/RegisterFile/n1657 ) );
  OAI22_X1 U1530 ( .A1(n946), .A2(n794), .B1(n940), .B2(\unit_decode/n1371 ), 
        .ZN(\unit_decode/RegisterFile/n1658 ) );
  OAI22_X1 U1531 ( .A1(n945), .A2(n791), .B1(n940), .B2(\unit_decode/n1372 ), 
        .ZN(\unit_decode/RegisterFile/n1659 ) );
  OAI22_X1 U1532 ( .A1(n945), .A2(n788), .B1(n940), .B2(\unit_decode/n1373 ), 
        .ZN(\unit_decode/RegisterFile/n1660 ) );
  OAI22_X1 U1533 ( .A1(n945), .A2(n785), .B1(n940), .B2(\unit_decode/n1374 ), 
        .ZN(\unit_decode/RegisterFile/n1661 ) );
  OAI22_X1 U1534 ( .A1(n945), .A2(n782), .B1(n940), .B2(\unit_decode/n1375 ), 
        .ZN(\unit_decode/RegisterFile/n1662 ) );
  OAI22_X1 U1535 ( .A1(n945), .A2(n779), .B1(n940), .B2(\unit_decode/n1376 ), 
        .ZN(\unit_decode/RegisterFile/n1663 ) );
  OAI22_X1 U1536 ( .A1(n944), .A2(n776), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1377 ), .ZN(\unit_decode/RegisterFile/n1664 ) );
  OAI22_X1 U1537 ( .A1(n944), .A2(n773), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1378 ), .ZN(\unit_decode/RegisterFile/n1665 ) );
  OAI22_X1 U1538 ( .A1(n944), .A2(n770), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1379 ), .ZN(\unit_decode/RegisterFile/n1666 ) );
  OAI22_X1 U1539 ( .A1(n944), .A2(n767), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1380 ), .ZN(\unit_decode/RegisterFile/n1667 ) );
  OAI22_X1 U1540 ( .A1(n944), .A2(n764), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1381 ), .ZN(\unit_decode/RegisterFile/n1668 ) );
  OAI22_X1 U1541 ( .A1(n943), .A2(n761), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1382 ), .ZN(\unit_decode/RegisterFile/n1669 ) );
  OAI22_X1 U1542 ( .A1(n943), .A2(n758), .B1(\unit_decode/n2253 ), .B2(
        \unit_decode/n1383 ), .ZN(\unit_decode/RegisterFile/n1670 ) );
  OAI22_X1 U1543 ( .A1(n943), .A2(n755), .B1(n940), .B2(\unit_decode/n1384 ), 
        .ZN(\unit_decode/RegisterFile/n1671 ) );
  OAI22_X1 U1544 ( .A1(n943), .A2(n752), .B1(n940), .B2(\unit_decode/n1385 ), 
        .ZN(\unit_decode/RegisterFile/n1672 ) );
  OAI22_X1 U1545 ( .A1(n943), .A2(n749), .B1(n940), .B2(\unit_decode/n1386 ), 
        .ZN(\unit_decode/RegisterFile/n1673 ) );
  OAI22_X1 U1546 ( .A1(n942), .A2(n746), .B1(n940), .B2(\unit_decode/n1387 ), 
        .ZN(\unit_decode/RegisterFile/n1674 ) );
  OAI22_X1 U1547 ( .A1(n938), .A2(n812), .B1(n931), .B2(\unit_decode/n1388 ), 
        .ZN(\unit_decode/RegisterFile/n1684 ) );
  OAI22_X1 U1548 ( .A1(n938), .A2(n809), .B1(n931), .B2(\unit_decode/n1389 ), 
        .ZN(\unit_decode/RegisterFile/n1685 ) );
  OAI22_X1 U1549 ( .A1(n937), .A2(n806), .B1(n931), .B2(\unit_decode/n1390 ), 
        .ZN(\unit_decode/RegisterFile/n1686 ) );
  OAI22_X1 U1550 ( .A1(n937), .A2(n803), .B1(n931), .B2(\unit_decode/n1391 ), 
        .ZN(\unit_decode/RegisterFile/n1687 ) );
  OAI22_X1 U1551 ( .A1(n937), .A2(n800), .B1(n931), .B2(\unit_decode/n1392 ), 
        .ZN(\unit_decode/RegisterFile/n1688 ) );
  OAI22_X1 U1552 ( .A1(n937), .A2(n797), .B1(n931), .B2(\unit_decode/n1393 ), 
        .ZN(\unit_decode/RegisterFile/n1689 ) );
  OAI22_X1 U1553 ( .A1(n937), .A2(n794), .B1(n931), .B2(\unit_decode/n1394 ), 
        .ZN(\unit_decode/RegisterFile/n1690 ) );
  OAI22_X1 U1554 ( .A1(n936), .A2(n791), .B1(n931), .B2(\unit_decode/n1395 ), 
        .ZN(\unit_decode/RegisterFile/n1691 ) );
  OAI22_X1 U1555 ( .A1(n936), .A2(n788), .B1(n931), .B2(\unit_decode/n1396 ), 
        .ZN(\unit_decode/RegisterFile/n1692 ) );
  OAI22_X1 U1556 ( .A1(n936), .A2(n785), .B1(n931), .B2(\unit_decode/n1397 ), 
        .ZN(\unit_decode/RegisterFile/n1693 ) );
  OAI22_X1 U1557 ( .A1(n936), .A2(n782), .B1(n931), .B2(\unit_decode/n1398 ), 
        .ZN(\unit_decode/RegisterFile/n1694 ) );
  OAI22_X1 U1558 ( .A1(n936), .A2(n779), .B1(n931), .B2(\unit_decode/n1399 ), 
        .ZN(\unit_decode/RegisterFile/n1695 ) );
  OAI22_X1 U1559 ( .A1(n935), .A2(n776), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1400 ), .ZN(\unit_decode/RegisterFile/n1696 ) );
  OAI22_X1 U1560 ( .A1(n935), .A2(n773), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1401 ), .ZN(\unit_decode/RegisterFile/n1697 ) );
  OAI22_X1 U1561 ( .A1(n935), .A2(n770), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1402 ), .ZN(\unit_decode/RegisterFile/n1698 ) );
  OAI22_X1 U1562 ( .A1(n935), .A2(n767), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1403 ), .ZN(\unit_decode/RegisterFile/n1699 ) );
  OAI22_X1 U1563 ( .A1(n935), .A2(n764), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1404 ), .ZN(\unit_decode/RegisterFile/n1700 ) );
  OAI22_X1 U1564 ( .A1(n934), .A2(n761), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1405 ), .ZN(\unit_decode/RegisterFile/n1701 ) );
  OAI22_X1 U1565 ( .A1(n934), .A2(n758), .B1(\unit_decode/n2252 ), .B2(
        \unit_decode/n1406 ), .ZN(\unit_decode/RegisterFile/n1702 ) );
  OAI22_X1 U1566 ( .A1(n934), .A2(n755), .B1(n931), .B2(\unit_decode/n1407 ), 
        .ZN(\unit_decode/RegisterFile/n1703 ) );
  OAI22_X1 U1567 ( .A1(n934), .A2(n752), .B1(n931), .B2(\unit_decode/n1408 ), 
        .ZN(\unit_decode/RegisterFile/n1704 ) );
  OAI22_X1 U1568 ( .A1(n934), .A2(n749), .B1(n931), .B2(\unit_decode/n1409 ), 
        .ZN(\unit_decode/RegisterFile/n1705 ) );
  OAI22_X1 U1569 ( .A1(n933), .A2(n746), .B1(n931), .B2(\unit_decode/n1410 ), 
        .ZN(\unit_decode/RegisterFile/n1706 ) );
  OAI22_X1 U1570 ( .A1(n933), .A2(n743), .B1(n931), .B2(\unit_decode/n1411 ), 
        .ZN(\unit_decode/RegisterFile/n1707 ) );
  OAI22_X1 U1571 ( .A1(n911), .A2(n811), .B1(n904), .B2(\unit_decode/n1460 ), 
        .ZN(\unit_decode/RegisterFile/n1780 ) );
  OAI22_X1 U1572 ( .A1(n911), .A2(n808), .B1(n904), .B2(\unit_decode/n1461 ), 
        .ZN(\unit_decode/RegisterFile/n1781 ) );
  OAI22_X1 U1573 ( .A1(n910), .A2(n805), .B1(n904), .B2(\unit_decode/n1462 ), 
        .ZN(\unit_decode/RegisterFile/n1782 ) );
  OAI22_X1 U1574 ( .A1(n910), .A2(n802), .B1(n904), .B2(\unit_decode/n1463 ), 
        .ZN(\unit_decode/RegisterFile/n1783 ) );
  OAI22_X1 U1575 ( .A1(n910), .A2(n799), .B1(n904), .B2(\unit_decode/n1464 ), 
        .ZN(\unit_decode/RegisterFile/n1784 ) );
  OAI22_X1 U1576 ( .A1(n910), .A2(n796), .B1(n904), .B2(\unit_decode/n1465 ), 
        .ZN(\unit_decode/RegisterFile/n1785 ) );
  OAI22_X1 U1577 ( .A1(n910), .A2(n793), .B1(n904), .B2(\unit_decode/n1466 ), 
        .ZN(\unit_decode/RegisterFile/n1786 ) );
  OAI22_X1 U1578 ( .A1(n909), .A2(n790), .B1(n904), .B2(\unit_decode/n1467 ), 
        .ZN(\unit_decode/RegisterFile/n1787 ) );
  OAI22_X1 U1579 ( .A1(n909), .A2(n787), .B1(n904), .B2(\unit_decode/n1468 ), 
        .ZN(\unit_decode/RegisterFile/n1788 ) );
  OAI22_X1 U1580 ( .A1(n909), .A2(n784), .B1(n904), .B2(\unit_decode/n1469 ), 
        .ZN(\unit_decode/RegisterFile/n1789 ) );
  OAI22_X1 U1581 ( .A1(n909), .A2(n781), .B1(n904), .B2(\unit_decode/n1470 ), 
        .ZN(\unit_decode/RegisterFile/n1790 ) );
  OAI22_X1 U1582 ( .A1(n909), .A2(n778), .B1(n904), .B2(\unit_decode/n1471 ), 
        .ZN(\unit_decode/RegisterFile/n1791 ) );
  OAI22_X1 U1583 ( .A1(n908), .A2(n775), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1472 ), .ZN(\unit_decode/RegisterFile/n1792 ) );
  OAI22_X1 U1584 ( .A1(n908), .A2(n772), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1473 ), .ZN(\unit_decode/RegisterFile/n1793 ) );
  OAI22_X1 U1585 ( .A1(n908), .A2(n769), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1474 ), .ZN(\unit_decode/RegisterFile/n1794 ) );
  OAI22_X1 U1586 ( .A1(n908), .A2(n766), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1475 ), .ZN(\unit_decode/RegisterFile/n1795 ) );
  OAI22_X1 U1587 ( .A1(n908), .A2(n763), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1476 ), .ZN(\unit_decode/RegisterFile/n1796 ) );
  OAI22_X1 U1588 ( .A1(n907), .A2(n760), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1477 ), .ZN(\unit_decode/RegisterFile/n1797 ) );
  OAI22_X1 U1589 ( .A1(n907), .A2(n757), .B1(\unit_decode/n2249 ), .B2(
        \unit_decode/n1478 ), .ZN(\unit_decode/RegisterFile/n1798 ) );
  OAI22_X1 U1590 ( .A1(n907), .A2(n754), .B1(n904), .B2(\unit_decode/n1479 ), 
        .ZN(\unit_decode/RegisterFile/n1799 ) );
  OAI22_X1 U1591 ( .A1(n907), .A2(n751), .B1(n904), .B2(\unit_decode/n1480 ), 
        .ZN(\unit_decode/RegisterFile/n1800 ) );
  OAI22_X1 U1592 ( .A1(n907), .A2(n748), .B1(n904), .B2(\unit_decode/n1481 ), 
        .ZN(\unit_decode/RegisterFile/n1801 ) );
  OAI22_X1 U1593 ( .A1(n906), .A2(n745), .B1(n904), .B2(\unit_decode/n1482 ), 
        .ZN(\unit_decode/RegisterFile/n1802 ) );
  OAI22_X1 U1594 ( .A1(n906), .A2(n742), .B1(n904), .B2(\unit_decode/n1483 ), 
        .ZN(\unit_decode/RegisterFile/n1803 ) );
  OAI22_X1 U1595 ( .A1(n902), .A2(n811), .B1(n895), .B2(\unit_decode/n1484 ), 
        .ZN(\unit_decode/RegisterFile/n1812 ) );
  OAI22_X1 U1596 ( .A1(n902), .A2(n808), .B1(n895), .B2(\unit_decode/n1485 ), 
        .ZN(\unit_decode/RegisterFile/n1813 ) );
  OAI22_X1 U1597 ( .A1(n901), .A2(n805), .B1(n895), .B2(\unit_decode/n1486 ), 
        .ZN(\unit_decode/RegisterFile/n1814 ) );
  OAI22_X1 U1598 ( .A1(n901), .A2(n802), .B1(n895), .B2(\unit_decode/n1487 ), 
        .ZN(\unit_decode/RegisterFile/n1815 ) );
  OAI22_X1 U1599 ( .A1(n901), .A2(n799), .B1(n895), .B2(\unit_decode/n1488 ), 
        .ZN(\unit_decode/RegisterFile/n1816 ) );
  OAI22_X1 U1600 ( .A1(n901), .A2(n796), .B1(n895), .B2(\unit_decode/n1489 ), 
        .ZN(\unit_decode/RegisterFile/n1817 ) );
  OAI22_X1 U1601 ( .A1(n901), .A2(n793), .B1(n895), .B2(\unit_decode/n1490 ), 
        .ZN(\unit_decode/RegisterFile/n1818 ) );
  OAI22_X1 U1602 ( .A1(n900), .A2(n790), .B1(n895), .B2(\unit_decode/n1491 ), 
        .ZN(\unit_decode/RegisterFile/n1819 ) );
  OAI22_X1 U1603 ( .A1(n900), .A2(n787), .B1(n895), .B2(\unit_decode/n1492 ), 
        .ZN(\unit_decode/RegisterFile/n1820 ) );
  OAI22_X1 U1604 ( .A1(n900), .A2(n784), .B1(n895), .B2(\unit_decode/n1493 ), 
        .ZN(\unit_decode/RegisterFile/n1821 ) );
  OAI22_X1 U1605 ( .A1(n900), .A2(n781), .B1(n895), .B2(\unit_decode/n1494 ), 
        .ZN(\unit_decode/RegisterFile/n1822 ) );
  OAI22_X1 U1606 ( .A1(n900), .A2(n778), .B1(n895), .B2(\unit_decode/n1495 ), 
        .ZN(\unit_decode/RegisterFile/n1823 ) );
  OAI22_X1 U1607 ( .A1(n899), .A2(n775), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1496 ), .ZN(\unit_decode/RegisterFile/n1824 ) );
  OAI22_X1 U1608 ( .A1(n899), .A2(n772), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1497 ), .ZN(\unit_decode/RegisterFile/n1825 ) );
  OAI22_X1 U1609 ( .A1(n899), .A2(n769), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1498 ), .ZN(\unit_decode/RegisterFile/n1826 ) );
  OAI22_X1 U1610 ( .A1(n899), .A2(n766), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1499 ), .ZN(\unit_decode/RegisterFile/n1827 ) );
  OAI22_X1 U1611 ( .A1(n899), .A2(n763), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1500 ), .ZN(\unit_decode/RegisterFile/n1828 ) );
  OAI22_X1 U1612 ( .A1(n898), .A2(n760), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1501 ), .ZN(\unit_decode/RegisterFile/n1829 ) );
  OAI22_X1 U1613 ( .A1(n898), .A2(n757), .B1(\unit_decode/n2248 ), .B2(
        \unit_decode/n1502 ), .ZN(\unit_decode/RegisterFile/n1830 ) );
  OAI22_X1 U1614 ( .A1(n898), .A2(n754), .B1(n895), .B2(\unit_decode/n1503 ), 
        .ZN(\unit_decode/RegisterFile/n1831 ) );
  OAI22_X1 U1615 ( .A1(n898), .A2(n751), .B1(n895), .B2(\unit_decode/n1504 ), 
        .ZN(\unit_decode/RegisterFile/n1832 ) );
  OAI22_X1 U1616 ( .A1(n898), .A2(n748), .B1(n895), .B2(\unit_decode/n1505 ), 
        .ZN(\unit_decode/RegisterFile/n1833 ) );
  OAI22_X1 U1617 ( .A1(n897), .A2(n745), .B1(n895), .B2(\unit_decode/n1506 ), 
        .ZN(\unit_decode/RegisterFile/n1834 ) );
  OAI22_X1 U1618 ( .A1(n897), .A2(n742), .B1(n895), .B2(\unit_decode/n1507 ), 
        .ZN(\unit_decode/RegisterFile/n1835 ) );
  OAI22_X1 U1619 ( .A1(n875), .A2(n811), .B1(n868), .B2(\unit_decode/n1556 ), 
        .ZN(\unit_decode/RegisterFile/n1908 ) );
  OAI22_X1 U1620 ( .A1(n875), .A2(n808), .B1(n868), .B2(\unit_decode/n1557 ), 
        .ZN(\unit_decode/RegisterFile/n1909 ) );
  OAI22_X1 U1621 ( .A1(n874), .A2(n805), .B1(n868), .B2(\unit_decode/n1558 ), 
        .ZN(\unit_decode/RegisterFile/n1910 ) );
  OAI22_X1 U1622 ( .A1(n874), .A2(n802), .B1(n868), .B2(\unit_decode/n1559 ), 
        .ZN(\unit_decode/RegisterFile/n1911 ) );
  OAI22_X1 U1623 ( .A1(n874), .A2(n799), .B1(n868), .B2(\unit_decode/n1560 ), 
        .ZN(\unit_decode/RegisterFile/n1912 ) );
  OAI22_X1 U1624 ( .A1(n874), .A2(n796), .B1(n868), .B2(\unit_decode/n1561 ), 
        .ZN(\unit_decode/RegisterFile/n1913 ) );
  OAI22_X1 U1625 ( .A1(n874), .A2(n793), .B1(n868), .B2(\unit_decode/n1562 ), 
        .ZN(\unit_decode/RegisterFile/n1914 ) );
  OAI22_X1 U1626 ( .A1(n873), .A2(n790), .B1(n868), .B2(\unit_decode/n1563 ), 
        .ZN(\unit_decode/RegisterFile/n1915 ) );
  OAI22_X1 U1627 ( .A1(n873), .A2(n787), .B1(n868), .B2(\unit_decode/n1564 ), 
        .ZN(\unit_decode/RegisterFile/n1916 ) );
  OAI22_X1 U1628 ( .A1(n873), .A2(n784), .B1(n868), .B2(\unit_decode/n1565 ), 
        .ZN(\unit_decode/RegisterFile/n1917 ) );
  OAI22_X1 U1629 ( .A1(n873), .A2(n781), .B1(n868), .B2(\unit_decode/n1566 ), 
        .ZN(\unit_decode/RegisterFile/n1918 ) );
  OAI22_X1 U1630 ( .A1(n873), .A2(n778), .B1(n868), .B2(\unit_decode/n1567 ), 
        .ZN(\unit_decode/RegisterFile/n1919 ) );
  OAI22_X1 U1631 ( .A1(n872), .A2(n775), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1568 ), .ZN(\unit_decode/RegisterFile/n1920 ) );
  OAI22_X1 U1632 ( .A1(n872), .A2(n772), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1569 ), .ZN(\unit_decode/RegisterFile/n1921 ) );
  OAI22_X1 U1633 ( .A1(n872), .A2(n769), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1570 ), .ZN(\unit_decode/RegisterFile/n1922 ) );
  OAI22_X1 U1634 ( .A1(n872), .A2(n766), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1571 ), .ZN(\unit_decode/RegisterFile/n1923 ) );
  OAI22_X1 U1635 ( .A1(n872), .A2(n763), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1572 ), .ZN(\unit_decode/RegisterFile/n1924 ) );
  OAI22_X1 U1636 ( .A1(n871), .A2(n760), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1573 ), .ZN(\unit_decode/RegisterFile/n1925 ) );
  OAI22_X1 U1637 ( .A1(n871), .A2(n757), .B1(\unit_decode/n2242 ), .B2(
        \unit_decode/n1574 ), .ZN(\unit_decode/RegisterFile/n1926 ) );
  OAI22_X1 U1638 ( .A1(n871), .A2(n754), .B1(n868), .B2(\unit_decode/n1575 ), 
        .ZN(\unit_decode/RegisterFile/n1927 ) );
  OAI22_X1 U1639 ( .A1(n871), .A2(n751), .B1(n868), .B2(\unit_decode/n1576 ), 
        .ZN(\unit_decode/RegisterFile/n1928 ) );
  OAI22_X1 U1640 ( .A1(n871), .A2(n748), .B1(n868), .B2(\unit_decode/n1577 ), 
        .ZN(\unit_decode/RegisterFile/n1929 ) );
  OAI22_X1 U1641 ( .A1(n870), .A2(n745), .B1(n868), .B2(\unit_decode/n1578 ), 
        .ZN(\unit_decode/RegisterFile/n1930 ) );
  OAI22_X1 U1642 ( .A1(n870), .A2(n742), .B1(n868), .B2(\unit_decode/n1579 ), 
        .ZN(\unit_decode/RegisterFile/n1931 ) );
  OAI22_X1 U1643 ( .A1(n866), .A2(n811), .B1(n859), .B2(\unit_decode/n1580 ), 
        .ZN(\unit_decode/RegisterFile/n1940 ) );
  OAI22_X1 U1644 ( .A1(n866), .A2(n808), .B1(n859), .B2(\unit_decode/n1581 ), 
        .ZN(\unit_decode/RegisterFile/n1941 ) );
  OAI22_X1 U1645 ( .A1(n865), .A2(n805), .B1(n859), .B2(\unit_decode/n1582 ), 
        .ZN(\unit_decode/RegisterFile/n1942 ) );
  OAI22_X1 U1646 ( .A1(n865), .A2(n802), .B1(n859), .B2(\unit_decode/n1583 ), 
        .ZN(\unit_decode/RegisterFile/n1943 ) );
  OAI22_X1 U1647 ( .A1(n865), .A2(n799), .B1(n859), .B2(\unit_decode/n1584 ), 
        .ZN(\unit_decode/RegisterFile/n1944 ) );
  OAI22_X1 U1648 ( .A1(n865), .A2(n796), .B1(n859), .B2(\unit_decode/n1585 ), 
        .ZN(\unit_decode/RegisterFile/n1945 ) );
  OAI22_X1 U1649 ( .A1(n865), .A2(n793), .B1(n859), .B2(\unit_decode/n1586 ), 
        .ZN(\unit_decode/RegisterFile/n1946 ) );
  OAI22_X1 U1650 ( .A1(n864), .A2(n790), .B1(n859), .B2(\unit_decode/n1587 ), 
        .ZN(\unit_decode/RegisterFile/n1947 ) );
  OAI22_X1 U1651 ( .A1(n864), .A2(n787), .B1(n859), .B2(\unit_decode/n1588 ), 
        .ZN(\unit_decode/RegisterFile/n1948 ) );
  OAI22_X1 U1652 ( .A1(n864), .A2(n784), .B1(n859), .B2(\unit_decode/n1589 ), 
        .ZN(\unit_decode/RegisterFile/n1949 ) );
  OAI22_X1 U1653 ( .A1(n864), .A2(n781), .B1(n859), .B2(\unit_decode/n1590 ), 
        .ZN(\unit_decode/RegisterFile/n1950 ) );
  OAI22_X1 U1654 ( .A1(n864), .A2(n778), .B1(n859), .B2(\unit_decode/n1591 ), 
        .ZN(\unit_decode/RegisterFile/n1951 ) );
  OAI22_X1 U1655 ( .A1(n863), .A2(n775), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1592 ), .ZN(\unit_decode/RegisterFile/n1952 ) );
  OAI22_X1 U1656 ( .A1(n863), .A2(n772), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1593 ), .ZN(\unit_decode/RegisterFile/n1953 ) );
  OAI22_X1 U1657 ( .A1(n863), .A2(n769), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1594 ), .ZN(\unit_decode/RegisterFile/n1954 ) );
  OAI22_X1 U1658 ( .A1(n863), .A2(n766), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1595 ), .ZN(\unit_decode/RegisterFile/n1955 ) );
  OAI22_X1 U1659 ( .A1(n863), .A2(n763), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1596 ), .ZN(\unit_decode/RegisterFile/n1956 ) );
  OAI22_X1 U1660 ( .A1(n862), .A2(n760), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1597 ), .ZN(\unit_decode/RegisterFile/n1957 ) );
  OAI22_X1 U1661 ( .A1(n862), .A2(n757), .B1(\unit_decode/n2240 ), .B2(
        \unit_decode/n1598 ), .ZN(\unit_decode/RegisterFile/n1958 ) );
  OAI22_X1 U1662 ( .A1(n862), .A2(n754), .B1(n859), .B2(\unit_decode/n1599 ), 
        .ZN(\unit_decode/RegisterFile/n1959 ) );
  OAI22_X1 U1663 ( .A1(n862), .A2(n751), .B1(n859), .B2(\unit_decode/n1600 ), 
        .ZN(\unit_decode/RegisterFile/n1960 ) );
  OAI22_X1 U1664 ( .A1(n862), .A2(n748), .B1(n859), .B2(\unit_decode/n1601 ), 
        .ZN(\unit_decode/RegisterFile/n1961 ) );
  OAI22_X1 U1665 ( .A1(n861), .A2(n745), .B1(n859), .B2(\unit_decode/n1602 ), 
        .ZN(\unit_decode/RegisterFile/n1962 ) );
  OAI22_X1 U1666 ( .A1(n861), .A2(n742), .B1(n859), .B2(\unit_decode/n1603 ), 
        .ZN(\unit_decode/RegisterFile/n1963 ) );
  OAI22_X1 U1667 ( .A1(n839), .A2(n811), .B1(n832), .B2(\unit_decode/n1652 ), 
        .ZN(\unit_decode/RegisterFile/n2036 ) );
  OAI22_X1 U1668 ( .A1(n839), .A2(n808), .B1(n832), .B2(\unit_decode/n1653 ), 
        .ZN(\unit_decode/RegisterFile/n2037 ) );
  OAI22_X1 U1669 ( .A1(n838), .A2(n805), .B1(n832), .B2(\unit_decode/n1654 ), 
        .ZN(\unit_decode/RegisterFile/n2038 ) );
  OAI22_X1 U1670 ( .A1(n838), .A2(n802), .B1(n832), .B2(\unit_decode/n1655 ), 
        .ZN(\unit_decode/RegisterFile/n2039 ) );
  OAI22_X1 U1671 ( .A1(n838), .A2(n799), .B1(n832), .B2(\unit_decode/n1656 ), 
        .ZN(\unit_decode/RegisterFile/n2040 ) );
  OAI22_X1 U1672 ( .A1(n838), .A2(n796), .B1(n832), .B2(\unit_decode/n1657 ), 
        .ZN(\unit_decode/RegisterFile/n2041 ) );
  OAI22_X1 U1673 ( .A1(n838), .A2(n793), .B1(n832), .B2(\unit_decode/n1658 ), 
        .ZN(\unit_decode/RegisterFile/n2042 ) );
  OAI22_X1 U1674 ( .A1(n837), .A2(n790), .B1(n832), .B2(\unit_decode/n1659 ), 
        .ZN(\unit_decode/RegisterFile/n2043 ) );
  OAI22_X1 U1675 ( .A1(n837), .A2(n787), .B1(n832), .B2(\unit_decode/n1660 ), 
        .ZN(\unit_decode/RegisterFile/n2044 ) );
  OAI22_X1 U1676 ( .A1(n837), .A2(n784), .B1(n832), .B2(\unit_decode/n1661 ), 
        .ZN(\unit_decode/RegisterFile/n2045 ) );
  OAI22_X1 U1677 ( .A1(n837), .A2(n781), .B1(n832), .B2(\unit_decode/n1662 ), 
        .ZN(\unit_decode/RegisterFile/n2046 ) );
  OAI22_X1 U1678 ( .A1(n837), .A2(n778), .B1(n832), .B2(\unit_decode/n1663 ), 
        .ZN(\unit_decode/RegisterFile/n2047 ) );
  OAI22_X1 U1679 ( .A1(n836), .A2(n775), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1664 ), .ZN(\unit_decode/RegisterFile/n2048 ) );
  OAI22_X1 U1680 ( .A1(n836), .A2(n772), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1665 ), .ZN(\unit_decode/RegisterFile/n2049 ) );
  OAI22_X1 U1681 ( .A1(n836), .A2(n769), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1666 ), .ZN(\unit_decode/RegisterFile/n2050 ) );
  OAI22_X1 U1682 ( .A1(n836), .A2(n766), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1667 ), .ZN(\unit_decode/RegisterFile/n2051 ) );
  OAI22_X1 U1683 ( .A1(n836), .A2(n763), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1668 ), .ZN(\unit_decode/RegisterFile/n2052 ) );
  OAI22_X1 U1684 ( .A1(n835), .A2(n760), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1669 ), .ZN(\unit_decode/RegisterFile/n2053 ) );
  OAI22_X1 U1685 ( .A1(n835), .A2(n757), .B1(\unit_decode/n2234 ), .B2(
        \unit_decode/n1670 ), .ZN(\unit_decode/RegisterFile/n2054 ) );
  OAI22_X1 U1686 ( .A1(n835), .A2(n754), .B1(n832), .B2(\unit_decode/n1671 ), 
        .ZN(\unit_decode/RegisterFile/n2055 ) );
  OAI22_X1 U1687 ( .A1(n835), .A2(n751), .B1(n832), .B2(\unit_decode/n1672 ), 
        .ZN(\unit_decode/RegisterFile/n2056 ) );
  OAI22_X1 U1688 ( .A1(n835), .A2(n748), .B1(n832), .B2(\unit_decode/n1673 ), 
        .ZN(\unit_decode/RegisterFile/n2057 ) );
  OAI22_X1 U1689 ( .A1(n834), .A2(n745), .B1(n832), .B2(\unit_decode/n1674 ), 
        .ZN(\unit_decode/RegisterFile/n2058 ) );
  OAI22_X1 U1690 ( .A1(n834), .A2(n742), .B1(n832), .B2(\unit_decode/n1675 ), 
        .ZN(\unit_decode/RegisterFile/n2059 ) );
  OAI22_X1 U1691 ( .A1(n830), .A2(n811), .B1(n823), .B2(\unit_decode/n1676 ), 
        .ZN(\unit_decode/RegisterFile/n2068 ) );
  OAI22_X1 U1692 ( .A1(n830), .A2(n808), .B1(n823), .B2(\unit_decode/n1677 ), 
        .ZN(\unit_decode/RegisterFile/n2069 ) );
  OAI22_X1 U1693 ( .A1(n829), .A2(n805), .B1(n823), .B2(\unit_decode/n1678 ), 
        .ZN(\unit_decode/RegisterFile/n2070 ) );
  OAI22_X1 U1694 ( .A1(n829), .A2(n802), .B1(n823), .B2(\unit_decode/n1679 ), 
        .ZN(\unit_decode/RegisterFile/n2071 ) );
  OAI22_X1 U1695 ( .A1(n829), .A2(n799), .B1(n823), .B2(\unit_decode/n1680 ), 
        .ZN(\unit_decode/RegisterFile/n2072 ) );
  OAI22_X1 U1696 ( .A1(n829), .A2(n796), .B1(n823), .B2(\unit_decode/n1681 ), 
        .ZN(\unit_decode/RegisterFile/n2073 ) );
  OAI22_X1 U1697 ( .A1(n829), .A2(n793), .B1(n823), .B2(\unit_decode/n1682 ), 
        .ZN(\unit_decode/RegisterFile/n2074 ) );
  OAI22_X1 U1698 ( .A1(n828), .A2(n790), .B1(n823), .B2(\unit_decode/n1683 ), 
        .ZN(\unit_decode/RegisterFile/n2075 ) );
  OAI22_X1 U1699 ( .A1(n828), .A2(n787), .B1(n823), .B2(\unit_decode/n1684 ), 
        .ZN(\unit_decode/RegisterFile/n2076 ) );
  OAI22_X1 U1700 ( .A1(n828), .A2(n784), .B1(n823), .B2(\unit_decode/n1685 ), 
        .ZN(\unit_decode/RegisterFile/n2077 ) );
  OAI22_X1 U1701 ( .A1(n828), .A2(n781), .B1(n823), .B2(\unit_decode/n1686 ), 
        .ZN(\unit_decode/RegisterFile/n2078 ) );
  OAI22_X1 U1702 ( .A1(n828), .A2(n778), .B1(n823), .B2(\unit_decode/n1687 ), 
        .ZN(\unit_decode/RegisterFile/n2079 ) );
  OAI22_X1 U1703 ( .A1(n827), .A2(n775), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1688 ), .ZN(\unit_decode/RegisterFile/n2080 ) );
  OAI22_X1 U1704 ( .A1(n827), .A2(n772), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1689 ), .ZN(\unit_decode/RegisterFile/n2081 ) );
  OAI22_X1 U1705 ( .A1(n827), .A2(n769), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1690 ), .ZN(\unit_decode/RegisterFile/n2082 ) );
  OAI22_X1 U1706 ( .A1(n827), .A2(n766), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1691 ), .ZN(\unit_decode/RegisterFile/n2083 ) );
  OAI22_X1 U1707 ( .A1(n827), .A2(n763), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1692 ), .ZN(\unit_decode/RegisterFile/n2084 ) );
  OAI22_X1 U1708 ( .A1(n826), .A2(n760), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1693 ), .ZN(\unit_decode/RegisterFile/n2085 ) );
  OAI22_X1 U1709 ( .A1(n826), .A2(n757), .B1(\unit_decode/n2232 ), .B2(
        \unit_decode/n1694 ), .ZN(\unit_decode/RegisterFile/n2086 ) );
  OAI22_X1 U1710 ( .A1(n826), .A2(n754), .B1(n823), .B2(\unit_decode/n1695 ), 
        .ZN(\unit_decode/RegisterFile/n2087 ) );
  OAI22_X1 U1711 ( .A1(n826), .A2(n751), .B1(n823), .B2(\unit_decode/n1696 ), 
        .ZN(\unit_decode/RegisterFile/n2088 ) );
  OAI22_X1 U1712 ( .A1(n826), .A2(n748), .B1(n823), .B2(\unit_decode/n1697 ), 
        .ZN(\unit_decode/RegisterFile/n2089 ) );
  OAI22_X1 U1713 ( .A1(n825), .A2(n745), .B1(n823), .B2(\unit_decode/n1698 ), 
        .ZN(\unit_decode/RegisterFile/n2090 ) );
  OAI22_X1 U1714 ( .A1(n825), .A2(n742), .B1(n823), .B2(\unit_decode/n1699 ), 
        .ZN(\unit_decode/RegisterFile/n2091 ) );
  OAI22_X1 U1715 ( .A1(n969), .A2(n743), .B1(n967), .B2(\unit_decode/n2012 ), 
        .ZN(\unit_decode/RegisterFile/n1579 ) );
  OAI22_X1 U1716 ( .A1(n969), .A2(n746), .B1(n967), .B2(\unit_decode/n2013 ), 
        .ZN(\unit_decode/RegisterFile/n1578 ) );
  OAI22_X1 U1717 ( .A1(n970), .A2(n749), .B1(n967), .B2(\unit_decode/n2014 ), 
        .ZN(\unit_decode/RegisterFile/n1577 ) );
  OAI22_X1 U1718 ( .A1(n970), .A2(n752), .B1(n967), .B2(\unit_decode/n2015 ), 
        .ZN(\unit_decode/RegisterFile/n1576 ) );
  OAI22_X1 U1719 ( .A1(n970), .A2(n755), .B1(n967), .B2(\unit_decode/n2016 ), 
        .ZN(\unit_decode/RegisterFile/n1575 ) );
  OAI22_X1 U1720 ( .A1(n970), .A2(n758), .B1(n967), .B2(\unit_decode/n2017 ), 
        .ZN(\unit_decode/RegisterFile/n1574 ) );
  OAI22_X1 U1721 ( .A1(n970), .A2(n761), .B1(n967), .B2(\unit_decode/n2018 ), 
        .ZN(\unit_decode/RegisterFile/n1573 ) );
  OAI22_X1 U1722 ( .A1(n971), .A2(n764), .B1(n967), .B2(\unit_decode/n2019 ), 
        .ZN(\unit_decode/RegisterFile/n1572 ) );
  OAI22_X1 U1723 ( .A1(n971), .A2(n767), .B1(n967), .B2(\unit_decode/n2020 ), 
        .ZN(\unit_decode/RegisterFile/n1571 ) );
  OAI22_X1 U1724 ( .A1(n971), .A2(n770), .B1(n967), .B2(\unit_decode/n2021 ), 
        .ZN(\unit_decode/RegisterFile/n1570 ) );
  OAI22_X1 U1725 ( .A1(n971), .A2(n773), .B1(n967), .B2(\unit_decode/n2022 ), 
        .ZN(\unit_decode/RegisterFile/n1569 ) );
  OAI22_X1 U1726 ( .A1(n971), .A2(n776), .B1(n967), .B2(\unit_decode/n2023 ), 
        .ZN(\unit_decode/RegisterFile/n1568 ) );
  OAI22_X1 U1727 ( .A1(n972), .A2(n779), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2024 ), .ZN(\unit_decode/RegisterFile/n1567 ) );
  OAI22_X1 U1728 ( .A1(n972), .A2(n782), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2025 ), .ZN(\unit_decode/RegisterFile/n1566 ) );
  OAI22_X1 U1729 ( .A1(n972), .A2(n785), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2026 ), .ZN(\unit_decode/RegisterFile/n1565 ) );
  OAI22_X1 U1730 ( .A1(n972), .A2(n788), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2027 ), .ZN(\unit_decode/RegisterFile/n1564 ) );
  OAI22_X1 U1731 ( .A1(n972), .A2(n791), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2028 ), .ZN(\unit_decode/RegisterFile/n1563 ) );
  OAI22_X1 U1732 ( .A1(n973), .A2(n794), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2029 ), .ZN(\unit_decode/RegisterFile/n1562 ) );
  OAI22_X1 U1733 ( .A1(n973), .A2(n797), .B1(\unit_decode/n2257 ), .B2(
        \unit_decode/n2030 ), .ZN(\unit_decode/RegisterFile/n1561 ) );
  OAI22_X1 U1734 ( .A1(n973), .A2(n800), .B1(n967), .B2(\unit_decode/n2031 ), 
        .ZN(\unit_decode/RegisterFile/n1560 ) );
  OAI22_X1 U1735 ( .A1(n973), .A2(n803), .B1(n967), .B2(\unit_decode/n2032 ), 
        .ZN(\unit_decode/RegisterFile/n1559 ) );
  OAI22_X1 U1736 ( .A1(n973), .A2(n806), .B1(n967), .B2(\unit_decode/n2033 ), 
        .ZN(\unit_decode/RegisterFile/n1558 ) );
  OAI22_X1 U1737 ( .A1(n974), .A2(n809), .B1(n967), .B2(\unit_decode/n2034 ), 
        .ZN(\unit_decode/RegisterFile/n1557 ) );
  OAI22_X1 U1738 ( .A1(n974), .A2(n812), .B1(n967), .B2(\unit_decode/n2035 ), 
        .ZN(\unit_decode/RegisterFile/n1556 ) );
  OAI22_X1 U1739 ( .A1(n942), .A2(n743), .B1(n940), .B2(\unit_decode/n2084 ), 
        .ZN(\unit_decode/RegisterFile/n1675 ) );
  BUF_X1 U1740 ( .A(\unit_memory/DRAM/n722 ), .Z(n251) );
  AND2_X2 U1741 ( .A1(n1353), .A2(n1697), .ZN(n104) );
  AND3_X1 U1742 ( .A1(n1697), .A2(n1655), .A3(n1539), .ZN(n105) );
  BUF_X1 U1743 ( .A(\unit_memory/DRAM/n724 ), .Z(n268) );
  BUF_X1 U1744 ( .A(\unit_memory/DRAM/n725 ), .Z(n271) );
  BUF_X1 U1745 ( .A(\unit_memory/DRAM/n726 ), .Z(n274) );
  BUF_X1 U1746 ( .A(\unit_memory/DRAM/n727 ), .Z(n277) );
  BUF_X1 U1747 ( .A(\unit_memory/DRAM/n728 ), .Z(n280) );
  BUF_X1 U1748 ( .A(\unit_memory/DRAM/n729 ), .Z(n283) );
  BUF_X1 U1749 ( .A(\unit_memory/DRAM/n730 ), .Z(n286) );
  BUF_X1 U1750 ( .A(\unit_memory/DRAM/n731 ), .Z(n289) );
  BUF_X1 U1751 ( .A(\unit_memory/DRAM/n732 ), .Z(n292) );
  BUF_X1 U1752 ( .A(\unit_memory/DRAM/n733 ), .Z(n295) );
  BUF_X1 U1753 ( .A(\unit_memory/DRAM/n734 ), .Z(n298) );
  BUF_X1 U1754 ( .A(\unit_memory/DRAM/n735 ), .Z(n301) );
  BUF_X1 U1755 ( .A(\unit_memory/DRAM/n736 ), .Z(n304) );
  BUF_X1 U1756 ( .A(\unit_memory/DRAM/n737 ), .Z(n307) );
  BUF_X1 U1757 ( .A(\unit_memory/DRAM/n738 ), .Z(n310) );
  BUF_X1 U1758 ( .A(\unit_memory/DRAM/n739 ), .Z(n313) );
  BUF_X1 U1759 ( .A(\unit_memory/DRAM/n740 ), .Z(n316) );
  BUF_X1 U1760 ( .A(\unit_memory/DRAM/n741 ), .Z(n319) );
  BUF_X1 U1761 ( .A(\unit_memory/DRAM/n742 ), .Z(n322) );
  BUF_X1 U1762 ( .A(\unit_memory/DRAM/n743 ), .Z(n325) );
  BUF_X1 U1763 ( .A(\unit_memory/DRAM/n744 ), .Z(n328) );
  BUF_X1 U1764 ( .A(\unit_memory/DRAM/n745 ), .Z(n331) );
  BUF_X1 U1765 ( .A(\unit_memory/DRAM/n746 ), .Z(n334) );
  BUF_X1 U1766 ( .A(\unit_memory/DRAM/n747 ), .Z(n337) );
  BUF_X1 U1767 ( .A(\unit_memory/DRAM/n748 ), .Z(n340) );
  BUF_X1 U1768 ( .A(\unit_memory/DRAM/n749 ), .Z(n343) );
  BUF_X1 U1769 ( .A(\unit_memory/DRAM/n750 ), .Z(n346) );
  BUF_X1 U1770 ( .A(\unit_memory/DRAM/n751 ), .Z(n349) );
  BUF_X1 U1771 ( .A(\unit_memory/DRAM/n752 ), .Z(n352) );
  BUF_X1 U1772 ( .A(\unit_memory/DRAM/n753 ), .Z(n355) );
  BUF_X1 U1773 ( .A(\unit_memory/DRAM/n754 ), .Z(n358) );
  NAND2_X1 U1774 ( .A1(\unit_memory/DRAM/n755 ), .A2(\unit_memory/DRAM/n756 ), 
        .ZN(\unit_memory/DRAM/n723 ) );
  NAND2_X1 U1775 ( .A1(\unit_decode/n2186 ), .A2(n1345), .ZN(
        \unit_decode/n3513 ) );
  AND2_X1 U1776 ( .A1(net130925), .A2(n114), .ZN(n106) );
  AND2_X1 U1777 ( .A1(net130925), .A2(n36), .ZN(n107) );
  INV_X1 U1778 ( .A(\unit_decode/n2270 ), .ZN(n1083) );
  OAI21_X1 U1779 ( .B1(\unit_decode/n2241 ), .B2(\unit_decode/n2264 ), .A(
        n1350), .ZN(\unit_decode/n2270 ) );
  INV_X1 U1780 ( .A(\unit_decode/n2269 ), .ZN(n1074) );
  OAI21_X1 U1781 ( .B1(\unit_decode/n2239 ), .B2(\unit_decode/n2264 ), .A(
        n1350), .ZN(\unit_decode/n2269 ) );
  INV_X1 U1782 ( .A(\unit_decode/n2268 ), .ZN(n1065) );
  OAI21_X1 U1783 ( .B1(\unit_decode/n2237 ), .B2(\unit_decode/n2264 ), .A(
        n1350), .ZN(\unit_decode/n2268 ) );
  INV_X1 U1784 ( .A(\unit_decode/n2267 ), .ZN(n1056) );
  OAI21_X1 U1785 ( .B1(\unit_decode/n2235 ), .B2(\unit_decode/n2264 ), .A(
        n1349), .ZN(\unit_decode/n2267 ) );
  INV_X1 U1786 ( .A(\unit_decode/n2266 ), .ZN(n1047) );
  OAI21_X1 U1787 ( .B1(\unit_decode/n2233 ), .B2(\unit_decode/n2264 ), .A(
        n1349), .ZN(\unit_decode/n2266 ) );
  INV_X1 U1788 ( .A(\unit_decode/n2265 ), .ZN(n1038) );
  OAI21_X1 U1789 ( .B1(\unit_decode/n2231 ), .B2(\unit_decode/n2264 ), .A(
        n1349), .ZN(\unit_decode/n2265 ) );
  INV_X1 U1790 ( .A(\unit_decode/n2263 ), .ZN(n1029) );
  OAI21_X1 U1791 ( .B1(\unit_decode/n2229 ), .B2(\unit_decode/n2264 ), .A(
        n1349), .ZN(\unit_decode/n2263 ) );
  INV_X1 U1792 ( .A(\unit_decode/n2242 ), .ZN(n876) );
  OAI21_X1 U1793 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2243 ), .A(
        n1348), .ZN(\unit_decode/n2242 ) );
  INV_X1 U1794 ( .A(\unit_decode/n2240 ), .ZN(n867) );
  OAI21_X1 U1795 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2241 ), .A(
        n1348), .ZN(\unit_decode/n2240 ) );
  INV_X1 U1796 ( .A(\unit_decode/n2238 ), .ZN(n858) );
  OAI21_X1 U1797 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2239 ), .A(
        n1348), .ZN(\unit_decode/n2238 ) );
  INV_X1 U1798 ( .A(\unit_decode/n2236 ), .ZN(n849) );
  OAI21_X1 U1799 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2237 ), .A(
        n1348), .ZN(\unit_decode/n2236 ) );
  INV_X1 U1800 ( .A(\unit_decode/n2234 ), .ZN(n840) );
  OAI21_X1 U1801 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2235 ), .A(
        n1347), .ZN(\unit_decode/n2234 ) );
  INV_X1 U1802 ( .A(\unit_decode/n2232 ), .ZN(n831) );
  OAI21_X1 U1803 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2233 ), .A(
        n1348), .ZN(\unit_decode/n2232 ) );
  INV_X1 U1804 ( .A(\unit_decode/n2230 ), .ZN(n822) );
  OAI21_X1 U1805 ( .B1(\unit_decode/n2228 ), .B2(\unit_decode/n2231 ), .A(
        n1347), .ZN(\unit_decode/n2230 ) );
  NAND2_X1 U1806 ( .A1(n137), .A2(n1345), .ZN(\unit_decode/n3512 ) );
  NOR2_X1 U1807 ( .A1(\unit_decode/n2094 ), .A2(\unit_decode/n2095 ), .ZN(
        \unit_decode/n3492 ) );
  NOR2_X1 U1808 ( .A1(\unit_decode/n2099 ), .A2(\unit_decode/n2100 ), .ZN(
        \unit_decode/n2872 ) );
  NOR3_X1 U1809 ( .A1(\unit_decode/n2097 ), .A2(\unit_decode/n2098 ), .A3(
        \unit_decode/n2096 ), .ZN(\unit_decode/n2879 ) );
  NOR3_X1 U1810 ( .A1(\unit_decode/n2092 ), .A2(\unit_decode/n2093 ), .A3(
        \unit_decode/n2091 ), .ZN(\unit_decode/n3499 ) );
  NOR2_X1 U1811 ( .A1(\unit_decode/n2095 ), .A2(IR_OUT[22]), .ZN(
        \unit_decode/n3490 ) );
  OAI221_X1 U1812 ( .B1(\unit_decode/n1769 ), .B2(n1167), .C1(
        \unit_decode/n1766 ), .C2(n1170), .A(\unit_decode/n2356 ), .ZN(
        \unit_decode/n2351 ) );
  AOI22_X1 U1813 ( .A1(n1173), .A2(\unit_decode/n1785 ), .B1(n1174), .B2(
        \unit_decode/n1777 ), .ZN(\unit_decode/n2356 ) );
  OAI221_X1 U1814 ( .B1(\unit_decode/n1768 ), .B2(n1167), .C1(
        \unit_decode/n1765 ), .C2(n1170), .A(\unit_decode/n2338 ), .ZN(
        \unit_decode/n2333 ) );
  AOI22_X1 U1815 ( .A1(n1173), .A2(\unit_decode/n1784 ), .B1(n1174), .B2(
        \unit_decode/n1776 ), .ZN(\unit_decode/n2338 ) );
  OAI221_X1 U1816 ( .B1(\unit_decode/n1767 ), .B2(n1167), .C1(
        \unit_decode/n1764 ), .C2(n1170), .A(\unit_decode/n2314 ), .ZN(
        \unit_decode/n2299 ) );
  AOI22_X1 U1817 ( .A1(n1173), .A2(\unit_decode/n1783 ), .B1(n1174), .B2(
        \unit_decode/n1775 ), .ZN(\unit_decode/n2314 ) );
  OAI221_X1 U1818 ( .B1(\unit_decode/n1769 ), .B2(n1263), .C1(
        \unit_decode/n1766 ), .C2(n1266), .A(\unit_decode/n2976 ), .ZN(
        \unit_decode/n2971 ) );
  AOI22_X1 U1819 ( .A1(n1269), .A2(\unit_decode/n1785 ), .B1(n1270), .B2(
        \unit_decode/n1777 ), .ZN(\unit_decode/n2976 ) );
  OAI221_X1 U1820 ( .B1(\unit_decode/n1768 ), .B2(n1263), .C1(
        \unit_decode/n1765 ), .C2(n1266), .A(\unit_decode/n2958 ), .ZN(
        \unit_decode/n2953 ) );
  AOI22_X1 U1821 ( .A1(n1269), .A2(\unit_decode/n1784 ), .B1(n1270), .B2(
        \unit_decode/n1776 ), .ZN(\unit_decode/n2958 ) );
  OAI221_X1 U1822 ( .B1(\unit_decode/n1767 ), .B2(n1263), .C1(
        \unit_decode/n1764 ), .C2(n1266), .A(\unit_decode/n2934 ), .ZN(
        \unit_decode/n2919 ) );
  AOI22_X1 U1823 ( .A1(n1269), .A2(\unit_decode/n1783 ), .B1(n1270), .B2(
        \unit_decode/n1775 ), .ZN(\unit_decode/n2934 ) );
  AOI22_X1 U1824 ( .A1(n1185), .A2(\unit_decode/n1891 ), .B1(n1186), .B2(
        \unit_decode/n1883 ), .ZN(\unit_decode/n2447 ) );
  AOI22_X1 U1825 ( .A1(n1185), .A2(\unit_decode/n1890 ), .B1(n1186), .B2(
        \unit_decode/n1882 ), .ZN(\unit_decode/n2429 ) );
  AOI22_X1 U1826 ( .A1(n1185), .A2(\unit_decode/n1889 ), .B1(n1186), .B2(
        \unit_decode/n1881 ), .ZN(\unit_decode/n2411 ) );
  AOI22_X1 U1827 ( .A1(n1185), .A2(\unit_decode/n1888 ), .B1(n1186), .B2(
        \unit_decode/n1880 ), .ZN(\unit_decode/n2393 ) );
  AOI22_X1 U1828 ( .A1(n1185), .A2(\unit_decode/n1887 ), .B1(n1186), .B2(
        \unit_decode/n1879 ), .ZN(\unit_decode/n2375 ) );
  AOI22_X1 U1829 ( .A1(n1185), .A2(\unit_decode/n1886 ), .B1(n1186), .B2(
        \unit_decode/n1878 ), .ZN(\unit_decode/n2357 ) );
  AOI22_X1 U1830 ( .A1(n1185), .A2(\unit_decode/n1885 ), .B1(n1186), .B2(
        \unit_decode/n1877 ), .ZN(\unit_decode/n2339 ) );
  AOI22_X1 U1831 ( .A1(n1185), .A2(\unit_decode/n1884 ), .B1(n1186), .B2(
        \unit_decode/n1876 ), .ZN(\unit_decode/n2319 ) );
  AOI22_X1 U1832 ( .A1(n1281), .A2(\unit_decode/n1891 ), .B1(n1282), .B2(
        \unit_decode/n1883 ), .ZN(\unit_decode/n3067 ) );
  AOI22_X1 U1833 ( .A1(n1281), .A2(\unit_decode/n1890 ), .B1(n1282), .B2(
        \unit_decode/n1882 ), .ZN(\unit_decode/n3049 ) );
  AOI22_X1 U1834 ( .A1(n1281), .A2(\unit_decode/n1889 ), .B1(n1282), .B2(
        \unit_decode/n1881 ), .ZN(\unit_decode/n3031 ) );
  AOI22_X1 U1835 ( .A1(n1281), .A2(\unit_decode/n1888 ), .B1(n1282), .B2(
        \unit_decode/n1880 ), .ZN(\unit_decode/n3013 ) );
  AOI22_X1 U1836 ( .A1(n1281), .A2(\unit_decode/n1887 ), .B1(n1282), .B2(
        \unit_decode/n1879 ), .ZN(\unit_decode/n2995 ) );
  AOI22_X1 U1837 ( .A1(n1281), .A2(\unit_decode/n1886 ), .B1(n1282), .B2(
        \unit_decode/n1878 ), .ZN(\unit_decode/n2977 ) );
  AOI22_X1 U1838 ( .A1(n1281), .A2(\unit_decode/n1885 ), .B1(n1282), .B2(
        \unit_decode/n1877 ), .ZN(\unit_decode/n2959 ) );
  AOI22_X1 U1839 ( .A1(n1281), .A2(\unit_decode/n1884 ), .B1(n1282), .B2(
        \unit_decode/n1876 ), .ZN(\unit_decode/n2939 ) );
  NAND2_X1 U1840 ( .A1(\unit_decode/n2879 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2293 ) );
  NAND2_X1 U1841 ( .A1(\unit_decode/n3499 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2913 ) );
  BUF_X1 U1842 ( .A(\unit_memory/DRAM/n579 ), .Z(n223) );
  BUF_X1 U1843 ( .A(\unit_memory/DRAM/n580 ), .Z(n236) );
  BUF_X1 U1844 ( .A(\unit_memory/DRAM/n576 ), .Z(n197) );
  BUF_X1 U1845 ( .A(\unit_memory/DRAM/n577 ), .Z(n210) );
  NAND2_X1 U1846 ( .A1(\unit_decode/n3489 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2899 ) );
  NAND2_X1 U1847 ( .A1(\unit_decode/n3489 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2898 ) );
  NAND2_X1 U1848 ( .A1(\unit_decode/n3495 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2904 ) );
  NAND2_X1 U1849 ( .A1(\unit_decode/n3495 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2903 ) );
  NAND2_X1 U1850 ( .A1(\unit_decode/n3505 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2923 ) );
  NAND2_X1 U1851 ( .A1(\unit_decode/n3505 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2922 ) );
  NAND2_X1 U1852 ( .A1(\unit_decode/n3507 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2928 ) );
  NAND2_X1 U1853 ( .A1(\unit_decode/n3507 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2927 ) );
  NAND2_X1 U1854 ( .A1(\unit_decode/n2869 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2279 ) );
  NAND2_X1 U1855 ( .A1(\unit_decode/n2869 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2278 ) );
  NAND2_X1 U1856 ( .A1(\unit_decode/n2875 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2284 ) );
  NAND2_X1 U1857 ( .A1(\unit_decode/n2875 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2283 ) );
  NAND2_X1 U1858 ( .A1(\unit_decode/n2877 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2289 ) );
  NAND2_X1 U1859 ( .A1(\unit_decode/n2877 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2288 ) );
  NAND2_X1 U1860 ( .A1(\unit_decode/n2885 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2303 ) );
  NAND2_X1 U1861 ( .A1(\unit_decode/n2885 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2302 ) );
  NAND2_X1 U1862 ( .A1(\unit_decode/n2887 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2308 ) );
  NAND2_X1 U1863 ( .A1(\unit_decode/n2887 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2307 ) );
  NAND2_X1 U1864 ( .A1(\unit_decode/n2889 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2313 ) );
  NAND2_X1 U1865 ( .A1(\unit_decode/n2889 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2312 ) );
  NAND2_X1 U1866 ( .A1(\unit_decode/n2891 ), .A2(\unit_decode/n2872 ), .ZN(
        \unit_decode/n2318 ) );
  NAND2_X1 U1867 ( .A1(\unit_decode/n2891 ), .A2(\unit_decode/n2873 ), .ZN(
        \unit_decode/n2317 ) );
  NAND2_X1 U1868 ( .A1(\unit_decode/n3497 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2909 ) );
  NAND2_X1 U1869 ( .A1(\unit_decode/n3497 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2908 ) );
  NAND2_X1 U1870 ( .A1(\unit_decode/n3509 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2933 ) );
  NAND2_X1 U1871 ( .A1(\unit_decode/n3509 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2932 ) );
  NAND2_X1 U1872 ( .A1(\unit_decode/n3511 ), .A2(\unit_decode/n3492 ), .ZN(
        \unit_decode/n2938 ) );
  NAND2_X1 U1873 ( .A1(\unit_decode/n3511 ), .A2(\unit_decode/n3493 ), .ZN(
        \unit_decode/n2937 ) );
  NAND2_X1 U1874 ( .A1(\unit_decode/n2870 ), .A2(\unit_decode/n2879 ), .ZN(
        \unit_decode/n2294 ) );
  INV_X1 U1875 ( .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n548 ) );
  BUF_X1 U1876 ( .A(\unit_memory/DRAM/n580 ), .Z(n237) );
  BUF_X1 U1877 ( .A(\unit_memory/DRAM/n579 ), .Z(n224) );
  BUF_X1 U1878 ( .A(\unit_memory/DRAM/n576 ), .Z(n198) );
  BUF_X1 U1879 ( .A(\unit_memory/DRAM/n577 ), .Z(n211) );
  AND2_X1 U1880 ( .A1(\unit_decode/n2873 ), .A2(\unit_decode/n2879 ), .ZN(
        \unit_decode/n2296 ) );
  AND2_X1 U1881 ( .A1(\unit_decode/n3493 ), .A2(\unit_decode/n3499 ), .ZN(
        \unit_decode/n2916 ) );
  INV_X1 U1882 ( .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n549 ) );
  BUF_X1 U1883 ( .A(\unit_decode/RegisterFile/N445 ), .Z(n703) );
  BUF_X1 U1884 ( .A(\unit_decode/RegisterFile/N445 ), .Z(n704) );
  BUF_X1 U1885 ( .A(\unit_decode/RegisterFile/N444 ), .Z(n707) );
  BUF_X1 U1886 ( .A(\unit_decode/RegisterFile/N444 ), .Z(n706) );
  AND2_X1 U1887 ( .A1(\unit_decode/n2869 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2282 ) );
  AND2_X1 U1888 ( .A1(\unit_decode/n2869 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2281 ) );
  AND2_X1 U1889 ( .A1(\unit_decode/n2875 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2287 ) );
  AND2_X1 U1890 ( .A1(\unit_decode/n2875 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2286 ) );
  AND2_X1 U1891 ( .A1(\unit_decode/n2877 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2292 ) );
  AND2_X1 U1892 ( .A1(\unit_decode/n2877 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2291 ) );
  AND2_X1 U1893 ( .A1(\unit_decode/n2885 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2306 ) );
  AND2_X1 U1894 ( .A1(\unit_decode/n2885 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2305 ) );
  AND2_X1 U1895 ( .A1(\unit_decode/n2887 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2311 ) );
  AND2_X1 U1896 ( .A1(\unit_decode/n2887 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2310 ) );
  AND2_X1 U1897 ( .A1(\unit_decode/n2889 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2316 ) );
  AND2_X1 U1898 ( .A1(\unit_decode/n2889 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2315 ) );
  AND2_X1 U1899 ( .A1(\unit_decode/n2891 ), .A2(\unit_decode/n2870 ), .ZN(
        \unit_decode/n2321 ) );
  AND2_X1 U1900 ( .A1(\unit_decode/n2891 ), .A2(\unit_decode/n2871 ), .ZN(
        \unit_decode/n2320 ) );
  AND2_X1 U1901 ( .A1(\unit_decode/n3489 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2902 ) );
  AND2_X1 U1902 ( .A1(\unit_decode/n3489 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2901 ) );
  AND2_X1 U1903 ( .A1(\unit_decode/n3495 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2907 ) );
  AND2_X1 U1904 ( .A1(\unit_decode/n3495 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2906 ) );
  AND2_X1 U1905 ( .A1(\unit_decode/n3497 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2912 ) );
  AND2_X1 U1906 ( .A1(\unit_decode/n3497 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2911 ) );
  AND2_X1 U1907 ( .A1(\unit_decode/n3505 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2926 ) );
  AND2_X1 U1908 ( .A1(\unit_decode/n3505 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2925 ) );
  AND2_X1 U1909 ( .A1(\unit_decode/n3507 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2931 ) );
  AND2_X1 U1910 ( .A1(\unit_decode/n3507 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2930 ) );
  AND2_X1 U1911 ( .A1(\unit_decode/n3509 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2936 ) );
  AND2_X1 U1912 ( .A1(\unit_decode/n3509 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2935 ) );
  AND2_X1 U1913 ( .A1(\unit_decode/n3511 ), .A2(\unit_decode/n3490 ), .ZN(
        \unit_decode/n2941 ) );
  AND2_X1 U1914 ( .A1(\unit_decode/n3511 ), .A2(\unit_decode/n3491 ), .ZN(
        \unit_decode/n2940 ) );
  BUF_X1 U1915 ( .A(\unit_decode/RegisterFile/N445 ), .Z(n705) );
  BUF_X1 U1916 ( .A(\unit_decode/RegisterFile/N444 ), .Z(n708) );
  NAND4_X1 U1917 ( .A1(\unit_memory/DRAM/n837 ), .A2(\unit_memory/DRAM/n838 ), 
        .A3(\unit_memory/DRAM/n839 ), .A4(\unit_memory/DRAM/n840 ), .ZN(
        \unit_memory/DRAM/N596 ) );
  OAI21_X1 U1918 ( .B1(\unit_memory/DRAM/n854 ), .B2(\unit_memory/DRAM/n855 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n837 ) );
  OAI21_X1 U1919 ( .B1(\unit_memory/DRAM/n850 ), .B2(\unit_memory/DRAM/n851 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n838 ) );
  NAND4_X1 U1920 ( .A1(\unit_memory/DRAM/n811 ), .A2(\unit_memory/DRAM/n812 ), 
        .A3(\unit_memory/DRAM/n813 ), .A4(\unit_memory/DRAM/n814 ), .ZN(
        \unit_memory/DRAM/N597 ) );
  OAI21_X1 U1921 ( .B1(\unit_memory/DRAM/n832 ), .B2(\unit_memory/DRAM/n833 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n811 ) );
  OAI21_X1 U1922 ( .B1(\unit_memory/DRAM/n827 ), .B2(\unit_memory/DRAM/n828 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n812 ) );
  NAND4_X1 U1923 ( .A1(\unit_memory/DRAM/n858 ), .A2(\unit_memory/DRAM/n859 ), 
        .A3(\unit_memory/DRAM/n860 ), .A4(\unit_memory/DRAM/n861 ), .ZN(
        \unit_memory/DRAM/N595 ) );
  OAI21_X1 U1924 ( .B1(\unit_memory/DRAM/n875 ), .B2(\unit_memory/DRAM/n876 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n858 ) );
  OAI21_X1 U1925 ( .B1(\unit_memory/DRAM/n871 ), .B2(\unit_memory/DRAM/n872 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n859 ) );
  NAND4_X1 U1926 ( .A1(\unit_memory/DRAM/n879 ), .A2(\unit_memory/DRAM/n880 ), 
        .A3(\unit_memory/DRAM/n881 ), .A4(\unit_memory/DRAM/n882 ), .ZN(
        \unit_memory/DRAM/N594 ) );
  OAI21_X1 U1927 ( .B1(\unit_memory/DRAM/n896 ), .B2(\unit_memory/DRAM/n897 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n879 ) );
  OAI21_X1 U1928 ( .B1(\unit_memory/DRAM/n892 ), .B2(\unit_memory/DRAM/n893 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n880 ) );
  NAND4_X1 U1929 ( .A1(\unit_memory/DRAM/n900 ), .A2(\unit_memory/DRAM/n901 ), 
        .A3(\unit_memory/DRAM/n902 ), .A4(\unit_memory/DRAM/n903 ), .ZN(
        \unit_memory/DRAM/N593 ) );
  OAI21_X1 U1930 ( .B1(\unit_memory/DRAM/n917 ), .B2(\unit_memory/DRAM/n918 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n900 ) );
  OAI21_X1 U1931 ( .B1(\unit_memory/DRAM/n913 ), .B2(\unit_memory/DRAM/n914 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n901 ) );
  NAND4_X1 U1932 ( .A1(\unit_memory/DRAM/n921 ), .A2(\unit_memory/DRAM/n922 ), 
        .A3(\unit_memory/DRAM/n923 ), .A4(\unit_memory/DRAM/n924 ), .ZN(
        \unit_memory/DRAM/N592 ) );
  OAI21_X1 U1933 ( .B1(\unit_memory/DRAM/n938 ), .B2(\unit_memory/DRAM/n939 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n921 ) );
  OAI21_X1 U1934 ( .B1(\unit_memory/DRAM/n934 ), .B2(\unit_memory/DRAM/n935 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n922 ) );
  NAND4_X1 U1935 ( .A1(\unit_memory/DRAM/n942 ), .A2(\unit_memory/DRAM/n943 ), 
        .A3(\unit_memory/DRAM/n944 ), .A4(\unit_memory/DRAM/n945 ), .ZN(
        \unit_memory/DRAM/N591 ) );
  OAI21_X1 U1936 ( .B1(\unit_memory/DRAM/n959 ), .B2(\unit_memory/DRAM/n960 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n942 ) );
  OAI21_X1 U1937 ( .B1(\unit_memory/DRAM/n955 ), .B2(\unit_memory/DRAM/n956 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n943 ) );
  NAND4_X1 U1938 ( .A1(\unit_memory/DRAM/n963 ), .A2(\unit_memory/DRAM/n964 ), 
        .A3(\unit_memory/DRAM/n965 ), .A4(\unit_memory/DRAM/n966 ), .ZN(
        \unit_memory/DRAM/N590 ) );
  OAI21_X1 U1939 ( .B1(\unit_memory/DRAM/n980 ), .B2(\unit_memory/DRAM/n981 ), 
        .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n963 ) );
  OAI21_X1 U1940 ( .B1(\unit_memory/DRAM/n976 ), .B2(\unit_memory/DRAM/n977 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n964 ) );
  NAND4_X1 U1941 ( .A1(\unit_memory/DRAM/n984 ), .A2(\unit_memory/DRAM/n985 ), 
        .A3(\unit_memory/DRAM/n986 ), .A4(\unit_memory/DRAM/n987 ), .ZN(
        \unit_memory/DRAM/N589 ) );
  OAI21_X1 U1942 ( .B1(\unit_memory/DRAM/n1001 ), .B2(\unit_memory/DRAM/n1002 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n984 ) );
  OAI21_X1 U1943 ( .B1(\unit_memory/DRAM/n997 ), .B2(\unit_memory/DRAM/n998 ), 
        .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n985 ) );
  NAND4_X1 U1944 ( .A1(\unit_memory/DRAM/n1005 ), .A2(\unit_memory/DRAM/n1006 ), .A3(\unit_memory/DRAM/n1007 ), .A4(\unit_memory/DRAM/n1008 ), .ZN(
        \unit_memory/DRAM/N588 ) );
  OAI21_X1 U1945 ( .B1(\unit_memory/DRAM/n1022 ), .B2(\unit_memory/DRAM/n1023 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1005 ) );
  OAI21_X1 U1946 ( .B1(\unit_memory/DRAM/n1018 ), .B2(\unit_memory/DRAM/n1019 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1006 ) );
  NAND4_X1 U1947 ( .A1(\unit_memory/DRAM/n1026 ), .A2(\unit_memory/DRAM/n1027 ), .A3(\unit_memory/DRAM/n1028 ), .A4(\unit_memory/DRAM/n1029 ), .ZN(
        \unit_memory/DRAM/N587 ) );
  OAI21_X1 U1948 ( .B1(\unit_memory/DRAM/n1043 ), .B2(\unit_memory/DRAM/n1044 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1026 ) );
  OAI21_X1 U1949 ( .B1(\unit_memory/DRAM/n1039 ), .B2(\unit_memory/DRAM/n1040 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1027 ) );
  NAND4_X1 U1950 ( .A1(\unit_memory/DRAM/n1047 ), .A2(\unit_memory/DRAM/n1048 ), .A3(\unit_memory/DRAM/n1049 ), .A4(\unit_memory/DRAM/n1050 ), .ZN(
        \unit_memory/DRAM/N586 ) );
  OAI21_X1 U1951 ( .B1(\unit_memory/DRAM/n1064 ), .B2(\unit_memory/DRAM/n1065 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1047 ) );
  OAI21_X1 U1952 ( .B1(\unit_memory/DRAM/n1060 ), .B2(\unit_memory/DRAM/n1061 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1048 ) );
  NAND4_X1 U1953 ( .A1(\unit_memory/DRAM/n1068 ), .A2(\unit_memory/DRAM/n1069 ), .A3(\unit_memory/DRAM/n1070 ), .A4(\unit_memory/DRAM/n1071 ), .ZN(
        \unit_memory/DRAM/N585 ) );
  OAI21_X1 U1954 ( .B1(\unit_memory/DRAM/n1085 ), .B2(\unit_memory/DRAM/n1086 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1068 ) );
  OAI21_X1 U1955 ( .B1(\unit_memory/DRAM/n1081 ), .B2(\unit_memory/DRAM/n1082 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1069 ) );
  NAND4_X1 U1956 ( .A1(\unit_memory/DRAM/n1089 ), .A2(\unit_memory/DRAM/n1090 ), .A3(\unit_memory/DRAM/n1091 ), .A4(\unit_memory/DRAM/n1092 ), .ZN(
        \unit_memory/DRAM/N584 ) );
  OAI21_X1 U1957 ( .B1(\unit_memory/DRAM/n1106 ), .B2(\unit_memory/DRAM/n1107 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1089 ) );
  OAI21_X1 U1958 ( .B1(\unit_memory/DRAM/n1102 ), .B2(\unit_memory/DRAM/n1103 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1090 ) );
  NAND4_X1 U1959 ( .A1(\unit_memory/DRAM/n1110 ), .A2(\unit_memory/DRAM/n1111 ), .A3(\unit_memory/DRAM/n1112 ), .A4(\unit_memory/DRAM/n1113 ), .ZN(
        \unit_memory/DRAM/N583 ) );
  OAI21_X1 U1960 ( .B1(\unit_memory/DRAM/n1127 ), .B2(\unit_memory/DRAM/n1128 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1110 ) );
  OAI21_X1 U1961 ( .B1(\unit_memory/DRAM/n1123 ), .B2(\unit_memory/DRAM/n1124 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1111 ) );
  NAND4_X1 U1962 ( .A1(\unit_memory/DRAM/n1131 ), .A2(\unit_memory/DRAM/n1132 ), .A3(\unit_memory/DRAM/n1133 ), .A4(\unit_memory/DRAM/n1134 ), .ZN(
        \unit_memory/DRAM/N582 ) );
  OAI21_X1 U1963 ( .B1(\unit_memory/DRAM/n2195 ), .B2(\unit_memory/DRAM/n2196 ), .A(\unit_memory/DRAM/n834 ), .ZN(\unit_memory/DRAM/n1131 ) );
  OAI21_X1 U1964 ( .B1(\unit_memory/DRAM/n2191 ), .B2(\unit_memory/DRAM/n2192 ), .A(\unit_memory/DRAM/n829 ), .ZN(\unit_memory/DRAM/n1132 ) );
  NAND2_X1 U1965 ( .A1(\unit_memory/DRAM/n782 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n574 ) );
  NAND2_X1 U1966 ( .A1(\unit_memory/DRAM/n772 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n575 ) );
  AND4_X1 U1967 ( .A1(\unit_memory/DRAM/n1137 ), .A2(\unit_memory/DRAM/n1138 ), 
        .A3(\unit_memory/DRAM/n1139 ), .A4(\unit_memory/DRAM/n1140 ), .ZN(
        \unit_memory/DRAM/n561 ) );
  OAI21_X1 U1968 ( .B1(\unit_memory/DRAM/n1155 ), .B2(\unit_memory/DRAM/n1156 ), .A(\unit_memory/DRAM/n548 ), .ZN(\unit_memory/DRAM/n1137 ) );
  OAI21_X1 U1969 ( .B1(\unit_memory/DRAM/n1151 ), .B2(\unit_memory/DRAM/n1152 ), .A(\unit_memory/DRAM/n549 ), .ZN(\unit_memory/DRAM/n1138 ) );
  OAI21_X1 U1970 ( .B1(\unit_memory/DRAM/n1146 ), .B2(\unit_memory/DRAM/n1147 ), .A(\unit_memory/DRAM/n1148 ), .ZN(\unit_memory/DRAM/n1139 ) );
  NAND2_X1 U1971 ( .A1(\unit_decode/n2862 ), .A2(\unit_decode/n2863 ), .ZN(
        \unit_decode/RegisterFile/N412 ) );
  NOR4_X1 U1972 ( .A1(\unit_decode/n2880 ), .A2(\unit_decode/n2881 ), .A3(
        \unit_decode/n2882 ), .A4(\unit_decode/n2883 ), .ZN(
        \unit_decode/n2862 ) );
  NOR4_X1 U1973 ( .A1(\unit_decode/n2864 ), .A2(\unit_decode/n2865 ), .A3(
        \unit_decode/n2866 ), .A4(\unit_decode/n2867 ), .ZN(
        \unit_decode/n2863 ) );
  OAI221_X1 U1974 ( .B1(\unit_decode/n1293 ), .B2(n1177), .C1(
        \unit_decode/n1269 ), .C2(n1180), .A(\unit_decode/n2890 ), .ZN(
        \unit_decode/n2880 ) );
  NAND2_X1 U1975 ( .A1(\unit_decode/n2844 ), .A2(\unit_decode/n2845 ), .ZN(
        \unit_decode/RegisterFile/N413 ) );
  NOR4_X1 U1976 ( .A1(\unit_decode/n2854 ), .A2(\unit_decode/n2855 ), .A3(
        \unit_decode/n2856 ), .A4(\unit_decode/n2857 ), .ZN(
        \unit_decode/n2844 ) );
  NOR4_X1 U1977 ( .A1(\unit_decode/n2846 ), .A2(\unit_decode/n2847 ), .A3(
        \unit_decode/n2848 ), .A4(\unit_decode/n2849 ), .ZN(
        \unit_decode/n2845 ) );
  OAI221_X1 U1978 ( .B1(\unit_decode/n1294 ), .B2(n1177), .C1(
        \unit_decode/n1270 ), .C2(n1180), .A(\unit_decode/n2861 ), .ZN(
        \unit_decode/n2854 ) );
  NAND2_X1 U1979 ( .A1(\unit_decode/n2826 ), .A2(\unit_decode/n2827 ), .ZN(
        \unit_decode/RegisterFile/N414 ) );
  NOR4_X1 U1980 ( .A1(\unit_decode/n2836 ), .A2(\unit_decode/n2837 ), .A3(
        \unit_decode/n2838 ), .A4(\unit_decode/n2839 ), .ZN(
        \unit_decode/n2826 ) );
  NOR4_X1 U1981 ( .A1(\unit_decode/n2828 ), .A2(\unit_decode/n2829 ), .A3(
        \unit_decode/n2830 ), .A4(\unit_decode/n2831 ), .ZN(
        \unit_decode/n2827 ) );
  OAI221_X1 U1982 ( .B1(\unit_decode/n1295 ), .B2(n1177), .C1(
        \unit_decode/n1271 ), .C2(n1180), .A(\unit_decode/n2843 ), .ZN(
        \unit_decode/n2836 ) );
  NAND2_X1 U1983 ( .A1(\unit_decode/n2808 ), .A2(\unit_decode/n2809 ), .ZN(
        \unit_decode/RegisterFile/N415 ) );
  NOR4_X1 U1984 ( .A1(\unit_decode/n2818 ), .A2(\unit_decode/n2819 ), .A3(
        \unit_decode/n2820 ), .A4(\unit_decode/n2821 ), .ZN(
        \unit_decode/n2808 ) );
  NOR4_X1 U1985 ( .A1(\unit_decode/n2810 ), .A2(\unit_decode/n2811 ), .A3(
        \unit_decode/n2812 ), .A4(\unit_decode/n2813 ), .ZN(
        \unit_decode/n2809 ) );
  OAI221_X1 U1986 ( .B1(\unit_decode/n1296 ), .B2(n1177), .C1(
        \unit_decode/n1272 ), .C2(n1180), .A(\unit_decode/n2825 ), .ZN(
        \unit_decode/n2818 ) );
  NAND2_X1 U1987 ( .A1(\unit_decode/n2790 ), .A2(\unit_decode/n2791 ), .ZN(
        \unit_decode/RegisterFile/N416 ) );
  NOR4_X1 U1988 ( .A1(\unit_decode/n2800 ), .A2(\unit_decode/n2801 ), .A3(
        \unit_decode/n2802 ), .A4(\unit_decode/n2803 ), .ZN(
        \unit_decode/n2790 ) );
  NOR4_X1 U1989 ( .A1(\unit_decode/n2792 ), .A2(\unit_decode/n2793 ), .A3(
        \unit_decode/n2794 ), .A4(\unit_decode/n2795 ), .ZN(
        \unit_decode/n2791 ) );
  OAI221_X1 U1990 ( .B1(\unit_decode/n1297 ), .B2(n1177), .C1(
        \unit_decode/n1273 ), .C2(n1180), .A(\unit_decode/n2807 ), .ZN(
        \unit_decode/n2800 ) );
  NAND2_X1 U1991 ( .A1(\unit_decode/n2772 ), .A2(\unit_decode/n2773 ), .ZN(
        \unit_decode/RegisterFile/N417 ) );
  NOR4_X1 U1992 ( .A1(\unit_decode/n2782 ), .A2(\unit_decode/n2783 ), .A3(
        \unit_decode/n2784 ), .A4(\unit_decode/n2785 ), .ZN(
        \unit_decode/n2772 ) );
  NOR4_X1 U1993 ( .A1(\unit_decode/n2774 ), .A2(\unit_decode/n2775 ), .A3(
        \unit_decode/n2776 ), .A4(\unit_decode/n2777 ), .ZN(
        \unit_decode/n2773 ) );
  OAI221_X1 U1994 ( .B1(\unit_decode/n1298 ), .B2(n1177), .C1(
        \unit_decode/n1274 ), .C2(n1180), .A(\unit_decode/n2789 ), .ZN(
        \unit_decode/n2782 ) );
  NAND2_X1 U1995 ( .A1(\unit_decode/n2754 ), .A2(\unit_decode/n2755 ), .ZN(
        \unit_decode/RegisterFile/N418 ) );
  NOR4_X1 U1996 ( .A1(\unit_decode/n2764 ), .A2(\unit_decode/n2765 ), .A3(
        \unit_decode/n2766 ), .A4(\unit_decode/n2767 ), .ZN(
        \unit_decode/n2754 ) );
  NOR4_X1 U1997 ( .A1(\unit_decode/n2756 ), .A2(\unit_decode/n2757 ), .A3(
        \unit_decode/n2758 ), .A4(\unit_decode/n2759 ), .ZN(
        \unit_decode/n2755 ) );
  OAI221_X1 U1998 ( .B1(\unit_decode/n1299 ), .B2(n1177), .C1(
        \unit_decode/n1275 ), .C2(n1180), .A(\unit_decode/n2771 ), .ZN(
        \unit_decode/n2764 ) );
  NAND2_X1 U1999 ( .A1(\unit_decode/n2736 ), .A2(\unit_decode/n2737 ), .ZN(
        \unit_decode/RegisterFile/N419 ) );
  NOR4_X1 U2000 ( .A1(\unit_decode/n2746 ), .A2(\unit_decode/n2747 ), .A3(
        \unit_decode/n2748 ), .A4(\unit_decode/n2749 ), .ZN(
        \unit_decode/n2736 ) );
  NOR4_X1 U2001 ( .A1(\unit_decode/n2738 ), .A2(\unit_decode/n2739 ), .A3(
        \unit_decode/n2740 ), .A4(\unit_decode/n2741 ), .ZN(
        \unit_decode/n2737 ) );
  OAI221_X1 U2002 ( .B1(\unit_decode/n1300 ), .B2(n1177), .C1(
        \unit_decode/n1276 ), .C2(n1180), .A(\unit_decode/n2753 ), .ZN(
        \unit_decode/n2746 ) );
  NAND2_X1 U2003 ( .A1(\unit_decode/n2718 ), .A2(\unit_decode/n2719 ), .ZN(
        \unit_decode/RegisterFile/N420 ) );
  NOR4_X1 U2004 ( .A1(\unit_decode/n2728 ), .A2(\unit_decode/n2729 ), .A3(
        \unit_decode/n2730 ), .A4(\unit_decode/n2731 ), .ZN(
        \unit_decode/n2718 ) );
  NOR4_X1 U2005 ( .A1(\unit_decode/n2720 ), .A2(\unit_decode/n2721 ), .A3(
        \unit_decode/n2722 ), .A4(\unit_decode/n2723 ), .ZN(
        \unit_decode/n2719 ) );
  OAI221_X1 U2006 ( .B1(\unit_decode/n1301 ), .B2(n1177), .C1(
        \unit_decode/n1277 ), .C2(n1180), .A(\unit_decode/n2735 ), .ZN(
        \unit_decode/n2728 ) );
  NAND2_X1 U2007 ( .A1(\unit_decode/n2700 ), .A2(\unit_decode/n2701 ), .ZN(
        \unit_decode/RegisterFile/N421 ) );
  NOR4_X1 U2008 ( .A1(\unit_decode/n2710 ), .A2(\unit_decode/n2711 ), .A3(
        \unit_decode/n2712 ), .A4(\unit_decode/n2713 ), .ZN(
        \unit_decode/n2700 ) );
  NOR4_X1 U2009 ( .A1(\unit_decode/n2702 ), .A2(\unit_decode/n2703 ), .A3(
        \unit_decode/n2704 ), .A4(\unit_decode/n2705 ), .ZN(
        \unit_decode/n2701 ) );
  OAI221_X1 U2010 ( .B1(\unit_decode/n1302 ), .B2(n1177), .C1(
        \unit_decode/n1278 ), .C2(n1180), .A(\unit_decode/n2717 ), .ZN(
        \unit_decode/n2710 ) );
  NAND2_X1 U2011 ( .A1(\unit_decode/n2682 ), .A2(\unit_decode/n2683 ), .ZN(
        \unit_decode/RegisterFile/N422 ) );
  NOR4_X1 U2012 ( .A1(\unit_decode/n2692 ), .A2(\unit_decode/n2693 ), .A3(
        \unit_decode/n2694 ), .A4(\unit_decode/n2695 ), .ZN(
        \unit_decode/n2682 ) );
  NOR4_X1 U2013 ( .A1(\unit_decode/n2684 ), .A2(\unit_decode/n2685 ), .A3(
        \unit_decode/n2686 ), .A4(\unit_decode/n2687 ), .ZN(
        \unit_decode/n2683 ) );
  OAI221_X1 U2014 ( .B1(\unit_decode/n1303 ), .B2(n1177), .C1(
        \unit_decode/n1279 ), .C2(n1180), .A(\unit_decode/n2699 ), .ZN(
        \unit_decode/n2692 ) );
  NAND2_X1 U2015 ( .A1(\unit_decode/n2664 ), .A2(\unit_decode/n2665 ), .ZN(
        \unit_decode/RegisterFile/N423 ) );
  NOR4_X1 U2016 ( .A1(\unit_decode/n2674 ), .A2(\unit_decode/n2675 ), .A3(
        \unit_decode/n2676 ), .A4(\unit_decode/n2677 ), .ZN(
        \unit_decode/n2664 ) );
  NOR4_X1 U2017 ( .A1(\unit_decode/n2666 ), .A2(\unit_decode/n2667 ), .A3(
        \unit_decode/n2668 ), .A4(\unit_decode/n2669 ), .ZN(
        \unit_decode/n2665 ) );
  OAI221_X1 U2018 ( .B1(\unit_decode/n1304 ), .B2(n1177), .C1(
        \unit_decode/n1280 ), .C2(n1180), .A(\unit_decode/n2681 ), .ZN(
        \unit_decode/n2674 ) );
  NAND2_X1 U2019 ( .A1(\unit_decode/n2646 ), .A2(\unit_decode/n2647 ), .ZN(
        \unit_decode/RegisterFile/N424 ) );
  NOR4_X1 U2020 ( .A1(\unit_decode/n2656 ), .A2(\unit_decode/n2657 ), .A3(
        \unit_decode/n2658 ), .A4(\unit_decode/n2659 ), .ZN(
        \unit_decode/n2646 ) );
  NOR4_X1 U2021 ( .A1(\unit_decode/n2648 ), .A2(\unit_decode/n2649 ), .A3(
        \unit_decode/n2650 ), .A4(\unit_decode/n2651 ), .ZN(
        \unit_decode/n2647 ) );
  OAI221_X1 U2022 ( .B1(\unit_decode/n1305 ), .B2(n1178), .C1(
        \unit_decode/n1281 ), .C2(n1181), .A(\unit_decode/n2663 ), .ZN(
        \unit_decode/n2656 ) );
  NAND2_X1 U2023 ( .A1(\unit_decode/n2628 ), .A2(\unit_decode/n2629 ), .ZN(
        \unit_decode/RegisterFile/N425 ) );
  NOR4_X1 U2024 ( .A1(\unit_decode/n2638 ), .A2(\unit_decode/n2639 ), .A3(
        \unit_decode/n2640 ), .A4(\unit_decode/n2641 ), .ZN(
        \unit_decode/n2628 ) );
  NOR4_X1 U2025 ( .A1(\unit_decode/n2630 ), .A2(\unit_decode/n2631 ), .A3(
        \unit_decode/n2632 ), .A4(\unit_decode/n2633 ), .ZN(
        \unit_decode/n2629 ) );
  OAI221_X1 U2026 ( .B1(\unit_decode/n1306 ), .B2(n1178), .C1(
        \unit_decode/n1282 ), .C2(n1181), .A(\unit_decode/n2645 ), .ZN(
        \unit_decode/n2638 ) );
  NAND2_X1 U2027 ( .A1(\unit_decode/n2610 ), .A2(\unit_decode/n2611 ), .ZN(
        \unit_decode/RegisterFile/N426 ) );
  NOR4_X1 U2028 ( .A1(\unit_decode/n2620 ), .A2(\unit_decode/n2621 ), .A3(
        \unit_decode/n2622 ), .A4(\unit_decode/n2623 ), .ZN(
        \unit_decode/n2610 ) );
  NOR4_X1 U2029 ( .A1(\unit_decode/n2612 ), .A2(\unit_decode/n2613 ), .A3(
        \unit_decode/n2614 ), .A4(\unit_decode/n2615 ), .ZN(
        \unit_decode/n2611 ) );
  OAI221_X1 U2030 ( .B1(\unit_decode/n1307 ), .B2(n1178), .C1(
        \unit_decode/n1283 ), .C2(n1181), .A(\unit_decode/n2627 ), .ZN(
        \unit_decode/n2620 ) );
  NAND2_X1 U2031 ( .A1(\unit_decode/n2592 ), .A2(\unit_decode/n2593 ), .ZN(
        \unit_decode/RegisterFile/N427 ) );
  NOR4_X1 U2032 ( .A1(\unit_decode/n2602 ), .A2(\unit_decode/n2603 ), .A3(
        \unit_decode/n2604 ), .A4(\unit_decode/n2605 ), .ZN(
        \unit_decode/n2592 ) );
  NOR4_X1 U2033 ( .A1(\unit_decode/n2594 ), .A2(\unit_decode/n2595 ), .A3(
        \unit_decode/n2596 ), .A4(\unit_decode/n2597 ), .ZN(
        \unit_decode/n2593 ) );
  OAI221_X1 U2034 ( .B1(\unit_decode/n1308 ), .B2(n1178), .C1(
        \unit_decode/n1284 ), .C2(n1181), .A(\unit_decode/n2609 ), .ZN(
        \unit_decode/n2602 ) );
  NAND2_X1 U2035 ( .A1(\unit_decode/n2574 ), .A2(\unit_decode/n2575 ), .ZN(
        \unit_decode/RegisterFile/N428 ) );
  NOR4_X1 U2036 ( .A1(\unit_decode/n2584 ), .A2(\unit_decode/n2585 ), .A3(
        \unit_decode/n2586 ), .A4(\unit_decode/n2587 ), .ZN(
        \unit_decode/n2574 ) );
  NOR4_X1 U2037 ( .A1(\unit_decode/n2576 ), .A2(\unit_decode/n2577 ), .A3(
        \unit_decode/n2578 ), .A4(\unit_decode/n2579 ), .ZN(
        \unit_decode/n2575 ) );
  OAI221_X1 U2038 ( .B1(\unit_decode/n1309 ), .B2(n1178), .C1(
        \unit_decode/n1285 ), .C2(n1181), .A(\unit_decode/n2591 ), .ZN(
        \unit_decode/n2584 ) );
  NAND2_X1 U2039 ( .A1(\unit_decode/n2556 ), .A2(\unit_decode/n2557 ), .ZN(
        \unit_decode/RegisterFile/N429 ) );
  NOR4_X1 U2040 ( .A1(\unit_decode/n2566 ), .A2(\unit_decode/n2567 ), .A3(
        \unit_decode/n2568 ), .A4(\unit_decode/n2569 ), .ZN(
        \unit_decode/n2556 ) );
  NOR4_X1 U2041 ( .A1(\unit_decode/n2558 ), .A2(\unit_decode/n2559 ), .A3(
        \unit_decode/n2560 ), .A4(\unit_decode/n2561 ), .ZN(
        \unit_decode/n2557 ) );
  OAI221_X1 U2042 ( .B1(\unit_decode/n1310 ), .B2(n1178), .C1(
        \unit_decode/n1286 ), .C2(n1181), .A(\unit_decode/n2573 ), .ZN(
        \unit_decode/n2566 ) );
  NAND2_X1 U2043 ( .A1(\unit_decode/n2538 ), .A2(\unit_decode/n2539 ), .ZN(
        \unit_decode/RegisterFile/N430 ) );
  NOR4_X1 U2044 ( .A1(\unit_decode/n2548 ), .A2(\unit_decode/n2549 ), .A3(
        \unit_decode/n2550 ), .A4(\unit_decode/n2551 ), .ZN(
        \unit_decode/n2538 ) );
  NOR4_X1 U2045 ( .A1(\unit_decode/n2540 ), .A2(\unit_decode/n2541 ), .A3(
        \unit_decode/n2542 ), .A4(\unit_decode/n2543 ), .ZN(
        \unit_decode/n2539 ) );
  OAI221_X1 U2046 ( .B1(\unit_decode/n1311 ), .B2(n1178), .C1(
        \unit_decode/n1287 ), .C2(n1181), .A(\unit_decode/n2555 ), .ZN(
        \unit_decode/n2548 ) );
  NAND2_X1 U2047 ( .A1(\unit_decode/n2520 ), .A2(\unit_decode/n2521 ), .ZN(
        \unit_decode/RegisterFile/N431 ) );
  NOR4_X1 U2048 ( .A1(\unit_decode/n2530 ), .A2(\unit_decode/n2531 ), .A3(
        \unit_decode/n2532 ), .A4(\unit_decode/n2533 ), .ZN(
        \unit_decode/n2520 ) );
  NOR4_X1 U2049 ( .A1(\unit_decode/n2522 ), .A2(\unit_decode/n2523 ), .A3(
        \unit_decode/n2524 ), .A4(\unit_decode/n2525 ), .ZN(
        \unit_decode/n2521 ) );
  OAI221_X1 U2050 ( .B1(\unit_decode/n1312 ), .B2(n1178), .C1(
        \unit_decode/n1288 ), .C2(n1181), .A(\unit_decode/n2537 ), .ZN(
        \unit_decode/n2530 ) );
  NAND2_X1 U2051 ( .A1(\unit_decode/n2502 ), .A2(\unit_decode/n2503 ), .ZN(
        \unit_decode/RegisterFile/N432 ) );
  NOR4_X1 U2052 ( .A1(\unit_decode/n2512 ), .A2(\unit_decode/n2513 ), .A3(
        \unit_decode/n2514 ), .A4(\unit_decode/n2515 ), .ZN(
        \unit_decode/n2502 ) );
  NOR4_X1 U2053 ( .A1(\unit_decode/n2504 ), .A2(\unit_decode/n2505 ), .A3(
        \unit_decode/n2506 ), .A4(\unit_decode/n2507 ), .ZN(
        \unit_decode/n2503 ) );
  OAI221_X1 U2054 ( .B1(\unit_decode/n1313 ), .B2(n1178), .C1(
        \unit_decode/n1289 ), .C2(n1181), .A(\unit_decode/n2519 ), .ZN(
        \unit_decode/n2512 ) );
  NAND2_X1 U2055 ( .A1(\unit_decode/n2484 ), .A2(\unit_decode/n2485 ), .ZN(
        \unit_decode/RegisterFile/N433 ) );
  NOR4_X1 U2056 ( .A1(\unit_decode/n2494 ), .A2(\unit_decode/n2495 ), .A3(
        \unit_decode/n2496 ), .A4(\unit_decode/n2497 ), .ZN(
        \unit_decode/n2484 ) );
  NOR4_X1 U2057 ( .A1(\unit_decode/n2486 ), .A2(\unit_decode/n2487 ), .A3(
        \unit_decode/n2488 ), .A4(\unit_decode/n2489 ), .ZN(
        \unit_decode/n2485 ) );
  OAI221_X1 U2058 ( .B1(\unit_decode/n1314 ), .B2(n1178), .C1(
        \unit_decode/n1290 ), .C2(n1181), .A(\unit_decode/n2501 ), .ZN(
        \unit_decode/n2494 ) );
  NAND2_X1 U2059 ( .A1(\unit_decode/n2466 ), .A2(\unit_decode/n2467 ), .ZN(
        \unit_decode/RegisterFile/N434 ) );
  NOR4_X1 U2060 ( .A1(\unit_decode/n2476 ), .A2(\unit_decode/n2477 ), .A3(
        \unit_decode/n2478 ), .A4(\unit_decode/n2479 ), .ZN(
        \unit_decode/n2466 ) );
  NOR4_X1 U2061 ( .A1(\unit_decode/n2468 ), .A2(\unit_decode/n2469 ), .A3(
        \unit_decode/n2470 ), .A4(\unit_decode/n2471 ), .ZN(
        \unit_decode/n2467 ) );
  OAI221_X1 U2062 ( .B1(\unit_decode/n1315 ), .B2(n1178), .C1(
        \unit_decode/n1291 ), .C2(n1181), .A(\unit_decode/n2483 ), .ZN(
        \unit_decode/n2476 ) );
  NAND2_X1 U2063 ( .A1(\unit_decode/n2448 ), .A2(\unit_decode/n2449 ), .ZN(
        \unit_decode/RegisterFile/N435 ) );
  NOR4_X1 U2064 ( .A1(\unit_decode/n2458 ), .A2(\unit_decode/n2459 ), .A3(
        \unit_decode/n2460 ), .A4(\unit_decode/n2461 ), .ZN(
        \unit_decode/n2448 ) );
  NOR4_X1 U2065 ( .A1(\unit_decode/n2450 ), .A2(\unit_decode/n2451 ), .A3(
        \unit_decode/n2452 ), .A4(\unit_decode/n2453 ), .ZN(
        \unit_decode/n2449 ) );
  OAI221_X1 U2066 ( .B1(\unit_decode/n1316 ), .B2(n1178), .C1(
        \unit_decode/n1292 ), .C2(n1181), .A(\unit_decode/n2465 ), .ZN(
        \unit_decode/n2458 ) );
  NAND2_X1 U2067 ( .A1(\unit_decode/n3482 ), .A2(\unit_decode/n3483 ), .ZN(
        \unit_decode/RegisterFile/N379 ) );
  NOR4_X1 U2068 ( .A1(\unit_decode/n3500 ), .A2(\unit_decode/n3501 ), .A3(
        \unit_decode/n3502 ), .A4(\unit_decode/n3503 ), .ZN(
        \unit_decode/n3482 ) );
  NOR4_X1 U2069 ( .A1(\unit_decode/n3484 ), .A2(\unit_decode/n3485 ), .A3(
        \unit_decode/n3486 ), .A4(\unit_decode/n3487 ), .ZN(
        \unit_decode/n3483 ) );
  OAI221_X1 U2070 ( .B1(\unit_decode/n1293 ), .B2(n1273), .C1(
        \unit_decode/n1269 ), .C2(n1276), .A(\unit_decode/n3510 ), .ZN(
        \unit_decode/n3500 ) );
  NAND2_X1 U2071 ( .A1(\unit_decode/n3464 ), .A2(\unit_decode/n3465 ), .ZN(
        \unit_decode/RegisterFile/N380 ) );
  NOR4_X1 U2072 ( .A1(\unit_decode/n3474 ), .A2(\unit_decode/n3475 ), .A3(
        \unit_decode/n3476 ), .A4(\unit_decode/n3477 ), .ZN(
        \unit_decode/n3464 ) );
  NOR4_X1 U2073 ( .A1(\unit_decode/n3466 ), .A2(\unit_decode/n3467 ), .A3(
        \unit_decode/n3468 ), .A4(\unit_decode/n3469 ), .ZN(
        \unit_decode/n3465 ) );
  OAI221_X1 U2074 ( .B1(\unit_decode/n1294 ), .B2(n1273), .C1(
        \unit_decode/n1270 ), .C2(n1276), .A(\unit_decode/n3481 ), .ZN(
        \unit_decode/n3474 ) );
  NAND2_X1 U2075 ( .A1(\unit_decode/n3446 ), .A2(\unit_decode/n3447 ), .ZN(
        \unit_decode/RegisterFile/N381 ) );
  NOR4_X1 U2076 ( .A1(\unit_decode/n3456 ), .A2(\unit_decode/n3457 ), .A3(
        \unit_decode/n3458 ), .A4(\unit_decode/n3459 ), .ZN(
        \unit_decode/n3446 ) );
  NOR4_X1 U2077 ( .A1(\unit_decode/n3448 ), .A2(\unit_decode/n3449 ), .A3(
        \unit_decode/n3450 ), .A4(\unit_decode/n3451 ), .ZN(
        \unit_decode/n3447 ) );
  OAI221_X1 U2078 ( .B1(\unit_decode/n1295 ), .B2(n1273), .C1(
        \unit_decode/n1271 ), .C2(n1276), .A(\unit_decode/n3463 ), .ZN(
        \unit_decode/n3456 ) );
  NAND2_X1 U2079 ( .A1(\unit_decode/n3428 ), .A2(\unit_decode/n3429 ), .ZN(
        \unit_decode/RegisterFile/N382 ) );
  NOR4_X1 U2080 ( .A1(\unit_decode/n3438 ), .A2(\unit_decode/n3439 ), .A3(
        \unit_decode/n3440 ), .A4(\unit_decode/n3441 ), .ZN(
        \unit_decode/n3428 ) );
  NOR4_X1 U2081 ( .A1(\unit_decode/n3430 ), .A2(\unit_decode/n3431 ), .A3(
        \unit_decode/n3432 ), .A4(\unit_decode/n3433 ), .ZN(
        \unit_decode/n3429 ) );
  OAI221_X1 U2082 ( .B1(\unit_decode/n1296 ), .B2(n1273), .C1(
        \unit_decode/n1272 ), .C2(n1276), .A(\unit_decode/n3445 ), .ZN(
        \unit_decode/n3438 ) );
  NAND2_X1 U2083 ( .A1(\unit_decode/n3410 ), .A2(\unit_decode/n3411 ), .ZN(
        \unit_decode/RegisterFile/N383 ) );
  NOR4_X1 U2084 ( .A1(\unit_decode/n3420 ), .A2(\unit_decode/n3421 ), .A3(
        \unit_decode/n3422 ), .A4(\unit_decode/n3423 ), .ZN(
        \unit_decode/n3410 ) );
  NOR4_X1 U2085 ( .A1(\unit_decode/n3412 ), .A2(\unit_decode/n3413 ), .A3(
        \unit_decode/n3414 ), .A4(\unit_decode/n3415 ), .ZN(
        \unit_decode/n3411 ) );
  OAI221_X1 U2086 ( .B1(\unit_decode/n1297 ), .B2(n1273), .C1(
        \unit_decode/n1273 ), .C2(n1276), .A(\unit_decode/n3427 ), .ZN(
        \unit_decode/n3420 ) );
  NAND2_X1 U2087 ( .A1(\unit_decode/n3392 ), .A2(\unit_decode/n3393 ), .ZN(
        \unit_decode/RegisterFile/N384 ) );
  NOR4_X1 U2088 ( .A1(\unit_decode/n3402 ), .A2(\unit_decode/n3403 ), .A3(
        \unit_decode/n3404 ), .A4(\unit_decode/n3405 ), .ZN(
        \unit_decode/n3392 ) );
  NOR4_X1 U2089 ( .A1(\unit_decode/n3394 ), .A2(\unit_decode/n3395 ), .A3(
        \unit_decode/n3396 ), .A4(\unit_decode/n3397 ), .ZN(
        \unit_decode/n3393 ) );
  OAI221_X1 U2090 ( .B1(\unit_decode/n1298 ), .B2(n1273), .C1(
        \unit_decode/n1274 ), .C2(n1276), .A(\unit_decode/n3409 ), .ZN(
        \unit_decode/n3402 ) );
  NAND2_X1 U2091 ( .A1(\unit_decode/n3374 ), .A2(\unit_decode/n3375 ), .ZN(
        \unit_decode/RegisterFile/N385 ) );
  NOR4_X1 U2092 ( .A1(\unit_decode/n3384 ), .A2(\unit_decode/n3385 ), .A3(
        \unit_decode/n3386 ), .A4(\unit_decode/n3387 ), .ZN(
        \unit_decode/n3374 ) );
  NOR4_X1 U2093 ( .A1(\unit_decode/n3376 ), .A2(\unit_decode/n3377 ), .A3(
        \unit_decode/n3378 ), .A4(\unit_decode/n3379 ), .ZN(
        \unit_decode/n3375 ) );
  OAI221_X1 U2094 ( .B1(\unit_decode/n1299 ), .B2(n1273), .C1(
        \unit_decode/n1275 ), .C2(n1276), .A(\unit_decode/n3391 ), .ZN(
        \unit_decode/n3384 ) );
  NAND2_X1 U2095 ( .A1(\unit_decode/n3356 ), .A2(\unit_decode/n3357 ), .ZN(
        \unit_decode/RegisterFile/N386 ) );
  NOR4_X1 U2096 ( .A1(\unit_decode/n3366 ), .A2(\unit_decode/n3367 ), .A3(
        \unit_decode/n3368 ), .A4(\unit_decode/n3369 ), .ZN(
        \unit_decode/n3356 ) );
  NOR4_X1 U2097 ( .A1(\unit_decode/n3358 ), .A2(\unit_decode/n3359 ), .A3(
        \unit_decode/n3360 ), .A4(\unit_decode/n3361 ), .ZN(
        \unit_decode/n3357 ) );
  OAI221_X1 U2098 ( .B1(\unit_decode/n1300 ), .B2(n1273), .C1(
        \unit_decode/n1276 ), .C2(n1276), .A(\unit_decode/n3373 ), .ZN(
        \unit_decode/n3366 ) );
  NAND2_X1 U2099 ( .A1(\unit_decode/n3338 ), .A2(\unit_decode/n3339 ), .ZN(
        \unit_decode/RegisterFile/N387 ) );
  NOR4_X1 U2100 ( .A1(\unit_decode/n3348 ), .A2(\unit_decode/n3349 ), .A3(
        \unit_decode/n3350 ), .A4(\unit_decode/n3351 ), .ZN(
        \unit_decode/n3338 ) );
  NOR4_X1 U2101 ( .A1(\unit_decode/n3340 ), .A2(\unit_decode/n3341 ), .A3(
        \unit_decode/n3342 ), .A4(\unit_decode/n3343 ), .ZN(
        \unit_decode/n3339 ) );
  OAI221_X1 U2102 ( .B1(\unit_decode/n1301 ), .B2(n1273), .C1(
        \unit_decode/n1277 ), .C2(n1276), .A(\unit_decode/n3355 ), .ZN(
        \unit_decode/n3348 ) );
  NAND2_X1 U2103 ( .A1(\unit_decode/n3320 ), .A2(\unit_decode/n3321 ), .ZN(
        \unit_decode/RegisterFile/N388 ) );
  NOR4_X1 U2104 ( .A1(\unit_decode/n3330 ), .A2(\unit_decode/n3331 ), .A3(
        \unit_decode/n3332 ), .A4(\unit_decode/n3333 ), .ZN(
        \unit_decode/n3320 ) );
  NOR4_X1 U2105 ( .A1(\unit_decode/n3322 ), .A2(\unit_decode/n3323 ), .A3(
        \unit_decode/n3324 ), .A4(\unit_decode/n3325 ), .ZN(
        \unit_decode/n3321 ) );
  OAI221_X1 U2106 ( .B1(\unit_decode/n1302 ), .B2(n1273), .C1(
        \unit_decode/n1278 ), .C2(n1276), .A(\unit_decode/n3337 ), .ZN(
        \unit_decode/n3330 ) );
  NAND2_X1 U2107 ( .A1(\unit_decode/n3302 ), .A2(\unit_decode/n3303 ), .ZN(
        \unit_decode/RegisterFile/N389 ) );
  NOR4_X1 U2108 ( .A1(\unit_decode/n3312 ), .A2(\unit_decode/n3313 ), .A3(
        \unit_decode/n3314 ), .A4(\unit_decode/n3315 ), .ZN(
        \unit_decode/n3302 ) );
  NOR4_X1 U2109 ( .A1(\unit_decode/n3304 ), .A2(\unit_decode/n3305 ), .A3(
        \unit_decode/n3306 ), .A4(\unit_decode/n3307 ), .ZN(
        \unit_decode/n3303 ) );
  OAI221_X1 U2110 ( .B1(\unit_decode/n1303 ), .B2(n1273), .C1(
        \unit_decode/n1279 ), .C2(n1276), .A(\unit_decode/n3319 ), .ZN(
        \unit_decode/n3312 ) );
  NAND2_X1 U2111 ( .A1(\unit_decode/n3284 ), .A2(\unit_decode/n3285 ), .ZN(
        \unit_decode/RegisterFile/N390 ) );
  NOR4_X1 U2112 ( .A1(\unit_decode/n3294 ), .A2(\unit_decode/n3295 ), .A3(
        \unit_decode/n3296 ), .A4(\unit_decode/n3297 ), .ZN(
        \unit_decode/n3284 ) );
  NOR4_X1 U2113 ( .A1(\unit_decode/n3286 ), .A2(\unit_decode/n3287 ), .A3(
        \unit_decode/n3288 ), .A4(\unit_decode/n3289 ), .ZN(
        \unit_decode/n3285 ) );
  OAI221_X1 U2114 ( .B1(\unit_decode/n1304 ), .B2(n1273), .C1(
        \unit_decode/n1280 ), .C2(n1276), .A(\unit_decode/n3301 ), .ZN(
        \unit_decode/n3294 ) );
  NAND2_X1 U2115 ( .A1(\unit_decode/n3266 ), .A2(\unit_decode/n3267 ), .ZN(
        \unit_decode/RegisterFile/N391 ) );
  NOR4_X1 U2116 ( .A1(\unit_decode/n3276 ), .A2(\unit_decode/n3277 ), .A3(
        \unit_decode/n3278 ), .A4(\unit_decode/n3279 ), .ZN(
        \unit_decode/n3266 ) );
  NOR4_X1 U2117 ( .A1(\unit_decode/n3268 ), .A2(\unit_decode/n3269 ), .A3(
        \unit_decode/n3270 ), .A4(\unit_decode/n3271 ), .ZN(
        \unit_decode/n3267 ) );
  OAI221_X1 U2118 ( .B1(\unit_decode/n1305 ), .B2(n1274), .C1(
        \unit_decode/n1281 ), .C2(n1277), .A(\unit_decode/n3283 ), .ZN(
        \unit_decode/n3276 ) );
  NAND2_X1 U2119 ( .A1(\unit_decode/n3248 ), .A2(\unit_decode/n3249 ), .ZN(
        \unit_decode/RegisterFile/N392 ) );
  NOR4_X1 U2120 ( .A1(\unit_decode/n3258 ), .A2(\unit_decode/n3259 ), .A3(
        \unit_decode/n3260 ), .A4(\unit_decode/n3261 ), .ZN(
        \unit_decode/n3248 ) );
  NOR4_X1 U2121 ( .A1(\unit_decode/n3250 ), .A2(\unit_decode/n3251 ), .A3(
        \unit_decode/n3252 ), .A4(\unit_decode/n3253 ), .ZN(
        \unit_decode/n3249 ) );
  OAI221_X1 U2122 ( .B1(\unit_decode/n1306 ), .B2(n1274), .C1(
        \unit_decode/n1282 ), .C2(n1277), .A(\unit_decode/n3265 ), .ZN(
        \unit_decode/n3258 ) );
  NAND2_X1 U2123 ( .A1(\unit_decode/n3230 ), .A2(\unit_decode/n3231 ), .ZN(
        \unit_decode/RegisterFile/N393 ) );
  NOR4_X1 U2124 ( .A1(\unit_decode/n3240 ), .A2(\unit_decode/n3241 ), .A3(
        \unit_decode/n3242 ), .A4(\unit_decode/n3243 ), .ZN(
        \unit_decode/n3230 ) );
  NOR4_X1 U2125 ( .A1(\unit_decode/n3232 ), .A2(\unit_decode/n3233 ), .A3(
        \unit_decode/n3234 ), .A4(\unit_decode/n3235 ), .ZN(
        \unit_decode/n3231 ) );
  OAI221_X1 U2126 ( .B1(\unit_decode/n1307 ), .B2(n1274), .C1(
        \unit_decode/n1283 ), .C2(n1277), .A(\unit_decode/n3247 ), .ZN(
        \unit_decode/n3240 ) );
  NAND2_X1 U2127 ( .A1(\unit_decode/n3212 ), .A2(\unit_decode/n3213 ), .ZN(
        \unit_decode/RegisterFile/N394 ) );
  NOR4_X1 U2128 ( .A1(\unit_decode/n3222 ), .A2(\unit_decode/n3223 ), .A3(
        \unit_decode/n3224 ), .A4(\unit_decode/n3225 ), .ZN(
        \unit_decode/n3212 ) );
  NOR4_X1 U2129 ( .A1(\unit_decode/n3214 ), .A2(\unit_decode/n3215 ), .A3(
        \unit_decode/n3216 ), .A4(\unit_decode/n3217 ), .ZN(
        \unit_decode/n3213 ) );
  OAI221_X1 U2130 ( .B1(\unit_decode/n1308 ), .B2(n1274), .C1(
        \unit_decode/n1284 ), .C2(n1277), .A(\unit_decode/n3229 ), .ZN(
        \unit_decode/n3222 ) );
  NAND2_X1 U2131 ( .A1(\unit_decode/n3194 ), .A2(\unit_decode/n3195 ), .ZN(
        \unit_decode/RegisterFile/N395 ) );
  NOR4_X1 U2132 ( .A1(\unit_decode/n3204 ), .A2(\unit_decode/n3205 ), .A3(
        \unit_decode/n3206 ), .A4(\unit_decode/n3207 ), .ZN(
        \unit_decode/n3194 ) );
  NOR4_X1 U2133 ( .A1(\unit_decode/n3196 ), .A2(\unit_decode/n3197 ), .A3(
        \unit_decode/n3198 ), .A4(\unit_decode/n3199 ), .ZN(
        \unit_decode/n3195 ) );
  OAI221_X1 U2134 ( .B1(\unit_decode/n1309 ), .B2(n1274), .C1(
        \unit_decode/n1285 ), .C2(n1277), .A(\unit_decode/n3211 ), .ZN(
        \unit_decode/n3204 ) );
  NAND2_X1 U2135 ( .A1(\unit_decode/n3176 ), .A2(\unit_decode/n3177 ), .ZN(
        \unit_decode/RegisterFile/N396 ) );
  NOR4_X1 U2136 ( .A1(\unit_decode/n3186 ), .A2(\unit_decode/n3187 ), .A3(
        \unit_decode/n3188 ), .A4(\unit_decode/n3189 ), .ZN(
        \unit_decode/n3176 ) );
  NOR4_X1 U2137 ( .A1(\unit_decode/n3178 ), .A2(\unit_decode/n3179 ), .A3(
        \unit_decode/n3180 ), .A4(\unit_decode/n3181 ), .ZN(
        \unit_decode/n3177 ) );
  OAI221_X1 U2138 ( .B1(\unit_decode/n1310 ), .B2(n1274), .C1(
        \unit_decode/n1286 ), .C2(n1277), .A(\unit_decode/n3193 ), .ZN(
        \unit_decode/n3186 ) );
  NAND2_X1 U2139 ( .A1(\unit_decode/n3158 ), .A2(\unit_decode/n3159 ), .ZN(
        \unit_decode/RegisterFile/N397 ) );
  NOR4_X1 U2140 ( .A1(\unit_decode/n3168 ), .A2(\unit_decode/n3169 ), .A3(
        \unit_decode/n3170 ), .A4(\unit_decode/n3171 ), .ZN(
        \unit_decode/n3158 ) );
  NOR4_X1 U2141 ( .A1(\unit_decode/n3160 ), .A2(\unit_decode/n3161 ), .A3(
        \unit_decode/n3162 ), .A4(\unit_decode/n3163 ), .ZN(
        \unit_decode/n3159 ) );
  OAI221_X1 U2142 ( .B1(\unit_decode/n1311 ), .B2(n1274), .C1(
        \unit_decode/n1287 ), .C2(n1277), .A(\unit_decode/n3175 ), .ZN(
        \unit_decode/n3168 ) );
  NAND2_X1 U2143 ( .A1(\unit_decode/n3140 ), .A2(\unit_decode/n3141 ), .ZN(
        \unit_decode/RegisterFile/N398 ) );
  NOR4_X1 U2144 ( .A1(\unit_decode/n3150 ), .A2(\unit_decode/n3151 ), .A3(
        \unit_decode/n3152 ), .A4(\unit_decode/n3153 ), .ZN(
        \unit_decode/n3140 ) );
  NOR4_X1 U2145 ( .A1(\unit_decode/n3142 ), .A2(\unit_decode/n3143 ), .A3(
        \unit_decode/n3144 ), .A4(\unit_decode/n3145 ), .ZN(
        \unit_decode/n3141 ) );
  OAI221_X1 U2146 ( .B1(\unit_decode/n1312 ), .B2(n1274), .C1(
        \unit_decode/n1288 ), .C2(n1277), .A(\unit_decode/n3157 ), .ZN(
        \unit_decode/n3150 ) );
  NAND2_X1 U2147 ( .A1(\unit_decode/n3122 ), .A2(\unit_decode/n3123 ), .ZN(
        \unit_decode/RegisterFile/N399 ) );
  NOR4_X1 U2148 ( .A1(\unit_decode/n3132 ), .A2(\unit_decode/n3133 ), .A3(
        \unit_decode/n3134 ), .A4(\unit_decode/n3135 ), .ZN(
        \unit_decode/n3122 ) );
  NOR4_X1 U2149 ( .A1(\unit_decode/n3124 ), .A2(\unit_decode/n3125 ), .A3(
        \unit_decode/n3126 ), .A4(\unit_decode/n3127 ), .ZN(
        \unit_decode/n3123 ) );
  OAI221_X1 U2150 ( .B1(\unit_decode/n1313 ), .B2(n1274), .C1(
        \unit_decode/n1289 ), .C2(n1277), .A(\unit_decode/n3139 ), .ZN(
        \unit_decode/n3132 ) );
  NAND2_X1 U2151 ( .A1(\unit_decode/n3104 ), .A2(\unit_decode/n3105 ), .ZN(
        \unit_decode/RegisterFile/N400 ) );
  NOR4_X1 U2152 ( .A1(\unit_decode/n3114 ), .A2(\unit_decode/n3115 ), .A3(
        \unit_decode/n3116 ), .A4(\unit_decode/n3117 ), .ZN(
        \unit_decode/n3104 ) );
  NOR4_X1 U2153 ( .A1(\unit_decode/n3106 ), .A2(\unit_decode/n3107 ), .A3(
        \unit_decode/n3108 ), .A4(\unit_decode/n3109 ), .ZN(
        \unit_decode/n3105 ) );
  OAI221_X1 U2154 ( .B1(\unit_decode/n1314 ), .B2(n1274), .C1(
        \unit_decode/n1290 ), .C2(n1277), .A(\unit_decode/n3121 ), .ZN(
        \unit_decode/n3114 ) );
  NAND2_X1 U2155 ( .A1(\unit_decode/n3086 ), .A2(\unit_decode/n3087 ), .ZN(
        \unit_decode/RegisterFile/N401 ) );
  NOR4_X1 U2156 ( .A1(\unit_decode/n3096 ), .A2(\unit_decode/n3097 ), .A3(
        \unit_decode/n3098 ), .A4(\unit_decode/n3099 ), .ZN(
        \unit_decode/n3086 ) );
  NOR4_X1 U2157 ( .A1(\unit_decode/n3088 ), .A2(\unit_decode/n3089 ), .A3(
        \unit_decode/n3090 ), .A4(\unit_decode/n3091 ), .ZN(
        \unit_decode/n3087 ) );
  OAI221_X1 U2158 ( .B1(\unit_decode/n1315 ), .B2(n1274), .C1(
        \unit_decode/n1291 ), .C2(n1277), .A(\unit_decode/n3103 ), .ZN(
        \unit_decode/n3096 ) );
  NAND2_X1 U2159 ( .A1(\unit_decode/n3068 ), .A2(\unit_decode/n3069 ), .ZN(
        \unit_decode/RegisterFile/N402 ) );
  NOR4_X1 U2160 ( .A1(\unit_decode/n3078 ), .A2(\unit_decode/n3079 ), .A3(
        \unit_decode/n3080 ), .A4(\unit_decode/n3081 ), .ZN(
        \unit_decode/n3068 ) );
  NOR4_X1 U2161 ( .A1(\unit_decode/n3070 ), .A2(\unit_decode/n3071 ), .A3(
        \unit_decode/n3072 ), .A4(\unit_decode/n3073 ), .ZN(
        \unit_decode/n3069 ) );
  OAI221_X1 U2162 ( .B1(\unit_decode/n1316 ), .B2(n1274), .C1(
        \unit_decode/n1292 ), .C2(n1277), .A(\unit_decode/n3085 ), .ZN(
        \unit_decode/n3078 ) );
  AND2_X1 U2163 ( .A1(\unit_memory/DRAM/n792 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n571 ) );
  AND2_X1 U2164 ( .A1(\unit_memory/DRAM/n809 ), .A2(\unit_memory/DRAM/n547 ), 
        .ZN(\unit_memory/DRAM/n572 ) );
  BUF_X1 U2165 ( .A(n1342), .Z(n1340) );
  BUF_X1 U2166 ( .A(n1343), .Z(n1338) );
  BUF_X1 U2167 ( .A(n1343), .Z(n1337) );
  BUF_X1 U2168 ( .A(n1342), .Z(n1339) );
  BUF_X1 U2169 ( .A(n1344), .Z(n1336) );
  BUF_X1 U2170 ( .A(n1342), .Z(n1341) );
  NAND2_X1 U2171 ( .A1(n1293), .A2(cw_dec[0]), .ZN(\unit_decode/n3522 ) );
  NAND2_X1 U2172 ( .A1(aluout_regn[1]), .A2(\unit_memory/DRAM/n552 ), .ZN(
        \unit_memory/DRAM/n583 ) );
  NOR2_X1 U2173 ( .A1(\unit_memory/DRAM/n550 ), .A2(aluout_regn[2]), .ZN(
        \unit_memory/DRAM/n758 ) );
  NOR2_X1 U2174 ( .A1(\unit_memory/DRAM/n551 ), .A2(aluout_regn[2]), .ZN(
        \unit_memory/DRAM/n755 ) );
  NOR2_X1 U2175 ( .A1(\unit_memory/DRAM/n583 ), .A2(aluout_regn[2]), .ZN(
        \unit_memory/DRAM/n760 ) );
  NOR2_X1 U2176 ( .A1(\unit_memory/DRAM/n570 ), .A2(aluout_regn[2]), .ZN(
        \unit_memory/DRAM/n762 ) );
  INV_X1 U2177 ( .A(cw_dec[2]), .ZN(\unit_decode/n2186 ) );
  NAND2_X1 U2178 ( .A1(aluout_regn[1]), .A2(aluout_regn[0]), .ZN(
        \unit_memory/DRAM/n570 ) );
  INV_X1 U2179 ( .A(aluout_regn[2]), .ZN(\unit_memory/DRAM/n547 ) );
  AOI221_X1 U2180 ( .B1(n136), .B2(\unit_decode/n2116 ), .C1(
        \unit_decode/n237 ), .C2(\unit_decode/n2186 ), .A(n1322), .ZN(
        \unit_decode/IMMreg/ffi_0/n5 ) );
  AOI221_X1 U2181 ( .B1(n134), .B2(\unit_decode/n2114 ), .C1(
        \unit_decode/n225 ), .C2(\unit_decode/n2186 ), .A(n1326), .ZN(
        \unit_decode/IMMreg/ffi_2/n5 ) );
  AOI221_X1 U2182 ( .B1(n131), .B2(\unit_decode/n2108 ), .C1(
        \unit_decode/n3621 ), .C2(\unit_decode/n2186 ), .A(n1327), .ZN(
        \unit_decode/IMMreg/ffi_8/n5 ) );
  AOI221_X1 U2183 ( .B1(n130), .B2(\unit_decode/n2107 ), .C1(
        \unit_decode/n3620 ), .C2(\unit_decode/n2186 ), .A(n1325), .ZN(
        \unit_decode/IMMreg/ffi_9/n5 ) );
  AOI221_X1 U2184 ( .B1(n136), .B2(\unit_decode/n2115 ), .C1(
        \unit_decode/n229 ), .C2(\unit_decode/n2186 ), .A(n1323), .ZN(
        \unit_decode/IMMreg/ffi_1/n5 ) );
  AOI221_X1 U2185 ( .B1(n133), .B2(\unit_decode/n2113 ), .C1(
        \unit_decode/n231 ), .C2(\unit_decode/n2186 ), .A(n1323), .ZN(
        \unit_decode/IMMreg/ffi_3/n5 ) );
  AOI221_X1 U2186 ( .B1(n132), .B2(\unit_decode/n2112 ), .C1(
        \unit_decode/n211 ), .C2(\unit_decode/n2186 ), .A(n1327), .ZN(
        \unit_decode/IMMreg/ffi_4/n5 ) );
  AOI221_X1 U2187 ( .B1(n131), .B2(\unit_decode/n2111 ), .C1(
        \unit_decode/n213 ), .C2(\unit_decode/n2186 ), .A(n1324), .ZN(
        \unit_decode/IMMreg/ffi_5/n5 ) );
  AOI221_X1 U2188 ( .B1(n133), .B2(\unit_decode/n2110 ), .C1(
        \unit_decode/n197 ), .C2(\unit_decode/n2186 ), .A(n1322), .ZN(
        \unit_decode/IMMreg/ffi_6/n5 ) );
  AOI221_X1 U2189 ( .B1(n132), .B2(\unit_decode/n2109 ), .C1(
        \unit_decode/n209 ), .C2(\unit_decode/n2186 ), .A(n1325), .ZN(
        \unit_decode/IMMreg/ffi_7/n5 ) );
  AOI221_X1 U2190 ( .B1(n135), .B2(\unit_decode/n2106 ), .C1(
        \unit_decode/n3619 ), .C2(\unit_decode/n2186 ), .A(n1325), .ZN(
        \unit_decode/IMMreg/ffi_10/n5 ) );
  AOI221_X1 U2191 ( .B1(n134), .B2(\unit_decode/n2105 ), .C1(
        \unit_decode/n3618 ), .C2(\unit_decode/n2186 ), .A(n1323), .ZN(
        \unit_decode/IMMreg/ffi_11/n5 ) );
  AOI221_X1 U2192 ( .B1(n137), .B2(\unit_decode/n2104 ), .C1(
        \unit_decode/n3617 ), .C2(\unit_decode/n2186 ), .A(n1326), .ZN(
        \unit_decode/IMMreg/ffi_12/n5 ) );
  AOI221_X1 U2193 ( .B1(n130), .B2(\unit_decode/n2103 ), .C1(
        \unit_decode/n3616 ), .C2(\unit_decode/n2186 ), .A(n1324), .ZN(
        \unit_decode/IMMreg/ffi_13/n5 ) );
  AOI221_X1 U2194 ( .B1(n137), .B2(\unit_decode/n2102 ), .C1(
        \unit_decode/n3615 ), .C2(\unit_decode/n2186 ), .A(n1326), .ZN(
        \unit_decode/IMMreg/ffi_14/n5 ) );
  AOI221_X1 U2195 ( .B1(n137), .B2(\unit_decode/n2101 ), .C1(
        \unit_decode/n3614 ), .C2(\unit_decode/n2186 ), .A(n1324), .ZN(
        \unit_decode/IMMreg/ffi_15/n5 ) );
  NOR2_X1 U2196 ( .A1(\unit_memory/DRAM/n552 ), .A2(aluout_regn[1]), .ZN(
        \unit_memory/DRAM/n1148 ) );
  NOR2_X1 U2197 ( .A1(aluout_regn[0]), .A2(aluout_regn[1]), .ZN(
        \unit_memory/DRAM/n1143 ) );
  OAI221_X1 U2198 ( .B1(\unit_decode/n2100 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3613 ), .C2(n1300), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_16/n5 ) );
  OAI221_X1 U2199 ( .B1(\unit_decode/n2099 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3612 ), .C2(n1300), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_17/n5 ) );
  OAI221_X1 U2200 ( .B1(\unit_decode/n2098 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3611 ), .C2(n1300), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_18/n5 ) );
  OAI221_X1 U2201 ( .B1(\unit_decode/n2097 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3610 ), .C2(n1300), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_19/n5 ) );
  OAI221_X1 U2202 ( .B1(\unit_decode/n2096 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3609 ), .C2(n1300), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_20/n5 ) );
  OAI221_X1 U2203 ( .B1(\unit_decode/n2095 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3608 ), .C2(n1299), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_21/n5 ) );
  OAI221_X1 U2204 ( .B1(\unit_decode/n2094 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3607 ), .C2(n1299), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_22/n5 ) );
  OAI221_X1 U2205 ( .B1(\unit_decode/n2093 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3606 ), .C2(n1299), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_23/n5 ) );
  OAI221_X1 U2206 ( .B1(\unit_decode/n2092 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3605 ), .C2(n1299), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_24/n5 ) );
  OAI221_X1 U2207 ( .B1(\unit_decode/n2091 ), .B2(\unit_decode/n3522 ), .C1(
        \unit_decode/n3604 ), .C2(n1299), .A(\unit_decode/n3520 ), .ZN(
        \unit_decode/IMMreg/ffi_25/n5 ) );
  NOR2_X1 U2208 ( .A1(\unit_memory/DRAM/n546 ), .A2(aluout_regn[4]), .ZN(
        \unit_memory/DRAM/n782 ) );
  NOR2_X1 U2209 ( .A1(aluout_regn[3]), .A2(aluout_regn[4]), .ZN(
        \unit_memory/DRAM/n772 ) );
  NAND4_X1 U2210 ( .A1(IR_OUT[27]), .A2(IR_OUT[26]), .A3(\unit_decode/n3517 ), 
        .A4(\unit_decode/n2090 ), .ZN(\unit_decode/n3516 ) );
  AND2_X1 U2211 ( .A1(\unit_decode/n3520 ), .A2(\unit_decode/n3521 ), .ZN(
        \unit_decode/n3519 ) );
  NAND4_X1 U2212 ( .A1(cw_dec[0]), .A2(n1293), .A3(IR_OUT[25]), .A4(
        \unit_decode/n2189 ), .ZN(\unit_decode/n3521 ) );
  OAI22_X1 U2213 ( .A1(n1285), .A2(\unit_decode/n1141 ), .B1(n1305), .B2(
        \unit_decode/n199 ), .ZN(\unit_decode/Areg/ffi_0/n5 ) );
  INV_X1 U2214 ( .A(\unit_decode/registerA[0] ), .ZN(\unit_decode/n1141 ) );
  OAI22_X1 U2215 ( .A1(n1286), .A2(\unit_decode/n1142 ), .B1(n1305), .B2(
        \unit_decode/n203 ), .ZN(\unit_decode/Areg/ffi_1/n5 ) );
  INV_X1 U2216 ( .A(\unit_decode/registerA[1] ), .ZN(\unit_decode/n1142 ) );
  OAI22_X1 U2217 ( .A1(n1285), .A2(\unit_decode/n1151 ), .B1(n1305), .B2(
        \unit_decode/n3531 ), .ZN(\unit_decode/Areg/ffi_10/n5 ) );
  INV_X1 U2218 ( .A(\unit_decode/registerA[10] ), .ZN(\unit_decode/n1151 ) );
  OAI22_X1 U2219 ( .A1(n1292), .A2(\unit_decode/n1152 ), .B1(n1305), .B2(
        \unit_decode/n3530 ), .ZN(\unit_decode/Areg/ffi_11/n5 ) );
  INV_X1 U2220 ( .A(\unit_decode/registerA[11] ), .ZN(\unit_decode/n1152 ) );
  OAI22_X1 U2221 ( .A1(n1291), .A2(\unit_decode/n1153 ), .B1(n1305), .B2(
        \unit_decode/n3529 ), .ZN(\unit_decode/Areg/ffi_12/n5 ) );
  INV_X1 U2222 ( .A(\unit_decode/registerA[12] ), .ZN(\unit_decode/n1153 ) );
  OR4_X1 U2223 ( .A1(\unit_decode/n2101 ), .A2(\unit_decode/n3512 ), .A3(
        cw_dec[0]), .A4(cw_dec[1]), .ZN(\unit_decode/n3520 ) );
  OAI22_X1 U2224 ( .A1(n950), .A2(n728), .B1(n949), .B2(\unit_decode/n1786 ), 
        .ZN(\unit_decode/RegisterFile/n1648 ) );
  OAI22_X1 U2225 ( .A1(n950), .A2(n731), .B1(n949), .B2(\unit_decode/n1787 ), 
        .ZN(\unit_decode/RegisterFile/n1647 ) );
  OAI22_X1 U2226 ( .A1(n951), .A2(n734), .B1(\unit_decode/n2254 ), .B2(
        \unit_decode/n1788 ), .ZN(\unit_decode/RegisterFile/n1646 ) );
  OAI22_X1 U2227 ( .A1(n951), .A2(n737), .B1(\unit_decode/n2254 ), .B2(
        \unit_decode/n1789 ), .ZN(\unit_decode/RegisterFile/n1645 ) );
  OAI22_X1 U2228 ( .A1(n951), .A2(n740), .B1(\unit_decode/n2254 ), .B2(
        \unit_decode/n1790 ), .ZN(\unit_decode/RegisterFile/n1644 ) );
  OAI22_X1 U2229 ( .A1(n951), .A2(n743), .B1(\unit_decode/n2254 ), .B2(
        \unit_decode/n2060 ), .ZN(\unit_decode/RegisterFile/n1643 ) );
  OAI22_X1 U2230 ( .A1(n923), .A2(n710), .B1(n922), .B2(\unit_decode/n1807 ), 
        .ZN(\unit_decode/RegisterFile/n1747 ) );
  OAI22_X1 U2231 ( .A1(n923), .A2(n722), .B1(n922), .B2(\unit_decode/n1808 ), 
        .ZN(\unit_decode/RegisterFile/n1746 ) );
  OAI22_X1 U2232 ( .A1(n923), .A2(n725), .B1(n922), .B2(\unit_decode/n1809 ), 
        .ZN(\unit_decode/RegisterFile/n1745 ) );
  OAI22_X1 U2233 ( .A1(n923), .A2(n728), .B1(n922), .B2(\unit_decode/n1810 ), 
        .ZN(\unit_decode/RegisterFile/n1744 ) );
  OAI22_X1 U2234 ( .A1(n923), .A2(n731), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1811 ), .ZN(\unit_decode/RegisterFile/n1743 ) );
  OAI22_X1 U2235 ( .A1(n924), .A2(n734), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1812 ), .ZN(\unit_decode/RegisterFile/n1742 ) );
  OAI22_X1 U2236 ( .A1(n924), .A2(n737), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1813 ), .ZN(\unit_decode/RegisterFile/n1741 ) );
  OAI22_X1 U2237 ( .A1(n924), .A2(n740), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1814 ), .ZN(\unit_decode/RegisterFile/n1740 ) );
  OAI22_X1 U2238 ( .A1(n914), .A2(n710), .B1(n913), .B2(\unit_decode/n1815 ), 
        .ZN(\unit_decode/RegisterFile/n1779 ) );
  OAI22_X1 U2239 ( .A1(n914), .A2(n722), .B1(n913), .B2(\unit_decode/n1816 ), 
        .ZN(\unit_decode/RegisterFile/n1778 ) );
  OAI22_X1 U2240 ( .A1(n914), .A2(n725), .B1(n913), .B2(\unit_decode/n1817 ), 
        .ZN(\unit_decode/RegisterFile/n1777 ) );
  OAI22_X1 U2241 ( .A1(n914), .A2(n728), .B1(n913), .B2(\unit_decode/n1818 ), 
        .ZN(\unit_decode/RegisterFile/n1776 ) );
  OAI22_X1 U2242 ( .A1(n914), .A2(n731), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1819 ), .ZN(\unit_decode/RegisterFile/n1775 ) );
  OAI22_X1 U2243 ( .A1(n915), .A2(n734), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1820 ), .ZN(\unit_decode/RegisterFile/n1774 ) );
  OAI22_X1 U2244 ( .A1(n915), .A2(n737), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1821 ), .ZN(\unit_decode/RegisterFile/n1773 ) );
  OAI22_X1 U2245 ( .A1(n915), .A2(n740), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1822 ), .ZN(\unit_decode/RegisterFile/n1772 ) );
  OAI22_X1 U2246 ( .A1(n887), .A2(n709), .B1(n886), .B2(\unit_decode/n1839 ), 
        .ZN(\unit_decode/RegisterFile/n1875 ) );
  OAI22_X1 U2247 ( .A1(n887), .A2(n721), .B1(n886), .B2(\unit_decode/n1840 ), 
        .ZN(\unit_decode/RegisterFile/n1874 ) );
  OAI22_X1 U2248 ( .A1(n887), .A2(n724), .B1(n886), .B2(\unit_decode/n1841 ), 
        .ZN(\unit_decode/RegisterFile/n1873 ) );
  OAI22_X1 U2249 ( .A1(n887), .A2(n727), .B1(n886), .B2(\unit_decode/n1842 ), 
        .ZN(\unit_decode/RegisterFile/n1872 ) );
  OAI22_X1 U2250 ( .A1(n887), .A2(n730), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1843 ), .ZN(\unit_decode/RegisterFile/n1871 ) );
  OAI22_X1 U2251 ( .A1(n888), .A2(n733), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1844 ), .ZN(\unit_decode/RegisterFile/n1870 ) );
  OAI22_X1 U2252 ( .A1(n888), .A2(n736), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1845 ), .ZN(\unit_decode/RegisterFile/n1869 ) );
  OAI22_X1 U2253 ( .A1(n888), .A2(n739), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1846 ), .ZN(\unit_decode/RegisterFile/n1868 ) );
  OAI22_X1 U2254 ( .A1(n878), .A2(n709), .B1(n877), .B2(\unit_decode/n1847 ), 
        .ZN(\unit_decode/RegisterFile/n1907 ) );
  OAI22_X1 U2255 ( .A1(n878), .A2(n721), .B1(n877), .B2(\unit_decode/n1848 ), 
        .ZN(\unit_decode/RegisterFile/n1906 ) );
  OAI22_X1 U2256 ( .A1(n878), .A2(n724), .B1(n877), .B2(\unit_decode/n1849 ), 
        .ZN(\unit_decode/RegisterFile/n1905 ) );
  OAI22_X1 U2257 ( .A1(n878), .A2(n727), .B1(n877), .B2(\unit_decode/n1850 ), 
        .ZN(\unit_decode/RegisterFile/n1904 ) );
  OAI22_X1 U2258 ( .A1(n878), .A2(n730), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1851 ), .ZN(\unit_decode/RegisterFile/n1903 ) );
  OAI22_X1 U2259 ( .A1(n879), .A2(n733), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1852 ), .ZN(\unit_decode/RegisterFile/n1902 ) );
  OAI22_X1 U2260 ( .A1(n879), .A2(n736), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1853 ), .ZN(\unit_decode/RegisterFile/n1901 ) );
  OAI22_X1 U2261 ( .A1(n879), .A2(n739), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1854 ), .ZN(\unit_decode/RegisterFile/n1900 ) );
  OAI22_X1 U2262 ( .A1(n1076), .A2(n711), .B1(n1075), .B2(\unit_decode/n1855 ), 
        .ZN(\unit_decode/RegisterFile/n1203 ) );
  OAI22_X1 U2263 ( .A1(n1076), .A2(n723), .B1(n1075), .B2(\unit_decode/n1856 ), 
        .ZN(\unit_decode/RegisterFile/n1202 ) );
  OAI22_X1 U2264 ( .A1(n1076), .A2(n726), .B1(n1075), .B2(\unit_decode/n1857 ), 
        .ZN(\unit_decode/RegisterFile/n1201 ) );
  OAI22_X1 U2265 ( .A1(n1076), .A2(n729), .B1(n1075), .B2(\unit_decode/n1858 ), 
        .ZN(\unit_decode/RegisterFile/n1200 ) );
  OAI22_X1 U2266 ( .A1(n1076), .A2(n732), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1859 ), .ZN(\unit_decode/RegisterFile/n1199 ) );
  OAI22_X1 U2267 ( .A1(n1077), .A2(n735), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1860 ), .ZN(\unit_decode/RegisterFile/n1198 ) );
  OAI22_X1 U2268 ( .A1(n1077), .A2(n738), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1861 ), .ZN(\unit_decode/RegisterFile/n1197 ) );
  OAI22_X1 U2269 ( .A1(n1077), .A2(n741), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1862 ), .ZN(\unit_decode/RegisterFile/n1196 ) );
  OAI22_X1 U2270 ( .A1(n851), .A2(n709), .B1(n850), .B2(\unit_decode/n1908 ), 
        .ZN(\unit_decode/RegisterFile/n2003 ) );
  OAI22_X1 U2271 ( .A1(n851), .A2(n721), .B1(n850), .B2(\unit_decode/n1909 ), 
        .ZN(\unit_decode/RegisterFile/n2002 ) );
  OAI22_X1 U2272 ( .A1(n851), .A2(n724), .B1(n850), .B2(\unit_decode/n1910 ), 
        .ZN(\unit_decode/RegisterFile/n2001 ) );
  OAI22_X1 U2273 ( .A1(n851), .A2(n727), .B1(n850), .B2(\unit_decode/n1911 ), 
        .ZN(\unit_decode/RegisterFile/n2000 ) );
  OAI22_X1 U2274 ( .A1(n851), .A2(n730), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1912 ), .ZN(\unit_decode/RegisterFile/n1999 ) );
  OAI22_X1 U2275 ( .A1(n852), .A2(n733), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1913 ), .ZN(\unit_decode/RegisterFile/n1998 ) );
  OAI22_X1 U2276 ( .A1(n852), .A2(n736), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1914 ), .ZN(\unit_decode/RegisterFile/n1997 ) );
  OAI22_X1 U2277 ( .A1(n852), .A2(n739), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1915 ), .ZN(\unit_decode/RegisterFile/n1996 ) );
  OAI22_X1 U2278 ( .A1(n842), .A2(n709), .B1(n841), .B2(\unit_decode/n1916 ), 
        .ZN(\unit_decode/RegisterFile/n2035 ) );
  OAI22_X1 U2279 ( .A1(n842), .A2(n721), .B1(n841), .B2(\unit_decode/n1917 ), 
        .ZN(\unit_decode/RegisterFile/n2034 ) );
  OAI22_X1 U2280 ( .A1(n842), .A2(n724), .B1(n841), .B2(\unit_decode/n1918 ), 
        .ZN(\unit_decode/RegisterFile/n2033 ) );
  OAI22_X1 U2281 ( .A1(n842), .A2(n727), .B1(n841), .B2(\unit_decode/n1919 ), 
        .ZN(\unit_decode/RegisterFile/n2032 ) );
  OAI22_X1 U2282 ( .A1(n842), .A2(n730), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1920 ), .ZN(\unit_decode/RegisterFile/n2031 ) );
  OAI22_X1 U2283 ( .A1(n843), .A2(n733), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1921 ), .ZN(\unit_decode/RegisterFile/n2030 ) );
  OAI22_X1 U2284 ( .A1(n843), .A2(n736), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1922 ), .ZN(\unit_decode/RegisterFile/n2029 ) );
  OAI22_X1 U2285 ( .A1(n843), .A2(n739), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1923 ), .ZN(\unit_decode/RegisterFile/n2028 ) );
  OAI22_X1 U2286 ( .A1(n815), .A2(n709), .B1(n814), .B2(\unit_decode/n1940 ), 
        .ZN(\unit_decode/RegisterFile/n2131 ) );
  OAI22_X1 U2287 ( .A1(n815), .A2(n721), .B1(n814), .B2(\unit_decode/n1941 ), 
        .ZN(\unit_decode/RegisterFile/n2130 ) );
  OAI22_X1 U2288 ( .A1(n815), .A2(n724), .B1(n814), .B2(\unit_decode/n1942 ), 
        .ZN(\unit_decode/RegisterFile/n2129 ) );
  OAI22_X1 U2289 ( .A1(n815), .A2(n727), .B1(n814), .B2(\unit_decode/n1943 ), 
        .ZN(\unit_decode/RegisterFile/n2128 ) );
  OAI22_X1 U2290 ( .A1(n815), .A2(n730), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1944 ), .ZN(\unit_decode/RegisterFile/n2127 ) );
  OAI22_X1 U2291 ( .A1(n816), .A2(n733), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1945 ), .ZN(\unit_decode/RegisterFile/n2126 ) );
  OAI22_X1 U2292 ( .A1(n816), .A2(n736), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1946 ), .ZN(\unit_decode/RegisterFile/n2125 ) );
  OAI22_X1 U2293 ( .A1(n816), .A2(n739), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1947 ), .ZN(\unit_decode/RegisterFile/n2124 ) );
  OAI22_X1 U2294 ( .A1(n713), .A2(n709), .B1(n712), .B2(\unit_decode/n1948 ), 
        .ZN(\unit_decode/RegisterFile/n2163 ) );
  OAI22_X1 U2295 ( .A1(n713), .A2(n721), .B1(n712), .B2(\unit_decode/n1949 ), 
        .ZN(\unit_decode/RegisterFile/n2162 ) );
  OAI22_X1 U2296 ( .A1(n713), .A2(n724), .B1(n712), .B2(\unit_decode/n1950 ), 
        .ZN(\unit_decode/RegisterFile/n2161 ) );
  OAI22_X1 U2297 ( .A1(n713), .A2(n727), .B1(n712), .B2(\unit_decode/n1951 ), 
        .ZN(\unit_decode/RegisterFile/n2160 ) );
  OAI22_X1 U2298 ( .A1(n713), .A2(n730), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1952 ), .ZN(\unit_decode/RegisterFile/n2159 ) );
  OAI22_X1 U2299 ( .A1(n714), .A2(n733), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1953 ), .ZN(\unit_decode/RegisterFile/n2158 ) );
  OAI22_X1 U2300 ( .A1(n714), .A2(n736), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1954 ), .ZN(\unit_decode/RegisterFile/n2157 ) );
  OAI22_X1 U2301 ( .A1(n714), .A2(n739), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1955 ), .ZN(\unit_decode/RegisterFile/n2156 ) );
  OAI22_X1 U2302 ( .A1(n1087), .A2(\unit_decode/n1189 ), .B1(n1085), .B2(n741), 
        .ZN(\unit_decode/RegisterFile/n1164 ) );
  OAI22_X1 U2303 ( .A1(n1087), .A2(\unit_decode/n1190 ), .B1(n1084), .B2(n738), 
        .ZN(\unit_decode/RegisterFile/n1165 ) );
  OAI22_X1 U2304 ( .A1(n1087), .A2(\unit_decode/n1191 ), .B1(n1085), .B2(n735), 
        .ZN(\unit_decode/RegisterFile/n1166 ) );
  OAI22_X1 U2305 ( .A1(n1086), .A2(\unit_decode/n1192 ), .B1(n1084), .B2(n732), 
        .ZN(\unit_decode/RegisterFile/n1167 ) );
  OAI22_X1 U2306 ( .A1(n1086), .A2(\unit_decode/n1193 ), .B1(n1085), .B2(n729), 
        .ZN(\unit_decode/RegisterFile/n1168 ) );
  OAI22_X1 U2307 ( .A1(n1086), .A2(\unit_decode/n1194 ), .B1(n1084), .B2(n726), 
        .ZN(\unit_decode/RegisterFile/n1169 ) );
  OAI22_X1 U2308 ( .A1(n1086), .A2(\unit_decode/n1195 ), .B1(n1085), .B2(n723), 
        .ZN(\unit_decode/RegisterFile/n1170 ) );
  OAI22_X1 U2309 ( .A1(n1086), .A2(\unit_decode/n1196 ), .B1(n1084), .B2(n711), 
        .ZN(\unit_decode/RegisterFile/n1171 ) );
  OAI22_X1 U2310 ( .A1(n1037), .A2(n813), .B1(\unit_decode/n2265 ), .B2(
        \unit_decode/n1317 ), .ZN(\unit_decode/RegisterFile/n1332 ) );
  OAI22_X1 U2311 ( .A1(n1037), .A2(n810), .B1(n1030), .B2(\unit_decode/n1318 ), 
        .ZN(\unit_decode/RegisterFile/n1333 ) );
  OAI22_X1 U2312 ( .A1(n1036), .A2(n807), .B1(\unit_decode/n2265 ), .B2(
        \unit_decode/n1319 ), .ZN(\unit_decode/RegisterFile/n1334 ) );
  OAI22_X1 U2313 ( .A1(n1036), .A2(n804), .B1(n1030), .B2(\unit_decode/n1320 ), 
        .ZN(\unit_decode/RegisterFile/n1335 ) );
  OAI22_X1 U2314 ( .A1(n1036), .A2(n801), .B1(\unit_decode/n2265 ), .B2(
        \unit_decode/n1321 ), .ZN(\unit_decode/RegisterFile/n1336 ) );
  OAI22_X1 U2315 ( .A1(n1036), .A2(n798), .B1(\unit_decode/n2265 ), .B2(
        \unit_decode/n1322 ), .ZN(\unit_decode/RegisterFile/n1337 ) );
  OAI22_X1 U2316 ( .A1(n1036), .A2(n795), .B1(\unit_decode/n2265 ), .B2(
        \unit_decode/n1323 ), .ZN(\unit_decode/RegisterFile/n1338 ) );
  OAI22_X1 U2317 ( .A1(n1028), .A2(n813), .B1(\unit_decode/n2263 ), .B2(
        \unit_decode/n1341 ), .ZN(\unit_decode/RegisterFile/n1364 ) );
  OAI22_X1 U2318 ( .A1(n1028), .A2(n810), .B1(n1021), .B2(\unit_decode/n1342 ), 
        .ZN(\unit_decode/RegisterFile/n1365 ) );
  OAI22_X1 U2319 ( .A1(n1027), .A2(n807), .B1(\unit_decode/n2263 ), .B2(
        \unit_decode/n1343 ), .ZN(\unit_decode/RegisterFile/n1366 ) );
  OAI22_X1 U2320 ( .A1(n1027), .A2(n804), .B1(n1021), .B2(\unit_decode/n1344 ), 
        .ZN(\unit_decode/RegisterFile/n1367 ) );
  OAI22_X1 U2321 ( .A1(n1027), .A2(n801), .B1(\unit_decode/n2263 ), .B2(
        \unit_decode/n1345 ), .ZN(\unit_decode/RegisterFile/n1368 ) );
  OAI22_X1 U2322 ( .A1(n1027), .A2(n798), .B1(\unit_decode/n2263 ), .B2(
        \unit_decode/n1346 ), .ZN(\unit_decode/RegisterFile/n1369 ) );
  OAI22_X1 U2323 ( .A1(n1027), .A2(n795), .B1(\unit_decode/n2263 ), .B2(
        \unit_decode/n1347 ), .ZN(\unit_decode/RegisterFile/n1370 ) );
  OAI22_X1 U2324 ( .A1(n964), .A2(n794), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n2053 ), .ZN(\unit_decode/RegisterFile/n1594 ) );
  OAI22_X1 U2325 ( .A1(n964), .A2(n797), .B1(n958), .B2(\unit_decode/n2054 ), 
        .ZN(\unit_decode/RegisterFile/n1593 ) );
  OAI22_X1 U2326 ( .A1(n964), .A2(n800), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n2055 ), .ZN(\unit_decode/RegisterFile/n1592 ) );
  OAI22_X1 U2327 ( .A1(n964), .A2(n803), .B1(n958), .B2(\unit_decode/n2056 ), 
        .ZN(\unit_decode/RegisterFile/n1591 ) );
  OAI22_X1 U2328 ( .A1(n964), .A2(n806), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n2057 ), .ZN(\unit_decode/RegisterFile/n1590 ) );
  OAI22_X1 U2329 ( .A1(n965), .A2(n809), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n2058 ), .ZN(\unit_decode/RegisterFile/n1589 ) );
  OAI22_X1 U2330 ( .A1(n965), .A2(n812), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n2059 ), .ZN(\unit_decode/RegisterFile/n1588 ) );
  OAI22_X1 U2331 ( .A1(n358), .A2(n694), .B1(\unit_memory/DRAM/n3390 ), .B2(
        n692), .ZN(\unit_memory/DRAM/n1157 ) );
  OAI22_X1 U2332 ( .A1(n1035), .A2(n792), .B1(n1030), .B2(\unit_decode/n1324 ), 
        .ZN(\unit_decode/RegisterFile/n1339 ) );
  OAI22_X1 U2333 ( .A1(n1035), .A2(n789), .B1(n1030), .B2(\unit_decode/n1325 ), 
        .ZN(\unit_decode/RegisterFile/n1340 ) );
  OAI22_X1 U2334 ( .A1(n1035), .A2(n786), .B1(n1030), .B2(\unit_decode/n1326 ), 
        .ZN(\unit_decode/RegisterFile/n1341 ) );
  OAI22_X1 U2335 ( .A1(n1035), .A2(n783), .B1(n1030), .B2(\unit_decode/n1327 ), 
        .ZN(\unit_decode/RegisterFile/n1342 ) );
  OAI22_X1 U2336 ( .A1(n1035), .A2(n780), .B1(n1030), .B2(\unit_decode/n1328 ), 
        .ZN(\unit_decode/RegisterFile/n1343 ) );
  OAI22_X1 U2337 ( .A1(n1034), .A2(n777), .B1(n1030), .B2(\unit_decode/n1329 ), 
        .ZN(\unit_decode/RegisterFile/n1344 ) );
  OAI22_X1 U2338 ( .A1(n1034), .A2(n774), .B1(n1030), .B2(\unit_decode/n1330 ), 
        .ZN(\unit_decode/RegisterFile/n1345 ) );
  OAI22_X1 U2339 ( .A1(n1034), .A2(n771), .B1(n1030), .B2(\unit_decode/n1331 ), 
        .ZN(\unit_decode/RegisterFile/n1346 ) );
  OAI22_X1 U2340 ( .A1(n1034), .A2(n768), .B1(n1030), .B2(\unit_decode/n1332 ), 
        .ZN(\unit_decode/RegisterFile/n1347 ) );
  OAI22_X1 U2341 ( .A1(n1034), .A2(n765), .B1(n1030), .B2(\unit_decode/n1333 ), 
        .ZN(\unit_decode/RegisterFile/n1348 ) );
  OAI22_X1 U2342 ( .A1(n1033), .A2(n762), .B1(n1030), .B2(\unit_decode/n1334 ), 
        .ZN(\unit_decode/RegisterFile/n1349 ) );
  OAI22_X1 U2343 ( .A1(n1033), .A2(n759), .B1(n1030), .B2(\unit_decode/n1335 ), 
        .ZN(\unit_decode/RegisterFile/n1350 ) );
  OAI22_X1 U2344 ( .A1(n1033), .A2(n756), .B1(n1030), .B2(\unit_decode/n1336 ), 
        .ZN(\unit_decode/RegisterFile/n1351 ) );
  OAI22_X1 U2345 ( .A1(n1026), .A2(n792), .B1(n1021), .B2(\unit_decode/n1348 ), 
        .ZN(\unit_decode/RegisterFile/n1371 ) );
  OAI22_X1 U2346 ( .A1(n1026), .A2(n789), .B1(n1021), .B2(\unit_decode/n1349 ), 
        .ZN(\unit_decode/RegisterFile/n1372 ) );
  OAI22_X1 U2347 ( .A1(n1026), .A2(n786), .B1(n1021), .B2(\unit_decode/n1350 ), 
        .ZN(\unit_decode/RegisterFile/n1373 ) );
  OAI22_X1 U2348 ( .A1(n1026), .A2(n783), .B1(n1021), .B2(\unit_decode/n1351 ), 
        .ZN(\unit_decode/RegisterFile/n1374 ) );
  OAI22_X1 U2349 ( .A1(n1026), .A2(n780), .B1(n1021), .B2(\unit_decode/n1352 ), 
        .ZN(\unit_decode/RegisterFile/n1375 ) );
  OAI22_X1 U2350 ( .A1(n1025), .A2(n777), .B1(n1021), .B2(\unit_decode/n1353 ), 
        .ZN(\unit_decode/RegisterFile/n1376 ) );
  OAI22_X1 U2351 ( .A1(n1025), .A2(n774), .B1(n1021), .B2(\unit_decode/n1354 ), 
        .ZN(\unit_decode/RegisterFile/n1377 ) );
  OAI22_X1 U2352 ( .A1(n1025), .A2(n771), .B1(n1021), .B2(\unit_decode/n1355 ), 
        .ZN(\unit_decode/RegisterFile/n1378 ) );
  OAI22_X1 U2353 ( .A1(n1025), .A2(n768), .B1(n1021), .B2(\unit_decode/n1356 ), 
        .ZN(\unit_decode/RegisterFile/n1379 ) );
  OAI22_X1 U2354 ( .A1(n1025), .A2(n765), .B1(n1021), .B2(\unit_decode/n1357 ), 
        .ZN(\unit_decode/RegisterFile/n1380 ) );
  OAI22_X1 U2355 ( .A1(n1024), .A2(n762), .B1(n1021), .B2(\unit_decode/n1358 ), 
        .ZN(\unit_decode/RegisterFile/n1381 ) );
  OAI22_X1 U2356 ( .A1(n1024), .A2(n759), .B1(n1021), .B2(\unit_decode/n1359 ), 
        .ZN(\unit_decode/RegisterFile/n1382 ) );
  OAI22_X1 U2357 ( .A1(n1024), .A2(n756), .B1(n1021), .B2(\unit_decode/n1360 ), 
        .ZN(\unit_decode/RegisterFile/n1383 ) );
  OAI22_X1 U2358 ( .A1(n961), .A2(n755), .B1(n958), .B2(\unit_decode/n2040 ), 
        .ZN(\unit_decode/RegisterFile/n1607 ) );
  OAI22_X1 U2359 ( .A1(n961), .A2(n758), .B1(n958), .B2(\unit_decode/n2041 ), 
        .ZN(\unit_decode/RegisterFile/n1606 ) );
  OAI22_X1 U2360 ( .A1(n961), .A2(n761), .B1(n958), .B2(\unit_decode/n2042 ), 
        .ZN(\unit_decode/RegisterFile/n1605 ) );
  OAI22_X1 U2361 ( .A1(n962), .A2(n764), .B1(n958), .B2(\unit_decode/n2043 ), 
        .ZN(\unit_decode/RegisterFile/n1604 ) );
  OAI22_X1 U2362 ( .A1(n962), .A2(n767), .B1(n958), .B2(\unit_decode/n2044 ), 
        .ZN(\unit_decode/RegisterFile/n1603 ) );
  OAI22_X1 U2363 ( .A1(n962), .A2(n770), .B1(n958), .B2(\unit_decode/n2045 ), 
        .ZN(\unit_decode/RegisterFile/n1602 ) );
  OAI22_X1 U2364 ( .A1(n962), .A2(n773), .B1(n958), .B2(\unit_decode/n2046 ), 
        .ZN(\unit_decode/RegisterFile/n1601 ) );
  OAI22_X1 U2365 ( .A1(n962), .A2(n776), .B1(n958), .B2(\unit_decode/n2047 ), 
        .ZN(\unit_decode/RegisterFile/n1600 ) );
  OAI22_X1 U2366 ( .A1(n963), .A2(n779), .B1(n958), .B2(\unit_decode/n2048 ), 
        .ZN(\unit_decode/RegisterFile/n1599 ) );
  OAI22_X1 U2367 ( .A1(n963), .A2(n782), .B1(n958), .B2(\unit_decode/n2049 ), 
        .ZN(\unit_decode/RegisterFile/n1598 ) );
  OAI22_X1 U2368 ( .A1(n963), .A2(n785), .B1(n958), .B2(\unit_decode/n2050 ), 
        .ZN(\unit_decode/RegisterFile/n1597 ) );
  OAI22_X1 U2369 ( .A1(n963), .A2(n788), .B1(n958), .B2(\unit_decode/n2051 ), 
        .ZN(\unit_decode/RegisterFile/n1596 ) );
  OAI22_X1 U2370 ( .A1(n963), .A2(n791), .B1(n958), .B2(\unit_decode/n2052 ), 
        .ZN(\unit_decode/RegisterFile/n1595 ) );
  OAI22_X1 U2371 ( .A1(n1013), .A2(n710), .B1(\unit_decode/RegisterFile/n3708 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1427 ) );
  OAI22_X1 U2372 ( .A1(n1013), .A2(n722), .B1(\unit_decode/RegisterFile/n3709 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1426 ) );
  OAI22_X1 U2373 ( .A1(n1013), .A2(n725), .B1(\unit_decode/RegisterFile/n3710 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1425 ) );
  OAI22_X1 U2374 ( .A1(n1013), .A2(n728), .B1(\unit_decode/RegisterFile/n3711 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1424 ) );
  OAI22_X1 U2375 ( .A1(n1013), .A2(n731), .B1(\unit_decode/RegisterFile/n3712 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1423 ) );
  OAI22_X1 U2376 ( .A1(n1014), .A2(n734), .B1(\unit_decode/RegisterFile/n3713 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1422 ) );
  OAI22_X1 U2377 ( .A1(n1014), .A2(n737), .B1(\unit_decode/RegisterFile/n3714 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1421 ) );
  OAI22_X1 U2378 ( .A1(n1014), .A2(n740), .B1(\unit_decode/RegisterFile/n3715 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1420 ) );
  OAI22_X1 U2379 ( .A1(n1004), .A2(n710), .B1(\unit_decode/RegisterFile/n3676 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1459 ) );
  OAI22_X1 U2380 ( .A1(n1004), .A2(n722), .B1(\unit_decode/RegisterFile/n3677 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1458 ) );
  OAI22_X1 U2381 ( .A1(n1004), .A2(n725), .B1(\unit_decode/RegisterFile/n3678 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1457 ) );
  OAI22_X1 U2382 ( .A1(n1004), .A2(n728), .B1(\unit_decode/RegisterFile/n3679 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1456 ) );
  OAI22_X1 U2383 ( .A1(n1004), .A2(n731), .B1(\unit_decode/RegisterFile/n3680 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1455 ) );
  OAI22_X1 U2384 ( .A1(n1005), .A2(n734), .B1(\unit_decode/RegisterFile/n3681 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1454 ) );
  OAI22_X1 U2385 ( .A1(n1005), .A2(n737), .B1(\unit_decode/RegisterFile/n3682 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1453 ) );
  OAI22_X1 U2386 ( .A1(n1005), .A2(n740), .B1(\unit_decode/RegisterFile/n3683 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1452 ) );
  OAI22_X1 U2387 ( .A1(n995), .A2(n710), .B1(\unit_decode/RegisterFile/n3644 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1491 ) );
  OAI22_X1 U2388 ( .A1(n995), .A2(n722), .B1(\unit_decode/RegisterFile/n3645 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1490 ) );
  OAI22_X1 U2389 ( .A1(n995), .A2(n725), .B1(\unit_decode/RegisterFile/n3646 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1489 ) );
  OAI22_X1 U2390 ( .A1(n995), .A2(n728), .B1(\unit_decode/RegisterFile/n3647 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1488 ) );
  OAI22_X1 U2391 ( .A1(n995), .A2(n731), .B1(\unit_decode/RegisterFile/n3648 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1487 ) );
  OAI22_X1 U2392 ( .A1(n996), .A2(n734), .B1(\unit_decode/RegisterFile/n3649 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1486 ) );
  OAI22_X1 U2393 ( .A1(n996), .A2(n737), .B1(\unit_decode/RegisterFile/n3650 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1485 ) );
  OAI22_X1 U2394 ( .A1(n996), .A2(n740), .B1(\unit_decode/RegisterFile/n3651 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1484 ) );
  OAI22_X1 U2395 ( .A1(n986), .A2(n710), .B1(\unit_decode/RegisterFile/n3612 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1523 ) );
  OAI22_X1 U2396 ( .A1(n986), .A2(n722), .B1(\unit_decode/RegisterFile/n3613 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1522 ) );
  OAI22_X1 U2397 ( .A1(n986), .A2(n725), .B1(\unit_decode/RegisterFile/n3614 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1521 ) );
  OAI22_X1 U2398 ( .A1(n986), .A2(n728), .B1(\unit_decode/RegisterFile/n3615 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1520 ) );
  OAI22_X1 U2399 ( .A1(n986), .A2(n731), .B1(\unit_decode/RegisterFile/n3616 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1519 ) );
  OAI22_X1 U2400 ( .A1(n987), .A2(n734), .B1(\unit_decode/RegisterFile/n3617 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1518 ) );
  OAI22_X1 U2401 ( .A1(n987), .A2(n737), .B1(\unit_decode/RegisterFile/n3618 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1517 ) );
  OAI22_X1 U2402 ( .A1(n987), .A2(n740), .B1(\unit_decode/RegisterFile/n3619 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1516 ) );
  OAI22_X1 U2403 ( .A1(n251), .A2(n257), .B1(\unit_memory/DRAM/n2367 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2180 ) );
  OAI22_X1 U2404 ( .A1(n257), .A2(n266), .B1(\unit_memory/DRAM/n2368 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2179 ) );
  OAI22_X1 U2405 ( .A1(n257), .A2(n269), .B1(\unit_memory/DRAM/n2369 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2178 ) );
  OAI22_X1 U2406 ( .A1(n257), .A2(n272), .B1(\unit_memory/DRAM/n2370 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2177 ) );
  OAI22_X1 U2407 ( .A1(n258), .A2(n275), .B1(\unit_memory/DRAM/n2371 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2176 ) );
  OAI22_X1 U2408 ( .A1(n258), .A2(n278), .B1(\unit_memory/DRAM/n2372 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2175 ) );
  OAI22_X1 U2409 ( .A1(n258), .A2(n281), .B1(\unit_memory/DRAM/n2373 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2174 ) );
  OAI22_X1 U2410 ( .A1(n258), .A2(n284), .B1(\unit_memory/DRAM/n2374 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2173 ) );
  OAI22_X1 U2411 ( .A1(n977), .A2(n728), .B1(\unit_decode/RegisterFile/n3583 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1552 ) );
  OAI22_X1 U2412 ( .A1(n977), .A2(n731), .B1(\unit_decode/RegisterFile/n3584 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1551 ) );
  OAI22_X1 U2413 ( .A1(n978), .A2(n734), .B1(\unit_decode/RegisterFile/n3585 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1550 ) );
  OAI22_X1 U2414 ( .A1(n978), .A2(n737), .B1(\unit_decode/RegisterFile/n3586 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1549 ) );
  OAI22_X1 U2415 ( .A1(n978), .A2(n740), .B1(\unit_decode/RegisterFile/n3587 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1548 ) );
  OAI22_X1 U2416 ( .A1(n955), .A2(n803), .B1(\unit_decode/RegisterFile/n3512 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1623 ) );
  OAI22_X1 U2417 ( .A1(n955), .A2(n806), .B1(\unit_decode/RegisterFile/n3513 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1622 ) );
  OAI22_X1 U2418 ( .A1(n1033), .A2(n753), .B1(n1030), .B2(\unit_decode/n1337 ), 
        .ZN(\unit_decode/RegisterFile/n1352 ) );
  OAI22_X1 U2419 ( .A1(n1033), .A2(n750), .B1(n1030), .B2(\unit_decode/n1338 ), 
        .ZN(\unit_decode/RegisterFile/n1353 ) );
  OAI22_X1 U2420 ( .A1(n1032), .A2(n747), .B1(n1030), .B2(\unit_decode/n1339 ), 
        .ZN(\unit_decode/RegisterFile/n1354 ) );
  OAI22_X1 U2421 ( .A1(n1032), .A2(n744), .B1(n1030), .B2(\unit_decode/n1340 ), 
        .ZN(\unit_decode/RegisterFile/n1355 ) );
  OAI22_X1 U2422 ( .A1(n1024), .A2(n753), .B1(n1021), .B2(\unit_decode/n1361 ), 
        .ZN(\unit_decode/RegisterFile/n1384 ) );
  OAI22_X1 U2423 ( .A1(n1024), .A2(n750), .B1(n1021), .B2(\unit_decode/n1362 ), 
        .ZN(\unit_decode/RegisterFile/n1385 ) );
  OAI22_X1 U2424 ( .A1(n1023), .A2(n747), .B1(n1021), .B2(\unit_decode/n1363 ), 
        .ZN(\unit_decode/RegisterFile/n1386 ) );
  OAI22_X1 U2425 ( .A1(n1023), .A2(n744), .B1(n1021), .B2(\unit_decode/n1364 ), 
        .ZN(\unit_decode/RegisterFile/n1387 ) );
  OAI22_X1 U2426 ( .A1(n959), .A2(n728), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n1778 ), .ZN(\unit_decode/RegisterFile/n1616 ) );
  OAI22_X1 U2427 ( .A1(n959), .A2(n731), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n1779 ), .ZN(\unit_decode/RegisterFile/n1615 ) );
  OAI22_X1 U2428 ( .A1(n960), .A2(n734), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n1780 ), .ZN(\unit_decode/RegisterFile/n1614 ) );
  OAI22_X1 U2429 ( .A1(n960), .A2(n737), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n1781 ), .ZN(\unit_decode/RegisterFile/n1613 ) );
  OAI22_X1 U2430 ( .A1(n960), .A2(n740), .B1(\unit_decode/n2256 ), .B2(
        \unit_decode/n1782 ), .ZN(\unit_decode/RegisterFile/n1612 ) );
  OAI22_X1 U2431 ( .A1(n960), .A2(n743), .B1(n958), .B2(\unit_decode/n2036 ), 
        .ZN(\unit_decode/RegisterFile/n1611 ) );
  OAI22_X1 U2432 ( .A1(n960), .A2(n746), .B1(n958), .B2(\unit_decode/n2037 ), 
        .ZN(\unit_decode/RegisterFile/n1610 ) );
  OAI22_X1 U2433 ( .A1(n961), .A2(n749), .B1(n958), .B2(\unit_decode/n2038 ), 
        .ZN(\unit_decode/RegisterFile/n1609 ) );
  OAI22_X1 U2434 ( .A1(n961), .A2(n752), .B1(n958), .B2(\unit_decode/n2039 ), 
        .ZN(\unit_decode/RegisterFile/n1608 ) );
  OAI22_X1 U2435 ( .A1(n1082), .A2(n813), .B1(n1075), .B2(\unit_decode/n1197 ), 
        .ZN(\unit_decode/RegisterFile/n1172 ) );
  OAI22_X1 U2436 ( .A1(n1082), .A2(n810), .B1(n1075), .B2(\unit_decode/n1198 ), 
        .ZN(\unit_decode/RegisterFile/n1173 ) );
  OAI22_X1 U2437 ( .A1(n1081), .A2(n807), .B1(n1075), .B2(\unit_decode/n1199 ), 
        .ZN(\unit_decode/RegisterFile/n1174 ) );
  OAI22_X1 U2438 ( .A1(n1081), .A2(n804), .B1(n1075), .B2(\unit_decode/n1200 ), 
        .ZN(\unit_decode/RegisterFile/n1175 ) );
  OAI22_X1 U2439 ( .A1(n1081), .A2(n801), .B1(n1075), .B2(\unit_decode/n1201 ), 
        .ZN(\unit_decode/RegisterFile/n1176 ) );
  OAI22_X1 U2440 ( .A1(n1081), .A2(n798), .B1(n1075), .B2(\unit_decode/n1202 ), 
        .ZN(\unit_decode/RegisterFile/n1177 ) );
  OAI22_X1 U2441 ( .A1(n1081), .A2(n795), .B1(n1075), .B2(\unit_decode/n1203 ), 
        .ZN(\unit_decode/RegisterFile/n1178 ) );
  OAI22_X1 U2442 ( .A1(n1080), .A2(n792), .B1(n1075), .B2(\unit_decode/n1204 ), 
        .ZN(\unit_decode/RegisterFile/n1179 ) );
  OAI22_X1 U2443 ( .A1(n1080), .A2(n789), .B1(n1075), .B2(\unit_decode/n1205 ), 
        .ZN(\unit_decode/RegisterFile/n1180 ) );
  OAI22_X1 U2444 ( .A1(n1080), .A2(n786), .B1(n1075), .B2(\unit_decode/n1206 ), 
        .ZN(\unit_decode/RegisterFile/n1181 ) );
  OAI22_X1 U2445 ( .A1(n1080), .A2(n783), .B1(n1075), .B2(\unit_decode/n1207 ), 
        .ZN(\unit_decode/RegisterFile/n1182 ) );
  OAI22_X1 U2446 ( .A1(n1080), .A2(n780), .B1(n1075), .B2(\unit_decode/n1208 ), 
        .ZN(\unit_decode/RegisterFile/n1183 ) );
  OAI22_X1 U2447 ( .A1(n1079), .A2(n777), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1209 ), .ZN(\unit_decode/RegisterFile/n1184 ) );
  OAI22_X1 U2448 ( .A1(n1079), .A2(n774), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1210 ), .ZN(\unit_decode/RegisterFile/n1185 ) );
  OAI22_X1 U2449 ( .A1(n1079), .A2(n771), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1211 ), .ZN(\unit_decode/RegisterFile/n1186 ) );
  OAI22_X1 U2450 ( .A1(n1079), .A2(n768), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1212 ), .ZN(\unit_decode/RegisterFile/n1187 ) );
  OAI22_X1 U2451 ( .A1(n1079), .A2(n765), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1213 ), .ZN(\unit_decode/RegisterFile/n1188 ) );
  OAI22_X1 U2452 ( .A1(n1078), .A2(n762), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1214 ), .ZN(\unit_decode/RegisterFile/n1189 ) );
  OAI22_X1 U2453 ( .A1(n1078), .A2(n759), .B1(\unit_decode/n2270 ), .B2(
        \unit_decode/n1215 ), .ZN(\unit_decode/RegisterFile/n1190 ) );
  OAI22_X1 U2454 ( .A1(n1078), .A2(n756), .B1(n1075), .B2(\unit_decode/n1216 ), 
        .ZN(\unit_decode/RegisterFile/n1191 ) );
  OAI22_X1 U2455 ( .A1(n1078), .A2(n753), .B1(n1075), .B2(\unit_decode/n1217 ), 
        .ZN(\unit_decode/RegisterFile/n1192 ) );
  OAI22_X1 U2456 ( .A1(n1078), .A2(n750), .B1(n1075), .B2(\unit_decode/n1218 ), 
        .ZN(\unit_decode/RegisterFile/n1193 ) );
  OAI22_X1 U2457 ( .A1(n1077), .A2(n747), .B1(n1075), .B2(\unit_decode/n1219 ), 
        .ZN(\unit_decode/RegisterFile/n1194 ) );
  OAI22_X1 U2458 ( .A1(n1077), .A2(n744), .B1(n1075), .B2(\unit_decode/n1220 ), 
        .ZN(\unit_decode/RegisterFile/n1195 ) );
  OAI22_X1 U2459 ( .A1(n929), .A2(n812), .B1(n922), .B2(\unit_decode/n1412 ), 
        .ZN(\unit_decode/RegisterFile/n1716 ) );
  OAI22_X1 U2460 ( .A1(n929), .A2(n809), .B1(n922), .B2(\unit_decode/n1413 ), 
        .ZN(\unit_decode/RegisterFile/n1717 ) );
  OAI22_X1 U2461 ( .A1(n928), .A2(n806), .B1(n922), .B2(\unit_decode/n1414 ), 
        .ZN(\unit_decode/RegisterFile/n1718 ) );
  OAI22_X1 U2462 ( .A1(n928), .A2(n803), .B1(n922), .B2(\unit_decode/n1415 ), 
        .ZN(\unit_decode/RegisterFile/n1719 ) );
  OAI22_X1 U2463 ( .A1(n928), .A2(n800), .B1(n922), .B2(\unit_decode/n1416 ), 
        .ZN(\unit_decode/RegisterFile/n1720 ) );
  OAI22_X1 U2464 ( .A1(n928), .A2(n797), .B1(n922), .B2(\unit_decode/n1417 ), 
        .ZN(\unit_decode/RegisterFile/n1721 ) );
  OAI22_X1 U2465 ( .A1(n928), .A2(n794), .B1(n922), .B2(\unit_decode/n1418 ), 
        .ZN(\unit_decode/RegisterFile/n1722 ) );
  OAI22_X1 U2466 ( .A1(n927), .A2(n791), .B1(n922), .B2(\unit_decode/n1419 ), 
        .ZN(\unit_decode/RegisterFile/n1723 ) );
  OAI22_X1 U2467 ( .A1(n927), .A2(n788), .B1(n922), .B2(\unit_decode/n1420 ), 
        .ZN(\unit_decode/RegisterFile/n1724 ) );
  OAI22_X1 U2468 ( .A1(n927), .A2(n785), .B1(n922), .B2(\unit_decode/n1421 ), 
        .ZN(\unit_decode/RegisterFile/n1725 ) );
  OAI22_X1 U2469 ( .A1(n927), .A2(n782), .B1(n922), .B2(\unit_decode/n1422 ), 
        .ZN(\unit_decode/RegisterFile/n1726 ) );
  OAI22_X1 U2470 ( .A1(n927), .A2(n779), .B1(n922), .B2(\unit_decode/n1423 ), 
        .ZN(\unit_decode/RegisterFile/n1727 ) );
  OAI22_X1 U2471 ( .A1(n926), .A2(n776), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1424 ), .ZN(\unit_decode/RegisterFile/n1728 ) );
  OAI22_X1 U2472 ( .A1(n926), .A2(n773), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1425 ), .ZN(\unit_decode/RegisterFile/n1729 ) );
  OAI22_X1 U2473 ( .A1(n926), .A2(n770), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1426 ), .ZN(\unit_decode/RegisterFile/n1730 ) );
  OAI22_X1 U2474 ( .A1(n926), .A2(n767), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1427 ), .ZN(\unit_decode/RegisterFile/n1731 ) );
  OAI22_X1 U2475 ( .A1(n926), .A2(n764), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1428 ), .ZN(\unit_decode/RegisterFile/n1732 ) );
  OAI22_X1 U2476 ( .A1(n925), .A2(n761), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1429 ), .ZN(\unit_decode/RegisterFile/n1733 ) );
  OAI22_X1 U2477 ( .A1(n925), .A2(n758), .B1(\unit_decode/n2251 ), .B2(
        \unit_decode/n1430 ), .ZN(\unit_decode/RegisterFile/n1734 ) );
  OAI22_X1 U2478 ( .A1(n925), .A2(n755), .B1(n922), .B2(\unit_decode/n1431 ), 
        .ZN(\unit_decode/RegisterFile/n1735 ) );
  OAI22_X1 U2479 ( .A1(n925), .A2(n752), .B1(n922), .B2(\unit_decode/n1432 ), 
        .ZN(\unit_decode/RegisterFile/n1736 ) );
  OAI22_X1 U2480 ( .A1(n925), .A2(n749), .B1(n922), .B2(\unit_decode/n1433 ), 
        .ZN(\unit_decode/RegisterFile/n1737 ) );
  OAI22_X1 U2481 ( .A1(n924), .A2(n746), .B1(n922), .B2(\unit_decode/n1434 ), 
        .ZN(\unit_decode/RegisterFile/n1738 ) );
  OAI22_X1 U2482 ( .A1(n924), .A2(n743), .B1(n922), .B2(\unit_decode/n1435 ), 
        .ZN(\unit_decode/RegisterFile/n1739 ) );
  OAI22_X1 U2483 ( .A1(n920), .A2(n812), .B1(n913), .B2(\unit_decode/n1436 ), 
        .ZN(\unit_decode/RegisterFile/n1748 ) );
  OAI22_X1 U2484 ( .A1(n920), .A2(n809), .B1(n913), .B2(\unit_decode/n1437 ), 
        .ZN(\unit_decode/RegisterFile/n1749 ) );
  OAI22_X1 U2485 ( .A1(n919), .A2(n806), .B1(n913), .B2(\unit_decode/n1438 ), 
        .ZN(\unit_decode/RegisterFile/n1750 ) );
  OAI22_X1 U2486 ( .A1(n919), .A2(n803), .B1(n913), .B2(\unit_decode/n1439 ), 
        .ZN(\unit_decode/RegisterFile/n1751 ) );
  OAI22_X1 U2487 ( .A1(n919), .A2(n800), .B1(n913), .B2(\unit_decode/n1440 ), 
        .ZN(\unit_decode/RegisterFile/n1752 ) );
  OAI22_X1 U2488 ( .A1(n919), .A2(n797), .B1(n913), .B2(\unit_decode/n1441 ), 
        .ZN(\unit_decode/RegisterFile/n1753 ) );
  OAI22_X1 U2489 ( .A1(n919), .A2(n794), .B1(n913), .B2(\unit_decode/n1442 ), 
        .ZN(\unit_decode/RegisterFile/n1754 ) );
  OAI22_X1 U2490 ( .A1(n918), .A2(n791), .B1(n913), .B2(\unit_decode/n1443 ), 
        .ZN(\unit_decode/RegisterFile/n1755 ) );
  OAI22_X1 U2491 ( .A1(n918), .A2(n788), .B1(n913), .B2(\unit_decode/n1444 ), 
        .ZN(\unit_decode/RegisterFile/n1756 ) );
  OAI22_X1 U2492 ( .A1(n918), .A2(n785), .B1(n913), .B2(\unit_decode/n1445 ), 
        .ZN(\unit_decode/RegisterFile/n1757 ) );
  OAI22_X1 U2493 ( .A1(n918), .A2(n782), .B1(n913), .B2(\unit_decode/n1446 ), 
        .ZN(\unit_decode/RegisterFile/n1758 ) );
  OAI22_X1 U2494 ( .A1(n918), .A2(n779), .B1(n913), .B2(\unit_decode/n1447 ), 
        .ZN(\unit_decode/RegisterFile/n1759 ) );
  OAI22_X1 U2495 ( .A1(n917), .A2(n776), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1448 ), .ZN(\unit_decode/RegisterFile/n1760 ) );
  OAI22_X1 U2496 ( .A1(n917), .A2(n773), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1449 ), .ZN(\unit_decode/RegisterFile/n1761 ) );
  OAI22_X1 U2497 ( .A1(n917), .A2(n770), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1450 ), .ZN(\unit_decode/RegisterFile/n1762 ) );
  OAI22_X1 U2498 ( .A1(n917), .A2(n767), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1451 ), .ZN(\unit_decode/RegisterFile/n1763 ) );
  OAI22_X1 U2499 ( .A1(n917), .A2(n764), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1452 ), .ZN(\unit_decode/RegisterFile/n1764 ) );
  OAI22_X1 U2500 ( .A1(n916), .A2(n761), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1453 ), .ZN(\unit_decode/RegisterFile/n1765 ) );
  OAI22_X1 U2501 ( .A1(n916), .A2(n758), .B1(\unit_decode/n2250 ), .B2(
        \unit_decode/n1454 ), .ZN(\unit_decode/RegisterFile/n1766 ) );
  OAI22_X1 U2502 ( .A1(n916), .A2(n755), .B1(n913), .B2(\unit_decode/n1455 ), 
        .ZN(\unit_decode/RegisterFile/n1767 ) );
  OAI22_X1 U2503 ( .A1(n916), .A2(n752), .B1(n913), .B2(\unit_decode/n1456 ), 
        .ZN(\unit_decode/RegisterFile/n1768 ) );
  OAI22_X1 U2504 ( .A1(n916), .A2(n749), .B1(n913), .B2(\unit_decode/n1457 ), 
        .ZN(\unit_decode/RegisterFile/n1769 ) );
  OAI22_X1 U2505 ( .A1(n915), .A2(n746), .B1(n913), .B2(\unit_decode/n1458 ), 
        .ZN(\unit_decode/RegisterFile/n1770 ) );
  OAI22_X1 U2506 ( .A1(n915), .A2(n743), .B1(n913), .B2(\unit_decode/n1459 ), 
        .ZN(\unit_decode/RegisterFile/n1771 ) );
  OAI22_X1 U2507 ( .A1(n893), .A2(n811), .B1(n886), .B2(\unit_decode/n1508 ), 
        .ZN(\unit_decode/RegisterFile/n1844 ) );
  OAI22_X1 U2508 ( .A1(n893), .A2(n808), .B1(n886), .B2(\unit_decode/n1509 ), 
        .ZN(\unit_decode/RegisterFile/n1845 ) );
  OAI22_X1 U2509 ( .A1(n892), .A2(n805), .B1(n886), .B2(\unit_decode/n1510 ), 
        .ZN(\unit_decode/RegisterFile/n1846 ) );
  OAI22_X1 U2510 ( .A1(n892), .A2(n802), .B1(n886), .B2(\unit_decode/n1511 ), 
        .ZN(\unit_decode/RegisterFile/n1847 ) );
  OAI22_X1 U2511 ( .A1(n892), .A2(n799), .B1(n886), .B2(\unit_decode/n1512 ), 
        .ZN(\unit_decode/RegisterFile/n1848 ) );
  OAI22_X1 U2512 ( .A1(n892), .A2(n796), .B1(n886), .B2(\unit_decode/n1513 ), 
        .ZN(\unit_decode/RegisterFile/n1849 ) );
  OAI22_X1 U2513 ( .A1(n892), .A2(n793), .B1(n886), .B2(\unit_decode/n1514 ), 
        .ZN(\unit_decode/RegisterFile/n1850 ) );
  OAI22_X1 U2514 ( .A1(n891), .A2(n790), .B1(n886), .B2(\unit_decode/n1515 ), 
        .ZN(\unit_decode/RegisterFile/n1851 ) );
  OAI22_X1 U2515 ( .A1(n891), .A2(n787), .B1(n886), .B2(\unit_decode/n1516 ), 
        .ZN(\unit_decode/RegisterFile/n1852 ) );
  OAI22_X1 U2516 ( .A1(n891), .A2(n784), .B1(n886), .B2(\unit_decode/n1517 ), 
        .ZN(\unit_decode/RegisterFile/n1853 ) );
  OAI22_X1 U2517 ( .A1(n891), .A2(n781), .B1(n886), .B2(\unit_decode/n1518 ), 
        .ZN(\unit_decode/RegisterFile/n1854 ) );
  OAI22_X1 U2518 ( .A1(n891), .A2(n778), .B1(n886), .B2(\unit_decode/n1519 ), 
        .ZN(\unit_decode/RegisterFile/n1855 ) );
  OAI22_X1 U2519 ( .A1(n890), .A2(n775), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1520 ), .ZN(\unit_decode/RegisterFile/n1856 ) );
  OAI22_X1 U2520 ( .A1(n890), .A2(n772), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1521 ), .ZN(\unit_decode/RegisterFile/n1857 ) );
  OAI22_X1 U2521 ( .A1(n890), .A2(n769), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1522 ), .ZN(\unit_decode/RegisterFile/n1858 ) );
  OAI22_X1 U2522 ( .A1(n890), .A2(n766), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1523 ), .ZN(\unit_decode/RegisterFile/n1859 ) );
  OAI22_X1 U2523 ( .A1(n890), .A2(n763), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1524 ), .ZN(\unit_decode/RegisterFile/n1860 ) );
  OAI22_X1 U2524 ( .A1(n889), .A2(n760), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1525 ), .ZN(\unit_decode/RegisterFile/n1861 ) );
  OAI22_X1 U2525 ( .A1(n889), .A2(n757), .B1(\unit_decode/n2247 ), .B2(
        \unit_decode/n1526 ), .ZN(\unit_decode/RegisterFile/n1862 ) );
  OAI22_X1 U2526 ( .A1(n889), .A2(n754), .B1(n886), .B2(\unit_decode/n1527 ), 
        .ZN(\unit_decode/RegisterFile/n1863 ) );
  OAI22_X1 U2527 ( .A1(n889), .A2(n751), .B1(n886), .B2(\unit_decode/n1528 ), 
        .ZN(\unit_decode/RegisterFile/n1864 ) );
  OAI22_X1 U2528 ( .A1(n889), .A2(n748), .B1(n886), .B2(\unit_decode/n1529 ), 
        .ZN(\unit_decode/RegisterFile/n1865 ) );
  OAI22_X1 U2529 ( .A1(n888), .A2(n745), .B1(n886), .B2(\unit_decode/n1530 ), 
        .ZN(\unit_decode/RegisterFile/n1866 ) );
  OAI22_X1 U2530 ( .A1(n888), .A2(n742), .B1(n886), .B2(\unit_decode/n1531 ), 
        .ZN(\unit_decode/RegisterFile/n1867 ) );
  OAI22_X1 U2531 ( .A1(n884), .A2(n811), .B1(n877), .B2(\unit_decode/n1532 ), 
        .ZN(\unit_decode/RegisterFile/n1876 ) );
  OAI22_X1 U2532 ( .A1(n884), .A2(n808), .B1(n877), .B2(\unit_decode/n1533 ), 
        .ZN(\unit_decode/RegisterFile/n1877 ) );
  OAI22_X1 U2533 ( .A1(n883), .A2(n805), .B1(n877), .B2(\unit_decode/n1534 ), 
        .ZN(\unit_decode/RegisterFile/n1878 ) );
  OAI22_X1 U2534 ( .A1(n883), .A2(n802), .B1(n877), .B2(\unit_decode/n1535 ), 
        .ZN(\unit_decode/RegisterFile/n1879 ) );
  OAI22_X1 U2535 ( .A1(n883), .A2(n799), .B1(n877), .B2(\unit_decode/n1536 ), 
        .ZN(\unit_decode/RegisterFile/n1880 ) );
  OAI22_X1 U2536 ( .A1(n883), .A2(n796), .B1(n877), .B2(\unit_decode/n1537 ), 
        .ZN(\unit_decode/RegisterFile/n1881 ) );
  OAI22_X1 U2537 ( .A1(n883), .A2(n793), .B1(n877), .B2(\unit_decode/n1538 ), 
        .ZN(\unit_decode/RegisterFile/n1882 ) );
  OAI22_X1 U2538 ( .A1(n882), .A2(n790), .B1(n877), .B2(\unit_decode/n1539 ), 
        .ZN(\unit_decode/RegisterFile/n1883 ) );
  OAI22_X1 U2539 ( .A1(n882), .A2(n787), .B1(n877), .B2(\unit_decode/n1540 ), 
        .ZN(\unit_decode/RegisterFile/n1884 ) );
  OAI22_X1 U2540 ( .A1(n882), .A2(n784), .B1(n877), .B2(\unit_decode/n1541 ), 
        .ZN(\unit_decode/RegisterFile/n1885 ) );
  OAI22_X1 U2541 ( .A1(n882), .A2(n781), .B1(n877), .B2(\unit_decode/n1542 ), 
        .ZN(\unit_decode/RegisterFile/n1886 ) );
  OAI22_X1 U2542 ( .A1(n882), .A2(n778), .B1(n877), .B2(\unit_decode/n1543 ), 
        .ZN(\unit_decode/RegisterFile/n1887 ) );
  OAI22_X1 U2543 ( .A1(n881), .A2(n775), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1544 ), .ZN(\unit_decode/RegisterFile/n1888 ) );
  OAI22_X1 U2544 ( .A1(n881), .A2(n772), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1545 ), .ZN(\unit_decode/RegisterFile/n1889 ) );
  OAI22_X1 U2545 ( .A1(n881), .A2(n769), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1546 ), .ZN(\unit_decode/RegisterFile/n1890 ) );
  OAI22_X1 U2546 ( .A1(n881), .A2(n766), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1547 ), .ZN(\unit_decode/RegisterFile/n1891 ) );
  OAI22_X1 U2547 ( .A1(n881), .A2(n763), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1548 ), .ZN(\unit_decode/RegisterFile/n1892 ) );
  OAI22_X1 U2548 ( .A1(n880), .A2(n760), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1549 ), .ZN(\unit_decode/RegisterFile/n1893 ) );
  OAI22_X1 U2549 ( .A1(n880), .A2(n757), .B1(\unit_decode/n2245 ), .B2(
        \unit_decode/n1550 ), .ZN(\unit_decode/RegisterFile/n1894 ) );
  OAI22_X1 U2550 ( .A1(n880), .A2(n754), .B1(n877), .B2(\unit_decode/n1551 ), 
        .ZN(\unit_decode/RegisterFile/n1895 ) );
  OAI22_X1 U2551 ( .A1(n880), .A2(n751), .B1(n877), .B2(\unit_decode/n1552 ), 
        .ZN(\unit_decode/RegisterFile/n1896 ) );
  OAI22_X1 U2552 ( .A1(n880), .A2(n748), .B1(n877), .B2(\unit_decode/n1553 ), 
        .ZN(\unit_decode/RegisterFile/n1897 ) );
  OAI22_X1 U2553 ( .A1(n879), .A2(n745), .B1(n877), .B2(\unit_decode/n1554 ), 
        .ZN(\unit_decode/RegisterFile/n1898 ) );
  OAI22_X1 U2554 ( .A1(n879), .A2(n742), .B1(n877), .B2(\unit_decode/n1555 ), 
        .ZN(\unit_decode/RegisterFile/n1899 ) );
  OAI22_X1 U2555 ( .A1(n857), .A2(n811), .B1(n850), .B2(\unit_decode/n1604 ), 
        .ZN(\unit_decode/RegisterFile/n1972 ) );
  OAI22_X1 U2556 ( .A1(n857), .A2(n808), .B1(n850), .B2(\unit_decode/n1605 ), 
        .ZN(\unit_decode/RegisterFile/n1973 ) );
  OAI22_X1 U2557 ( .A1(n856), .A2(n805), .B1(n850), .B2(\unit_decode/n1606 ), 
        .ZN(\unit_decode/RegisterFile/n1974 ) );
  OAI22_X1 U2558 ( .A1(n856), .A2(n802), .B1(n850), .B2(\unit_decode/n1607 ), 
        .ZN(\unit_decode/RegisterFile/n1975 ) );
  OAI22_X1 U2559 ( .A1(n856), .A2(n799), .B1(n850), .B2(\unit_decode/n1608 ), 
        .ZN(\unit_decode/RegisterFile/n1976 ) );
  OAI22_X1 U2560 ( .A1(n856), .A2(n796), .B1(n850), .B2(\unit_decode/n1609 ), 
        .ZN(\unit_decode/RegisterFile/n1977 ) );
  OAI22_X1 U2561 ( .A1(n856), .A2(n793), .B1(n850), .B2(\unit_decode/n1610 ), 
        .ZN(\unit_decode/RegisterFile/n1978 ) );
  OAI22_X1 U2562 ( .A1(n855), .A2(n790), .B1(n850), .B2(\unit_decode/n1611 ), 
        .ZN(\unit_decode/RegisterFile/n1979 ) );
  OAI22_X1 U2563 ( .A1(n855), .A2(n787), .B1(n850), .B2(\unit_decode/n1612 ), 
        .ZN(\unit_decode/RegisterFile/n1980 ) );
  OAI22_X1 U2564 ( .A1(n855), .A2(n784), .B1(n850), .B2(\unit_decode/n1613 ), 
        .ZN(\unit_decode/RegisterFile/n1981 ) );
  OAI22_X1 U2565 ( .A1(n855), .A2(n781), .B1(n850), .B2(\unit_decode/n1614 ), 
        .ZN(\unit_decode/RegisterFile/n1982 ) );
  OAI22_X1 U2566 ( .A1(n855), .A2(n778), .B1(n850), .B2(\unit_decode/n1615 ), 
        .ZN(\unit_decode/RegisterFile/n1983 ) );
  OAI22_X1 U2567 ( .A1(n854), .A2(n775), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1616 ), .ZN(\unit_decode/RegisterFile/n1984 ) );
  OAI22_X1 U2568 ( .A1(n854), .A2(n772), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1617 ), .ZN(\unit_decode/RegisterFile/n1985 ) );
  OAI22_X1 U2569 ( .A1(n854), .A2(n769), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1618 ), .ZN(\unit_decode/RegisterFile/n1986 ) );
  OAI22_X1 U2570 ( .A1(n854), .A2(n766), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1619 ), .ZN(\unit_decode/RegisterFile/n1987 ) );
  OAI22_X1 U2571 ( .A1(n854), .A2(n763), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1620 ), .ZN(\unit_decode/RegisterFile/n1988 ) );
  OAI22_X1 U2572 ( .A1(n853), .A2(n760), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1621 ), .ZN(\unit_decode/RegisterFile/n1989 ) );
  OAI22_X1 U2573 ( .A1(n853), .A2(n757), .B1(\unit_decode/n2238 ), .B2(
        \unit_decode/n1622 ), .ZN(\unit_decode/RegisterFile/n1990 ) );
  OAI22_X1 U2574 ( .A1(n853), .A2(n754), .B1(n850), .B2(\unit_decode/n1623 ), 
        .ZN(\unit_decode/RegisterFile/n1991 ) );
  OAI22_X1 U2575 ( .A1(n853), .A2(n751), .B1(n850), .B2(\unit_decode/n1624 ), 
        .ZN(\unit_decode/RegisterFile/n1992 ) );
  OAI22_X1 U2576 ( .A1(n853), .A2(n748), .B1(n850), .B2(\unit_decode/n1625 ), 
        .ZN(\unit_decode/RegisterFile/n1993 ) );
  OAI22_X1 U2577 ( .A1(n852), .A2(n745), .B1(n850), .B2(\unit_decode/n1626 ), 
        .ZN(\unit_decode/RegisterFile/n1994 ) );
  OAI22_X1 U2578 ( .A1(n852), .A2(n742), .B1(n850), .B2(\unit_decode/n1627 ), 
        .ZN(\unit_decode/RegisterFile/n1995 ) );
  OAI22_X1 U2579 ( .A1(n848), .A2(n811), .B1(n841), .B2(\unit_decode/n1628 ), 
        .ZN(\unit_decode/RegisterFile/n2004 ) );
  OAI22_X1 U2580 ( .A1(n848), .A2(n808), .B1(n841), .B2(\unit_decode/n1629 ), 
        .ZN(\unit_decode/RegisterFile/n2005 ) );
  OAI22_X1 U2581 ( .A1(n847), .A2(n805), .B1(n841), .B2(\unit_decode/n1630 ), 
        .ZN(\unit_decode/RegisterFile/n2006 ) );
  OAI22_X1 U2582 ( .A1(n847), .A2(n802), .B1(n841), .B2(\unit_decode/n1631 ), 
        .ZN(\unit_decode/RegisterFile/n2007 ) );
  OAI22_X1 U2583 ( .A1(n847), .A2(n799), .B1(n841), .B2(\unit_decode/n1632 ), 
        .ZN(\unit_decode/RegisterFile/n2008 ) );
  OAI22_X1 U2584 ( .A1(n847), .A2(n796), .B1(n841), .B2(\unit_decode/n1633 ), 
        .ZN(\unit_decode/RegisterFile/n2009 ) );
  OAI22_X1 U2585 ( .A1(n847), .A2(n793), .B1(n841), .B2(\unit_decode/n1634 ), 
        .ZN(\unit_decode/RegisterFile/n2010 ) );
  OAI22_X1 U2586 ( .A1(n846), .A2(n790), .B1(n841), .B2(\unit_decode/n1635 ), 
        .ZN(\unit_decode/RegisterFile/n2011 ) );
  OAI22_X1 U2587 ( .A1(n846), .A2(n787), .B1(n841), .B2(\unit_decode/n1636 ), 
        .ZN(\unit_decode/RegisterFile/n2012 ) );
  OAI22_X1 U2588 ( .A1(n846), .A2(n784), .B1(n841), .B2(\unit_decode/n1637 ), 
        .ZN(\unit_decode/RegisterFile/n2013 ) );
  OAI22_X1 U2589 ( .A1(n846), .A2(n781), .B1(n841), .B2(\unit_decode/n1638 ), 
        .ZN(\unit_decode/RegisterFile/n2014 ) );
  OAI22_X1 U2590 ( .A1(n846), .A2(n778), .B1(n841), .B2(\unit_decode/n1639 ), 
        .ZN(\unit_decode/RegisterFile/n2015 ) );
  OAI22_X1 U2591 ( .A1(n845), .A2(n775), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1640 ), .ZN(\unit_decode/RegisterFile/n2016 ) );
  OAI22_X1 U2592 ( .A1(n845), .A2(n772), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1641 ), .ZN(\unit_decode/RegisterFile/n2017 ) );
  OAI22_X1 U2593 ( .A1(n845), .A2(n769), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1642 ), .ZN(\unit_decode/RegisterFile/n2018 ) );
  OAI22_X1 U2594 ( .A1(n845), .A2(n766), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1643 ), .ZN(\unit_decode/RegisterFile/n2019 ) );
  OAI22_X1 U2595 ( .A1(n845), .A2(n763), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1644 ), .ZN(\unit_decode/RegisterFile/n2020 ) );
  OAI22_X1 U2596 ( .A1(n844), .A2(n760), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1645 ), .ZN(\unit_decode/RegisterFile/n2021 ) );
  OAI22_X1 U2597 ( .A1(n844), .A2(n757), .B1(\unit_decode/n2236 ), .B2(
        \unit_decode/n1646 ), .ZN(\unit_decode/RegisterFile/n2022 ) );
  OAI22_X1 U2598 ( .A1(n844), .A2(n754), .B1(n841), .B2(\unit_decode/n1647 ), 
        .ZN(\unit_decode/RegisterFile/n2023 ) );
  OAI22_X1 U2599 ( .A1(n844), .A2(n751), .B1(n841), .B2(\unit_decode/n1648 ), 
        .ZN(\unit_decode/RegisterFile/n2024 ) );
  OAI22_X1 U2600 ( .A1(n844), .A2(n748), .B1(n841), .B2(\unit_decode/n1649 ), 
        .ZN(\unit_decode/RegisterFile/n2025 ) );
  OAI22_X1 U2601 ( .A1(n843), .A2(n745), .B1(n841), .B2(\unit_decode/n1650 ), 
        .ZN(\unit_decode/RegisterFile/n2026 ) );
  OAI22_X1 U2602 ( .A1(n843), .A2(n742), .B1(n841), .B2(\unit_decode/n1651 ), 
        .ZN(\unit_decode/RegisterFile/n2027 ) );
  OAI22_X1 U2603 ( .A1(n821), .A2(n811), .B1(n814), .B2(\unit_decode/n1700 ), 
        .ZN(\unit_decode/RegisterFile/n2100 ) );
  OAI22_X1 U2604 ( .A1(n821), .A2(n808), .B1(n814), .B2(\unit_decode/n1701 ), 
        .ZN(\unit_decode/RegisterFile/n2101 ) );
  OAI22_X1 U2605 ( .A1(n820), .A2(n805), .B1(n814), .B2(\unit_decode/n1702 ), 
        .ZN(\unit_decode/RegisterFile/n2102 ) );
  OAI22_X1 U2606 ( .A1(n820), .A2(n802), .B1(n814), .B2(\unit_decode/n1703 ), 
        .ZN(\unit_decode/RegisterFile/n2103 ) );
  OAI22_X1 U2607 ( .A1(n820), .A2(n799), .B1(n814), .B2(\unit_decode/n1704 ), 
        .ZN(\unit_decode/RegisterFile/n2104 ) );
  OAI22_X1 U2608 ( .A1(n820), .A2(n796), .B1(n814), .B2(\unit_decode/n1705 ), 
        .ZN(\unit_decode/RegisterFile/n2105 ) );
  OAI22_X1 U2609 ( .A1(n820), .A2(n793), .B1(n814), .B2(\unit_decode/n1706 ), 
        .ZN(\unit_decode/RegisterFile/n2106 ) );
  OAI22_X1 U2610 ( .A1(n819), .A2(n790), .B1(n814), .B2(\unit_decode/n1707 ), 
        .ZN(\unit_decode/RegisterFile/n2107 ) );
  OAI22_X1 U2611 ( .A1(n819), .A2(n787), .B1(n814), .B2(\unit_decode/n1708 ), 
        .ZN(\unit_decode/RegisterFile/n2108 ) );
  OAI22_X1 U2612 ( .A1(n819), .A2(n784), .B1(n814), .B2(\unit_decode/n1709 ), 
        .ZN(\unit_decode/RegisterFile/n2109 ) );
  OAI22_X1 U2613 ( .A1(n819), .A2(n781), .B1(n814), .B2(\unit_decode/n1710 ), 
        .ZN(\unit_decode/RegisterFile/n2110 ) );
  OAI22_X1 U2614 ( .A1(n819), .A2(n778), .B1(n814), .B2(\unit_decode/n1711 ), 
        .ZN(\unit_decode/RegisterFile/n2111 ) );
  OAI22_X1 U2615 ( .A1(n818), .A2(n775), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1712 ), .ZN(\unit_decode/RegisterFile/n2112 ) );
  OAI22_X1 U2616 ( .A1(n818), .A2(n772), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1713 ), .ZN(\unit_decode/RegisterFile/n2113 ) );
  OAI22_X1 U2617 ( .A1(n818), .A2(n769), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1714 ), .ZN(\unit_decode/RegisterFile/n2114 ) );
  OAI22_X1 U2618 ( .A1(n818), .A2(n766), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1715 ), .ZN(\unit_decode/RegisterFile/n2115 ) );
  OAI22_X1 U2619 ( .A1(n818), .A2(n763), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1716 ), .ZN(\unit_decode/RegisterFile/n2116 ) );
  OAI22_X1 U2620 ( .A1(n817), .A2(n760), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1717 ), .ZN(\unit_decode/RegisterFile/n2117 ) );
  OAI22_X1 U2621 ( .A1(n817), .A2(n757), .B1(\unit_decode/n2230 ), .B2(
        \unit_decode/n1718 ), .ZN(\unit_decode/RegisterFile/n2118 ) );
  OAI22_X1 U2622 ( .A1(n817), .A2(n754), .B1(n814), .B2(\unit_decode/n1719 ), 
        .ZN(\unit_decode/RegisterFile/n2119 ) );
  OAI22_X1 U2623 ( .A1(n817), .A2(n751), .B1(n814), .B2(\unit_decode/n1720 ), 
        .ZN(\unit_decode/RegisterFile/n2120 ) );
  OAI22_X1 U2624 ( .A1(n817), .A2(n748), .B1(n814), .B2(\unit_decode/n1721 ), 
        .ZN(\unit_decode/RegisterFile/n2121 ) );
  OAI22_X1 U2625 ( .A1(n816), .A2(n745), .B1(n814), .B2(\unit_decode/n1722 ), 
        .ZN(\unit_decode/RegisterFile/n2122 ) );
  OAI22_X1 U2626 ( .A1(n816), .A2(n742), .B1(n814), .B2(\unit_decode/n1723 ), 
        .ZN(\unit_decode/RegisterFile/n2123 ) );
  OAI22_X1 U2627 ( .A1(n719), .A2(n811), .B1(n712), .B2(\unit_decode/n1724 ), 
        .ZN(\unit_decode/RegisterFile/n2132 ) );
  OAI22_X1 U2628 ( .A1(n719), .A2(n808), .B1(n712), .B2(\unit_decode/n1725 ), 
        .ZN(\unit_decode/RegisterFile/n2133 ) );
  OAI22_X1 U2629 ( .A1(n718), .A2(n805), .B1(n712), .B2(\unit_decode/n1726 ), 
        .ZN(\unit_decode/RegisterFile/n2134 ) );
  OAI22_X1 U2630 ( .A1(n718), .A2(n802), .B1(n712), .B2(\unit_decode/n1727 ), 
        .ZN(\unit_decode/RegisterFile/n2135 ) );
  OAI22_X1 U2631 ( .A1(n718), .A2(n799), .B1(n712), .B2(\unit_decode/n1728 ), 
        .ZN(\unit_decode/RegisterFile/n2136 ) );
  OAI22_X1 U2632 ( .A1(n718), .A2(n796), .B1(n712), .B2(\unit_decode/n1729 ), 
        .ZN(\unit_decode/RegisterFile/n2137 ) );
  OAI22_X1 U2633 ( .A1(n718), .A2(n793), .B1(n712), .B2(\unit_decode/n1730 ), 
        .ZN(\unit_decode/RegisterFile/n2138 ) );
  OAI22_X1 U2634 ( .A1(n717), .A2(n790), .B1(n712), .B2(\unit_decode/n1731 ), 
        .ZN(\unit_decode/RegisterFile/n2139 ) );
  OAI22_X1 U2635 ( .A1(n717), .A2(n787), .B1(n712), .B2(\unit_decode/n1732 ), 
        .ZN(\unit_decode/RegisterFile/n2140 ) );
  OAI22_X1 U2636 ( .A1(n717), .A2(n784), .B1(n712), .B2(\unit_decode/n1733 ), 
        .ZN(\unit_decode/RegisterFile/n2141 ) );
  OAI22_X1 U2637 ( .A1(n717), .A2(n781), .B1(n712), .B2(\unit_decode/n1734 ), 
        .ZN(\unit_decode/RegisterFile/n2142 ) );
  OAI22_X1 U2638 ( .A1(n717), .A2(n778), .B1(n712), .B2(\unit_decode/n1735 ), 
        .ZN(\unit_decode/RegisterFile/n2143 ) );
  OAI22_X1 U2639 ( .A1(n716), .A2(n775), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1736 ), .ZN(\unit_decode/RegisterFile/n2144 ) );
  OAI22_X1 U2640 ( .A1(n716), .A2(n772), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1737 ), .ZN(\unit_decode/RegisterFile/n2145 ) );
  OAI22_X1 U2641 ( .A1(n716), .A2(n769), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1738 ), .ZN(\unit_decode/RegisterFile/n2146 ) );
  OAI22_X1 U2642 ( .A1(n716), .A2(n766), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1739 ), .ZN(\unit_decode/RegisterFile/n2147 ) );
  OAI22_X1 U2643 ( .A1(n716), .A2(n763), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1740 ), .ZN(\unit_decode/RegisterFile/n2148 ) );
  OAI22_X1 U2644 ( .A1(n715), .A2(n760), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1741 ), .ZN(\unit_decode/RegisterFile/n2149 ) );
  OAI22_X1 U2645 ( .A1(n715), .A2(n757), .B1(\unit_decode/n2196 ), .B2(
        \unit_decode/n1742 ), .ZN(\unit_decode/RegisterFile/n2150 ) );
  OAI22_X1 U2646 ( .A1(n715), .A2(n754), .B1(n712), .B2(\unit_decode/n1743 ), 
        .ZN(\unit_decode/RegisterFile/n2151 ) );
  OAI22_X1 U2647 ( .A1(n715), .A2(n751), .B1(n712), .B2(\unit_decode/n1744 ), 
        .ZN(\unit_decode/RegisterFile/n2152 ) );
  OAI22_X1 U2648 ( .A1(n715), .A2(n748), .B1(n712), .B2(\unit_decode/n1745 ), 
        .ZN(\unit_decode/RegisterFile/n2153 ) );
  OAI22_X1 U2649 ( .A1(n714), .A2(n745), .B1(n712), .B2(\unit_decode/n1746 ), 
        .ZN(\unit_decode/RegisterFile/n2154 ) );
  OAI22_X1 U2650 ( .A1(n714), .A2(n742), .B1(n712), .B2(\unit_decode/n1747 ), 
        .ZN(\unit_decode/RegisterFile/n2155 ) );
  OAI22_X1 U2651 ( .A1(n1090), .A2(\unit_decode/n1173 ), .B1(n1084), .B2(n789), 
        .ZN(\unit_decode/RegisterFile/n1148 ) );
  OAI22_X1 U2652 ( .A1(n1090), .A2(\unit_decode/n1174 ), .B1(n1084), .B2(n786), 
        .ZN(\unit_decode/RegisterFile/n1149 ) );
  OAI22_X1 U2653 ( .A1(n1090), .A2(\unit_decode/n1175 ), .B1(n1084), .B2(n783), 
        .ZN(\unit_decode/RegisterFile/n1150 ) );
  OAI22_X1 U2654 ( .A1(n1090), .A2(\unit_decode/n1176 ), .B1(n1084), .B2(n780), 
        .ZN(\unit_decode/RegisterFile/n1151 ) );
  OAI22_X1 U2655 ( .A1(n1089), .A2(\unit_decode/n1177 ), .B1(n1085), .B2(n777), 
        .ZN(\unit_decode/RegisterFile/n1152 ) );
  OAI22_X1 U2656 ( .A1(n1089), .A2(\unit_decode/n1178 ), .B1(n1085), .B2(n774), 
        .ZN(\unit_decode/RegisterFile/n1153 ) );
  OAI22_X1 U2657 ( .A1(n1089), .A2(\unit_decode/n1179 ), .B1(n1085), .B2(n771), 
        .ZN(\unit_decode/RegisterFile/n1154 ) );
  OAI22_X1 U2658 ( .A1(n1089), .A2(\unit_decode/n1180 ), .B1(n1085), .B2(n768), 
        .ZN(\unit_decode/RegisterFile/n1155 ) );
  OAI22_X1 U2659 ( .A1(n1089), .A2(\unit_decode/n1181 ), .B1(n1085), .B2(n765), 
        .ZN(\unit_decode/RegisterFile/n1156 ) );
  OAI22_X1 U2660 ( .A1(n1088), .A2(\unit_decode/n1182 ), .B1(n1085), .B2(n762), 
        .ZN(\unit_decode/RegisterFile/n1157 ) );
  OAI22_X1 U2661 ( .A1(n1088), .A2(\unit_decode/n1183 ), .B1(n1085), .B2(n759), 
        .ZN(\unit_decode/RegisterFile/n1158 ) );
  OAI22_X1 U2662 ( .A1(n1088), .A2(\unit_decode/n1184 ), .B1(n1085), .B2(n756), 
        .ZN(\unit_decode/RegisterFile/n1159 ) );
  OAI22_X1 U2663 ( .A1(n1088), .A2(\unit_decode/n1185 ), .B1(n1085), .B2(n753), 
        .ZN(\unit_decode/RegisterFile/n1160 ) );
  OAI22_X1 U2664 ( .A1(n1088), .A2(\unit_decode/n1186 ), .B1(n1085), .B2(n750), 
        .ZN(\unit_decode/RegisterFile/n1161 ) );
  OAI22_X1 U2665 ( .A1(n1087), .A2(\unit_decode/n1187 ), .B1(n1085), .B2(n747), 
        .ZN(\unit_decode/RegisterFile/n1162 ) );
  OAI22_X1 U2666 ( .A1(n1087), .A2(\unit_decode/n1188 ), .B1(n1085), .B2(n744), 
        .ZN(\unit_decode/RegisterFile/n1163 ) );
  OAI22_X1 U2667 ( .A1(n1090), .A2(\unit_decode/n1956 ), .B1(n1084), .B2(n792), 
        .ZN(\unit_decode/RegisterFile/n1147 ) );
  OAI22_X1 U2668 ( .A1(n1091), .A2(\unit_decode/n1957 ), .B1(n1084), .B2(n795), 
        .ZN(\unit_decode/RegisterFile/n1146 ) );
  OAI22_X1 U2669 ( .A1(n1091), .A2(\unit_decode/n1958 ), .B1(n1084), .B2(n798), 
        .ZN(\unit_decode/RegisterFile/n1145 ) );
  OAI22_X1 U2670 ( .A1(n1091), .A2(\unit_decode/n1959 ), .B1(n1084), .B2(n801), 
        .ZN(\unit_decode/RegisterFile/n1144 ) );
  OAI22_X1 U2671 ( .A1(n1091), .A2(\unit_decode/n1960 ), .B1(n1084), .B2(n804), 
        .ZN(\unit_decode/RegisterFile/n1143 ) );
  OAI22_X1 U2672 ( .A1(n1091), .A2(\unit_decode/n1961 ), .B1(n1084), .B2(n807), 
        .ZN(\unit_decode/RegisterFile/n1142 ) );
  OAI22_X1 U2673 ( .A1(n1092), .A2(\unit_decode/n1962 ), .B1(n1084), .B2(n810), 
        .ZN(\unit_decode/RegisterFile/n1141 ) );
  OAI22_X1 U2674 ( .A1(n1092), .A2(\unit_decode/n1963 ), .B1(n1084), .B2(n813), 
        .ZN(\unit_decode/RegisterFile/n1140 ) );
  OAI22_X1 U2675 ( .A1(n1058), .A2(n711), .B1(\unit_decode/RegisterFile/n3868 ), .B2(n1057), .ZN(\unit_decode/RegisterFile/n1267 ) );
  OAI22_X1 U2676 ( .A1(n1058), .A2(n723), .B1(\unit_decode/RegisterFile/n3869 ), .B2(n1057), .ZN(\unit_decode/RegisterFile/n1266 ) );
  OAI22_X1 U2677 ( .A1(n1058), .A2(n726), .B1(\unit_decode/RegisterFile/n3870 ), .B2(\unit_decode/n2268 ), .ZN(\unit_decode/RegisterFile/n1265 ) );
  OAI22_X1 U2678 ( .A1(n1040), .A2(n711), .B1(\unit_decode/RegisterFile/n3804 ), .B2(n1039), .ZN(\unit_decode/RegisterFile/n1331 ) );
  OAI22_X1 U2679 ( .A1(n1040), .A2(n723), .B1(\unit_decode/RegisterFile/n3805 ), .B2(n1039), .ZN(\unit_decode/RegisterFile/n1330 ) );
  OAI22_X1 U2680 ( .A1(n1040), .A2(n726), .B1(\unit_decode/RegisterFile/n3806 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1329 ) );
  OAI22_X1 U2681 ( .A1(n1040), .A2(n729), .B1(\unit_decode/RegisterFile/n3807 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1328 ) );
  OAI22_X1 U2682 ( .A1(n1040), .A2(n732), .B1(\unit_decode/RegisterFile/n3808 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1327 ) );
  OAI22_X1 U2683 ( .A1(n1041), .A2(n735), .B1(\unit_decode/RegisterFile/n3809 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1326 ) );
  OAI22_X1 U2684 ( .A1(n1041), .A2(n738), .B1(\unit_decode/RegisterFile/n3810 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1325 ) );
  OAI22_X1 U2685 ( .A1(n1041), .A2(n741), .B1(\unit_decode/RegisterFile/n3811 ), .B2(\unit_decode/n2266 ), .ZN(\unit_decode/RegisterFile/n1324 ) );
  OAI22_X1 U2686 ( .A1(n1005), .A2(n743), .B1(\unit_decode/RegisterFile/n3684 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1451 ) );
  OAI22_X1 U2687 ( .A1(n1005), .A2(n746), .B1(\unit_decode/RegisterFile/n3685 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1450 ) );
  OAI22_X1 U2688 ( .A1(n1006), .A2(n749), .B1(\unit_decode/RegisterFile/n3686 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1449 ) );
  OAI22_X1 U2689 ( .A1(n1006), .A2(n752), .B1(\unit_decode/RegisterFile/n3687 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1448 ) );
  OAI22_X1 U2690 ( .A1(n1006), .A2(n755), .B1(\unit_decode/RegisterFile/n3688 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1447 ) );
  OAI22_X1 U2691 ( .A1(n1006), .A2(n758), .B1(\unit_decode/RegisterFile/n3689 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1446 ) );
  OAI22_X1 U2692 ( .A1(n1006), .A2(n761), .B1(\unit_decode/RegisterFile/n3690 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1445 ) );
  OAI22_X1 U2693 ( .A1(n1007), .A2(n764), .B1(\unit_decode/RegisterFile/n3691 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1444 ) );
  OAI22_X1 U2694 ( .A1(n1007), .A2(n767), .B1(\unit_decode/RegisterFile/n3692 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1443 ) );
  OAI22_X1 U2695 ( .A1(n1007), .A2(n770), .B1(\unit_decode/RegisterFile/n3693 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1442 ) );
  OAI22_X1 U2696 ( .A1(n1007), .A2(n773), .B1(\unit_decode/RegisterFile/n3694 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1441 ) );
  OAI22_X1 U2697 ( .A1(n1007), .A2(n776), .B1(\unit_decode/RegisterFile/n3695 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1440 ) );
  OAI22_X1 U2698 ( .A1(n1008), .A2(n779), .B1(\unit_decode/RegisterFile/n3696 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1439 ) );
  OAI22_X1 U2699 ( .A1(n1008), .A2(n782), .B1(\unit_decode/RegisterFile/n3697 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1438 ) );
  OAI22_X1 U2700 ( .A1(n1008), .A2(n785), .B1(\unit_decode/RegisterFile/n3698 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1437 ) );
  OAI22_X1 U2701 ( .A1(n1008), .A2(n788), .B1(\unit_decode/RegisterFile/n3699 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1436 ) );
  OAI22_X1 U2702 ( .A1(n1008), .A2(n791), .B1(\unit_decode/RegisterFile/n3700 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1435 ) );
  OAI22_X1 U2703 ( .A1(n1009), .A2(n794), .B1(\unit_decode/RegisterFile/n3701 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1434 ) );
  OAI22_X1 U2704 ( .A1(n1009), .A2(n797), .B1(\unit_decode/RegisterFile/n3702 ), .B2(\unit_decode/n2261 ), .ZN(\unit_decode/RegisterFile/n1433 ) );
  OAI22_X1 U2705 ( .A1(n1009), .A2(n800), .B1(\unit_decode/RegisterFile/n3703 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1432 ) );
  OAI22_X1 U2706 ( .A1(n1009), .A2(n803), .B1(\unit_decode/RegisterFile/n3704 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1431 ) );
  OAI22_X1 U2707 ( .A1(n1009), .A2(n806), .B1(\unit_decode/RegisterFile/n3705 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1430 ) );
  OAI22_X1 U2708 ( .A1(n1010), .A2(n809), .B1(\unit_decode/RegisterFile/n3706 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1429 ) );
  OAI22_X1 U2709 ( .A1(n1010), .A2(n812), .B1(\unit_decode/RegisterFile/n3707 ), .B2(n1003), .ZN(\unit_decode/RegisterFile/n1428 ) );
  OAI22_X1 U2710 ( .A1(n950), .A2(n710), .B1(\unit_decode/RegisterFile/n3484 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1651 ) );
  OAI22_X1 U2711 ( .A1(n950), .A2(n722), .B1(\unit_decode/RegisterFile/n3485 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1650 ) );
  OAI22_X1 U2712 ( .A1(n950), .A2(n725), .B1(\unit_decode/RegisterFile/n3486 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1649 ) );
  OAI22_X1 U2713 ( .A1(n1014), .A2(n743), .B1(\unit_decode/RegisterFile/n3716 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1419 ) );
  OAI22_X1 U2714 ( .A1(n1014), .A2(n746), .B1(\unit_decode/RegisterFile/n3717 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1418 ) );
  OAI22_X1 U2715 ( .A1(n1015), .A2(n749), .B1(\unit_decode/RegisterFile/n3718 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1417 ) );
  OAI22_X1 U2716 ( .A1(n1015), .A2(n752), .B1(\unit_decode/RegisterFile/n3719 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1416 ) );
  OAI22_X1 U2717 ( .A1(n1015), .A2(n755), .B1(\unit_decode/RegisterFile/n3720 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1415 ) );
  OAI22_X1 U2718 ( .A1(n1015), .A2(n758), .B1(\unit_decode/RegisterFile/n3721 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1414 ) );
  OAI22_X1 U2719 ( .A1(n1015), .A2(n761), .B1(\unit_decode/RegisterFile/n3722 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1413 ) );
  OAI22_X1 U2720 ( .A1(n1016), .A2(n764), .B1(\unit_decode/RegisterFile/n3723 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1412 ) );
  OAI22_X1 U2721 ( .A1(n1016), .A2(n767), .B1(\unit_decode/RegisterFile/n3724 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1411 ) );
  OAI22_X1 U2722 ( .A1(n1016), .A2(n770), .B1(\unit_decode/RegisterFile/n3725 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1410 ) );
  OAI22_X1 U2723 ( .A1(n1016), .A2(n773), .B1(\unit_decode/RegisterFile/n3726 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1409 ) );
  OAI22_X1 U2724 ( .A1(n1016), .A2(n776), .B1(\unit_decode/RegisterFile/n3727 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1408 ) );
  OAI22_X1 U2725 ( .A1(n1017), .A2(n779), .B1(\unit_decode/RegisterFile/n3728 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1407 ) );
  OAI22_X1 U2726 ( .A1(n1017), .A2(n782), .B1(\unit_decode/RegisterFile/n3729 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1406 ) );
  OAI22_X1 U2727 ( .A1(n1017), .A2(n785), .B1(\unit_decode/RegisterFile/n3730 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1405 ) );
  OAI22_X1 U2728 ( .A1(n1017), .A2(n788), .B1(\unit_decode/RegisterFile/n3731 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1404 ) );
  OAI22_X1 U2729 ( .A1(n1017), .A2(n791), .B1(\unit_decode/RegisterFile/n3732 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1403 ) );
  OAI22_X1 U2730 ( .A1(n1018), .A2(n794), .B1(\unit_decode/RegisterFile/n3733 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1402 ) );
  OAI22_X1 U2731 ( .A1(n1018), .A2(n797), .B1(\unit_decode/RegisterFile/n3734 ), .B2(\unit_decode/n2262 ), .ZN(\unit_decode/RegisterFile/n1401 ) );
  OAI22_X1 U2732 ( .A1(n1018), .A2(n800), .B1(\unit_decode/RegisterFile/n3735 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1400 ) );
  OAI22_X1 U2733 ( .A1(n1018), .A2(n803), .B1(\unit_decode/RegisterFile/n3736 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1399 ) );
  OAI22_X1 U2734 ( .A1(n1018), .A2(n806), .B1(\unit_decode/RegisterFile/n3737 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1398 ) );
  OAI22_X1 U2735 ( .A1(n1019), .A2(n809), .B1(\unit_decode/RegisterFile/n3738 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1397 ) );
  OAI22_X1 U2736 ( .A1(n1019), .A2(n812), .B1(\unit_decode/RegisterFile/n3739 ), .B2(n1012), .ZN(\unit_decode/RegisterFile/n1396 ) );
  OAI22_X1 U2737 ( .A1(n996), .A2(n743), .B1(\unit_decode/RegisterFile/n3652 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1483 ) );
  OAI22_X1 U2738 ( .A1(n996), .A2(n746), .B1(\unit_decode/RegisterFile/n3653 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1482 ) );
  OAI22_X1 U2739 ( .A1(n997), .A2(n749), .B1(\unit_decode/RegisterFile/n3654 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1481 ) );
  OAI22_X1 U2740 ( .A1(n997), .A2(n752), .B1(\unit_decode/RegisterFile/n3655 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1480 ) );
  OAI22_X1 U2741 ( .A1(n997), .A2(n755), .B1(\unit_decode/RegisterFile/n3656 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1479 ) );
  OAI22_X1 U2742 ( .A1(n997), .A2(n758), .B1(\unit_decode/RegisterFile/n3657 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1478 ) );
  OAI22_X1 U2743 ( .A1(n997), .A2(n761), .B1(\unit_decode/RegisterFile/n3658 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1477 ) );
  OAI22_X1 U2744 ( .A1(n998), .A2(n764), .B1(\unit_decode/RegisterFile/n3659 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1476 ) );
  OAI22_X1 U2745 ( .A1(n998), .A2(n767), .B1(\unit_decode/RegisterFile/n3660 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1475 ) );
  OAI22_X1 U2746 ( .A1(n998), .A2(n770), .B1(\unit_decode/RegisterFile/n3661 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1474 ) );
  OAI22_X1 U2747 ( .A1(n998), .A2(n773), .B1(\unit_decode/RegisterFile/n3662 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1473 ) );
  OAI22_X1 U2748 ( .A1(n998), .A2(n776), .B1(\unit_decode/RegisterFile/n3663 ), 
        .B2(n994), .ZN(\unit_decode/RegisterFile/n1472 ) );
  OAI22_X1 U2749 ( .A1(n999), .A2(n779), .B1(\unit_decode/RegisterFile/n3664 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1471 ) );
  OAI22_X1 U2750 ( .A1(n999), .A2(n782), .B1(\unit_decode/RegisterFile/n3665 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1470 ) );
  OAI22_X1 U2751 ( .A1(n999), .A2(n785), .B1(\unit_decode/RegisterFile/n3666 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1469 ) );
  OAI22_X1 U2752 ( .A1(n999), .A2(n788), .B1(\unit_decode/RegisterFile/n3667 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1468 ) );
  OAI22_X1 U2753 ( .A1(n999), .A2(n791), .B1(\unit_decode/RegisterFile/n3668 ), 
        .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1467 ) );
  OAI22_X1 U2754 ( .A1(n1000), .A2(n794), .B1(\unit_decode/RegisterFile/n3669 ), .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1466 ) );
  OAI22_X1 U2755 ( .A1(n1000), .A2(n797), .B1(\unit_decode/RegisterFile/n3670 ), .B2(\unit_decode/n2260 ), .ZN(\unit_decode/RegisterFile/n1465 ) );
  OAI22_X1 U2756 ( .A1(n1000), .A2(n800), .B1(\unit_decode/RegisterFile/n3671 ), .B2(n994), .ZN(\unit_decode/RegisterFile/n1464 ) );
  OAI22_X1 U2757 ( .A1(n1000), .A2(n803), .B1(\unit_decode/RegisterFile/n3672 ), .B2(n994), .ZN(\unit_decode/RegisterFile/n1463 ) );
  OAI22_X1 U2758 ( .A1(n1000), .A2(n806), .B1(\unit_decode/RegisterFile/n3673 ), .B2(n994), .ZN(\unit_decode/RegisterFile/n1462 ) );
  OAI22_X1 U2759 ( .A1(n1001), .A2(n809), .B1(\unit_decode/RegisterFile/n3674 ), .B2(n994), .ZN(\unit_decode/RegisterFile/n1461 ) );
  OAI22_X1 U2760 ( .A1(n1001), .A2(n812), .B1(\unit_decode/RegisterFile/n3675 ), .B2(n994), .ZN(\unit_decode/RegisterFile/n1460 ) );
  OAI22_X1 U2761 ( .A1(n987), .A2(n743), .B1(\unit_decode/RegisterFile/n3620 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1515 ) );
  OAI22_X1 U2762 ( .A1(n987), .A2(n746), .B1(\unit_decode/RegisterFile/n3621 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1514 ) );
  OAI22_X1 U2763 ( .A1(n988), .A2(n749), .B1(\unit_decode/RegisterFile/n3622 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1513 ) );
  OAI22_X1 U2764 ( .A1(n988), .A2(n752), .B1(\unit_decode/RegisterFile/n3623 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1512 ) );
  OAI22_X1 U2765 ( .A1(n988), .A2(n755), .B1(\unit_decode/RegisterFile/n3624 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1511 ) );
  OAI22_X1 U2766 ( .A1(n988), .A2(n758), .B1(\unit_decode/RegisterFile/n3625 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1510 ) );
  OAI22_X1 U2767 ( .A1(n988), .A2(n761), .B1(\unit_decode/RegisterFile/n3626 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1509 ) );
  OAI22_X1 U2768 ( .A1(n989), .A2(n764), .B1(\unit_decode/RegisterFile/n3627 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1508 ) );
  OAI22_X1 U2769 ( .A1(n989), .A2(n767), .B1(\unit_decode/RegisterFile/n3628 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1507 ) );
  OAI22_X1 U2770 ( .A1(n989), .A2(n770), .B1(\unit_decode/RegisterFile/n3629 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1506 ) );
  OAI22_X1 U2771 ( .A1(n989), .A2(n773), .B1(\unit_decode/RegisterFile/n3630 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1505 ) );
  OAI22_X1 U2772 ( .A1(n989), .A2(n776), .B1(\unit_decode/RegisterFile/n3631 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1504 ) );
  OAI22_X1 U2773 ( .A1(n990), .A2(n779), .B1(\unit_decode/RegisterFile/n3632 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1503 ) );
  OAI22_X1 U2774 ( .A1(n990), .A2(n782), .B1(\unit_decode/RegisterFile/n3633 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1502 ) );
  OAI22_X1 U2775 ( .A1(n990), .A2(n785), .B1(\unit_decode/RegisterFile/n3634 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1501 ) );
  OAI22_X1 U2776 ( .A1(n990), .A2(n788), .B1(\unit_decode/RegisterFile/n3635 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1500 ) );
  OAI22_X1 U2777 ( .A1(n990), .A2(n791), .B1(\unit_decode/RegisterFile/n3636 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1499 ) );
  OAI22_X1 U2778 ( .A1(n991), .A2(n794), .B1(\unit_decode/RegisterFile/n3637 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1498 ) );
  OAI22_X1 U2779 ( .A1(n991), .A2(n797), .B1(\unit_decode/RegisterFile/n3638 ), 
        .B2(\unit_decode/n2259 ), .ZN(\unit_decode/RegisterFile/n1497 ) );
  OAI22_X1 U2780 ( .A1(n991), .A2(n800), .B1(\unit_decode/RegisterFile/n3639 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1496 ) );
  OAI22_X1 U2781 ( .A1(n991), .A2(n803), .B1(\unit_decode/RegisterFile/n3640 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1495 ) );
  OAI22_X1 U2782 ( .A1(n991), .A2(n806), .B1(\unit_decode/RegisterFile/n3641 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1494 ) );
  OAI22_X1 U2783 ( .A1(n992), .A2(n809), .B1(\unit_decode/RegisterFile/n3642 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1493 ) );
  OAI22_X1 U2784 ( .A1(n992), .A2(n812), .B1(\unit_decode/RegisterFile/n3643 ), 
        .B2(n985), .ZN(\unit_decode/RegisterFile/n1492 ) );
  OAI22_X1 U2785 ( .A1(n978), .A2(n743), .B1(\unit_decode/RegisterFile/n3588 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1547 ) );
  OAI22_X1 U2786 ( .A1(n978), .A2(n746), .B1(\unit_decode/RegisterFile/n3589 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1546 ) );
  OAI22_X1 U2787 ( .A1(n979), .A2(n749), .B1(\unit_decode/RegisterFile/n3590 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1545 ) );
  OAI22_X1 U2788 ( .A1(n979), .A2(n752), .B1(\unit_decode/RegisterFile/n3591 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1544 ) );
  OAI22_X1 U2789 ( .A1(n979), .A2(n755), .B1(\unit_decode/RegisterFile/n3592 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1543 ) );
  OAI22_X1 U2790 ( .A1(n979), .A2(n758), .B1(\unit_decode/RegisterFile/n3593 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1542 ) );
  OAI22_X1 U2791 ( .A1(n979), .A2(n761), .B1(\unit_decode/RegisterFile/n3594 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1541 ) );
  OAI22_X1 U2792 ( .A1(n980), .A2(n764), .B1(\unit_decode/RegisterFile/n3595 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1540 ) );
  OAI22_X1 U2793 ( .A1(n980), .A2(n767), .B1(\unit_decode/RegisterFile/n3596 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1539 ) );
  OAI22_X1 U2794 ( .A1(n980), .A2(n770), .B1(\unit_decode/RegisterFile/n3597 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1538 ) );
  OAI22_X1 U2795 ( .A1(n980), .A2(n773), .B1(\unit_decode/RegisterFile/n3598 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1537 ) );
  OAI22_X1 U2796 ( .A1(n980), .A2(n776), .B1(\unit_decode/RegisterFile/n3599 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1536 ) );
  OAI22_X1 U2797 ( .A1(n981), .A2(n779), .B1(\unit_decode/RegisterFile/n3600 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1535 ) );
  OAI22_X1 U2798 ( .A1(n981), .A2(n782), .B1(\unit_decode/RegisterFile/n3601 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1534 ) );
  OAI22_X1 U2799 ( .A1(n981), .A2(n785), .B1(\unit_decode/RegisterFile/n3602 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1533 ) );
  OAI22_X1 U2800 ( .A1(n981), .A2(n788), .B1(\unit_decode/RegisterFile/n3603 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1532 ) );
  OAI22_X1 U2801 ( .A1(n981), .A2(n791), .B1(\unit_decode/RegisterFile/n3604 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1531 ) );
  OAI22_X1 U2802 ( .A1(n982), .A2(n794), .B1(\unit_decode/RegisterFile/n3605 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1530 ) );
  OAI22_X1 U2803 ( .A1(n982), .A2(n797), .B1(\unit_decode/RegisterFile/n3606 ), 
        .B2(\unit_decode/n2258 ), .ZN(\unit_decode/RegisterFile/n1529 ) );
  OAI22_X1 U2804 ( .A1(n982), .A2(n800), .B1(\unit_decode/RegisterFile/n3607 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1528 ) );
  OAI22_X1 U2805 ( .A1(n982), .A2(n803), .B1(\unit_decode/RegisterFile/n3608 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1527 ) );
  OAI22_X1 U2806 ( .A1(n982), .A2(n806), .B1(\unit_decode/RegisterFile/n3609 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1526 ) );
  OAI22_X1 U2807 ( .A1(n983), .A2(n809), .B1(\unit_decode/RegisterFile/n3610 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1525 ) );
  OAI22_X1 U2808 ( .A1(n983), .A2(n812), .B1(\unit_decode/RegisterFile/n3611 ), 
        .B2(n976), .ZN(\unit_decode/RegisterFile/n1524 ) );
  OAI22_X1 U2809 ( .A1(n951), .A2(n746), .B1(\unit_decode/RegisterFile/n3493 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1642 ) );
  OAI22_X1 U2810 ( .A1(n952), .A2(n749), .B1(\unit_decode/RegisterFile/n3494 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1641 ) );
  OAI22_X1 U2811 ( .A1(n952), .A2(n752), .B1(\unit_decode/RegisterFile/n3495 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1640 ) );
  OAI22_X1 U2812 ( .A1(n952), .A2(n755), .B1(\unit_decode/RegisterFile/n3496 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1639 ) );
  OAI22_X1 U2813 ( .A1(n952), .A2(n758), .B1(\unit_decode/RegisterFile/n3497 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1638 ) );
  OAI22_X1 U2814 ( .A1(n952), .A2(n761), .B1(\unit_decode/RegisterFile/n3498 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1637 ) );
  OAI22_X1 U2815 ( .A1(n953), .A2(n764), .B1(\unit_decode/RegisterFile/n3499 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1636 ) );
  OAI22_X1 U2816 ( .A1(n953), .A2(n767), .B1(\unit_decode/RegisterFile/n3500 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1635 ) );
  OAI22_X1 U2817 ( .A1(n953), .A2(n770), .B1(\unit_decode/RegisterFile/n3501 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1634 ) );
  OAI22_X1 U2818 ( .A1(n953), .A2(n773), .B1(\unit_decode/RegisterFile/n3502 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1633 ) );
  OAI22_X1 U2819 ( .A1(n953), .A2(n776), .B1(\unit_decode/RegisterFile/n3503 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1632 ) );
  OAI22_X1 U2820 ( .A1(n954), .A2(n779), .B1(\unit_decode/RegisterFile/n3504 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1631 ) );
  OAI22_X1 U2821 ( .A1(n954), .A2(n782), .B1(\unit_decode/RegisterFile/n3505 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1630 ) );
  OAI22_X1 U2822 ( .A1(n954), .A2(n785), .B1(\unit_decode/RegisterFile/n3506 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1629 ) );
  OAI22_X1 U2823 ( .A1(n954), .A2(n788), .B1(\unit_decode/RegisterFile/n3507 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1628 ) );
  OAI22_X1 U2824 ( .A1(n954), .A2(n791), .B1(\unit_decode/RegisterFile/n3508 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1627 ) );
  OAI22_X1 U2825 ( .A1(n955), .A2(n794), .B1(\unit_decode/RegisterFile/n3509 ), 
        .B2(\unit_decode/n2254 ), .ZN(\unit_decode/RegisterFile/n1626 ) );
  OAI22_X1 U2826 ( .A1(n955), .A2(n797), .B1(\unit_decode/RegisterFile/n3510 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1625 ) );
  OAI22_X1 U2827 ( .A1(n955), .A2(n800), .B1(\unit_decode/RegisterFile/n3511 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1624 ) );
  OAI22_X1 U2828 ( .A1(n956), .A2(n809), .B1(\unit_decode/RegisterFile/n3514 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1621 ) );
  OAI22_X1 U2829 ( .A1(n956), .A2(n812), .B1(\unit_decode/RegisterFile/n3515 ), 
        .B2(n949), .ZN(\unit_decode/RegisterFile/n1620 ) );
  OAI22_X1 U2830 ( .A1(n1049), .A2(n711), .B1(\unit_decode/RegisterFile/n3836 ), .B2(n1048), .ZN(\unit_decode/RegisterFile/n1299 ) );
  OAI22_X1 U2831 ( .A1(n1049), .A2(n723), .B1(\unit_decode/RegisterFile/n3837 ), .B2(n1048), .ZN(\unit_decode/RegisterFile/n1298 ) );
  OAI22_X1 U2832 ( .A1(n1049), .A2(n726), .B1(\unit_decode/RegisterFile/n3838 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1297 ) );
  OAI22_X1 U2833 ( .A1(n1049), .A2(n729), .B1(\unit_decode/RegisterFile/n3839 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1296 ) );
  OAI22_X1 U2834 ( .A1(n1049), .A2(n732), .B1(\unit_decode/RegisterFile/n3840 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1295 ) );
  OAI22_X1 U2835 ( .A1(n1050), .A2(n735), .B1(\unit_decode/RegisterFile/n3841 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1294 ) );
  OAI22_X1 U2836 ( .A1(n1050), .A2(n738), .B1(\unit_decode/RegisterFile/n3842 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1293 ) );
  OAI22_X1 U2837 ( .A1(n1050), .A2(n741), .B1(\unit_decode/RegisterFile/n3843 ), .B2(\unit_decode/n2267 ), .ZN(\unit_decode/RegisterFile/n1292 ) );
  OAI22_X1 U2838 ( .A1(n1031), .A2(n711), .B1(\unit_decode/RegisterFile/n3772 ), .B2(n1030), .ZN(\unit_decode/RegisterFile/n1363 ) );
  OAI22_X1 U2839 ( .A1(n1031), .A2(n723), .B1(\unit_decode/RegisterFile/n3773 ), .B2(n1030), .ZN(\unit_decode/RegisterFile/n1362 ) );
  OAI22_X1 U2840 ( .A1(n1031), .A2(n726), .B1(\unit_decode/RegisterFile/n3774 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1361 ) );
  OAI22_X1 U2841 ( .A1(n1031), .A2(n729), .B1(\unit_decode/RegisterFile/n3775 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1360 ) );
  OAI22_X1 U2842 ( .A1(n1031), .A2(n732), .B1(\unit_decode/RegisterFile/n3776 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1359 ) );
  OAI22_X1 U2843 ( .A1(n1032), .A2(n735), .B1(\unit_decode/RegisterFile/n3777 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1358 ) );
  OAI22_X1 U2844 ( .A1(n1032), .A2(n738), .B1(\unit_decode/RegisterFile/n3778 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1357 ) );
  OAI22_X1 U2845 ( .A1(n1032), .A2(n741), .B1(\unit_decode/RegisterFile/n3779 ), .B2(\unit_decode/n2265 ), .ZN(\unit_decode/RegisterFile/n1356 ) );
  OAI22_X1 U2846 ( .A1(n1022), .A2(n711), .B1(\unit_decode/RegisterFile/n3740 ), .B2(n1021), .ZN(\unit_decode/RegisterFile/n1395 ) );
  OAI22_X1 U2847 ( .A1(n1022), .A2(n723), .B1(\unit_decode/RegisterFile/n3741 ), .B2(n1021), .ZN(\unit_decode/RegisterFile/n1394 ) );
  OAI22_X1 U2848 ( .A1(n1022), .A2(n726), .B1(\unit_decode/RegisterFile/n3742 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1393 ) );
  OAI22_X1 U2849 ( .A1(n1022), .A2(n729), .B1(\unit_decode/RegisterFile/n3743 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1392 ) );
  OAI22_X1 U2850 ( .A1(n1022), .A2(n732), .B1(\unit_decode/RegisterFile/n3744 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1391 ) );
  OAI22_X1 U2851 ( .A1(n1023), .A2(n735), .B1(\unit_decode/RegisterFile/n3745 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1390 ) );
  OAI22_X1 U2852 ( .A1(n1023), .A2(n738), .B1(\unit_decode/RegisterFile/n3746 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1389 ) );
  OAI22_X1 U2853 ( .A1(n1023), .A2(n741), .B1(\unit_decode/RegisterFile/n3747 ), .B2(\unit_decode/n2263 ), .ZN(\unit_decode/RegisterFile/n1388 ) );
  OAI22_X1 U2854 ( .A1(n959), .A2(n710), .B1(\unit_decode/RegisterFile/n3516 ), 
        .B2(n958), .ZN(\unit_decode/RegisterFile/n1619 ) );
  OAI22_X1 U2855 ( .A1(n959), .A2(n722), .B1(\unit_decode/RegisterFile/n3517 ), 
        .B2(n958), .ZN(\unit_decode/RegisterFile/n1618 ) );
  OAI22_X1 U2856 ( .A1(n959), .A2(n725), .B1(\unit_decode/RegisterFile/n3518 ), 
        .B2(\unit_decode/n2256 ), .ZN(\unit_decode/RegisterFile/n1617 ) );
  OAI22_X1 U2857 ( .A1(n251), .A2(n359), .B1(\unit_memory/DRAM/n2399 ), .B2(
        n361), .ZN(\unit_memory/DRAM/n2148 ) );
  OAI22_X1 U2858 ( .A1(n266), .A2(n360), .B1(\unit_memory/DRAM/n2400 ), .B2(
        n361), .ZN(\unit_memory/DRAM/n2147 ) );
  OAI22_X1 U2859 ( .A1(n269), .A2(n359), .B1(\unit_memory/DRAM/n2401 ), .B2(
        n361), .ZN(\unit_memory/DRAM/n2146 ) );
  OAI22_X1 U2860 ( .A1(n272), .A2(n360), .B1(\unit_memory/DRAM/n2402 ), .B2(
        n361), .ZN(\unit_memory/DRAM/n2145 ) );
  OAI22_X1 U2861 ( .A1(n275), .A2(n359), .B1(\unit_memory/DRAM/n2403 ), .B2(
        n362), .ZN(\unit_memory/DRAM/n2144 ) );
  OAI22_X1 U2862 ( .A1(n278), .A2(n360), .B1(\unit_memory/DRAM/n2404 ), .B2(
        n362), .ZN(\unit_memory/DRAM/n2143 ) );
  OAI22_X1 U2863 ( .A1(n281), .A2(n359), .B1(\unit_memory/DRAM/n2405 ), .B2(
        n362), .ZN(\unit_memory/DRAM/n2142 ) );
  OAI22_X1 U2864 ( .A1(n284), .A2(n360), .B1(\unit_memory/DRAM/n2406 ), .B2(
        n362), .ZN(\unit_memory/DRAM/n2141 ) );
  OAI22_X1 U2865 ( .A1(n287), .A2(n360), .B1(\unit_memory/DRAM/n2407 ), .B2(
        n363), .ZN(\unit_memory/DRAM/n2140 ) );
  OAI22_X1 U2866 ( .A1(n290), .A2(n360), .B1(\unit_memory/DRAM/n2408 ), .B2(
        n363), .ZN(\unit_memory/DRAM/n2139 ) );
  OAI22_X1 U2867 ( .A1(n293), .A2(n360), .B1(\unit_memory/DRAM/n2409 ), .B2(
        n363), .ZN(\unit_memory/DRAM/n2138 ) );
  OAI22_X1 U2868 ( .A1(n296), .A2(n360), .B1(\unit_memory/DRAM/n2410 ), .B2(
        n363), .ZN(\unit_memory/DRAM/n2137 ) );
  OAI22_X1 U2869 ( .A1(n299), .A2(n360), .B1(\unit_memory/DRAM/n2411 ), .B2(
        n364), .ZN(\unit_memory/DRAM/n2136 ) );
  OAI22_X1 U2870 ( .A1(n302), .A2(n360), .B1(\unit_memory/DRAM/n2412 ), .B2(
        n364), .ZN(\unit_memory/DRAM/n2135 ) );
  OAI22_X1 U2871 ( .A1(n305), .A2(n360), .B1(\unit_memory/DRAM/n2413 ), .B2(
        n364), .ZN(\unit_memory/DRAM/n2134 ) );
  OAI22_X1 U2872 ( .A1(n308), .A2(n360), .B1(\unit_memory/DRAM/n2414 ), .B2(
        n364), .ZN(\unit_memory/DRAM/n2133 ) );
  OAI22_X1 U2873 ( .A1(n311), .A2(n360), .B1(\unit_memory/DRAM/n2415 ), .B2(
        n365), .ZN(\unit_memory/DRAM/n2132 ) );
  OAI22_X1 U2874 ( .A1(n335), .A2(n359), .B1(\unit_memory/DRAM/n2423 ), .B2(
        n367), .ZN(\unit_memory/DRAM/n2124 ) );
  OAI22_X1 U2875 ( .A1(n251), .A2(n403), .B1(\unit_memory/DRAM/n2527 ), .B2(
        n405), .ZN(\unit_memory/DRAM/n2020 ) );
  OAI22_X1 U2876 ( .A1(n266), .A2(n404), .B1(\unit_memory/DRAM/n2528 ), .B2(
        n405), .ZN(\unit_memory/DRAM/n2019 ) );
  OAI22_X1 U2877 ( .A1(n269), .A2(n403), .B1(\unit_memory/DRAM/n2529 ), .B2(
        n405), .ZN(\unit_memory/DRAM/n2018 ) );
  OAI22_X1 U2878 ( .A1(n272), .A2(n404), .B1(\unit_memory/DRAM/n2530 ), .B2(
        n405), .ZN(\unit_memory/DRAM/n2017 ) );
  OAI22_X1 U2879 ( .A1(n275), .A2(n403), .B1(\unit_memory/DRAM/n2531 ), .B2(
        n406), .ZN(\unit_memory/DRAM/n2016 ) );
  OAI22_X1 U2880 ( .A1(n278), .A2(n404), .B1(\unit_memory/DRAM/n2532 ), .B2(
        n406), .ZN(\unit_memory/DRAM/n2015 ) );
  OAI22_X1 U2881 ( .A1(n281), .A2(n403), .B1(\unit_memory/DRAM/n2533 ), .B2(
        n406), .ZN(\unit_memory/DRAM/n2014 ) );
  OAI22_X1 U2882 ( .A1(n284), .A2(n404), .B1(\unit_memory/DRAM/n2534 ), .B2(
        n406), .ZN(\unit_memory/DRAM/n2013 ) );
  OAI22_X1 U2883 ( .A1(n287), .A2(n404), .B1(\unit_memory/DRAM/n2535 ), .B2(
        n407), .ZN(\unit_memory/DRAM/n2012 ) );
  OAI22_X1 U2884 ( .A1(n290), .A2(n404), .B1(\unit_memory/DRAM/n2536 ), .B2(
        n407), .ZN(\unit_memory/DRAM/n2011 ) );
  OAI22_X1 U2885 ( .A1(n293), .A2(n404), .B1(\unit_memory/DRAM/n2537 ), .B2(
        n407), .ZN(\unit_memory/DRAM/n2010 ) );
  OAI22_X1 U2886 ( .A1(n296), .A2(n404), .B1(\unit_memory/DRAM/n2538 ), .B2(
        n407), .ZN(\unit_memory/DRAM/n2009 ) );
  OAI22_X1 U2887 ( .A1(n299), .A2(n404), .B1(\unit_memory/DRAM/n2539 ), .B2(
        n408), .ZN(\unit_memory/DRAM/n2008 ) );
  OAI22_X1 U2888 ( .A1(n302), .A2(n404), .B1(\unit_memory/DRAM/n2540 ), .B2(
        n408), .ZN(\unit_memory/DRAM/n2007 ) );
  OAI22_X1 U2889 ( .A1(n305), .A2(n404), .B1(\unit_memory/DRAM/n2541 ), .B2(
        n408), .ZN(\unit_memory/DRAM/n2006 ) );
  OAI22_X1 U2890 ( .A1(n308), .A2(n404), .B1(\unit_memory/DRAM/n2542 ), .B2(
        n408), .ZN(\unit_memory/DRAM/n2005 ) );
  OAI22_X1 U2891 ( .A1(n311), .A2(n404), .B1(\unit_memory/DRAM/n2543 ), .B2(
        n409), .ZN(\unit_memory/DRAM/n2004 ) );
  OAI22_X1 U2892 ( .A1(n335), .A2(n403), .B1(\unit_memory/DRAM/n2551 ), .B2(
        n411), .ZN(\unit_memory/DRAM/n1996 ) );
  OAI22_X1 U2893 ( .A1(n259), .A2(n287), .B1(\unit_memory/DRAM/n2375 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2172 ) );
  OAI22_X1 U2894 ( .A1(n259), .A2(n290), .B1(\unit_memory/DRAM/n2376 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2171 ) );
  OAI22_X1 U2895 ( .A1(n259), .A2(n293), .B1(\unit_memory/DRAM/n2377 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2170 ) );
  OAI22_X1 U2896 ( .A1(n259), .A2(n296), .B1(\unit_memory/DRAM/n2378 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2169 ) );
  OAI22_X1 U2897 ( .A1(n260), .A2(n299), .B1(\unit_memory/DRAM/n2379 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2168 ) );
  OAI22_X1 U2898 ( .A1(n260), .A2(n302), .B1(\unit_memory/DRAM/n2380 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2167 ) );
  OAI22_X1 U2899 ( .A1(n260), .A2(n305), .B1(\unit_memory/DRAM/n2381 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2166 ) );
  OAI22_X1 U2900 ( .A1(n260), .A2(n308), .B1(\unit_memory/DRAM/n2382 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2165 ) );
  OAI22_X1 U2901 ( .A1(n261), .A2(n311), .B1(\unit_memory/DRAM/n2383 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2164 ) );
  OAI22_X1 U2902 ( .A1(n263), .A2(n335), .B1(\unit_memory/DRAM/n2391 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2156 ) );
  OAI22_X1 U2903 ( .A1(n251), .A2(n370), .B1(\unit_memory/DRAM/n2431 ), .B2(
        n372), .ZN(\unit_memory/DRAM/n2116 ) );
  OAI22_X1 U2904 ( .A1(n266), .A2(n371), .B1(\unit_memory/DRAM/n2432 ), .B2(
        n372), .ZN(\unit_memory/DRAM/n2115 ) );
  OAI22_X1 U2905 ( .A1(n269), .A2(n370), .B1(\unit_memory/DRAM/n2433 ), .B2(
        n372), .ZN(\unit_memory/DRAM/n2114 ) );
  OAI22_X1 U2906 ( .A1(n272), .A2(n371), .B1(\unit_memory/DRAM/n2434 ), .B2(
        n372), .ZN(\unit_memory/DRAM/n2113 ) );
  OAI22_X1 U2907 ( .A1(n275), .A2(n370), .B1(\unit_memory/DRAM/n2435 ), .B2(
        n373), .ZN(\unit_memory/DRAM/n2112 ) );
  OAI22_X1 U2908 ( .A1(n278), .A2(n371), .B1(\unit_memory/DRAM/n2436 ), .B2(
        n373), .ZN(\unit_memory/DRAM/n2111 ) );
  OAI22_X1 U2909 ( .A1(n281), .A2(n370), .B1(\unit_memory/DRAM/n2437 ), .B2(
        n373), .ZN(\unit_memory/DRAM/n2110 ) );
  OAI22_X1 U2910 ( .A1(n284), .A2(n371), .B1(\unit_memory/DRAM/n2438 ), .B2(
        n373), .ZN(\unit_memory/DRAM/n2109 ) );
  OAI22_X1 U2911 ( .A1(n287), .A2(n371), .B1(\unit_memory/DRAM/n2439 ), .B2(
        n374), .ZN(\unit_memory/DRAM/n2108 ) );
  OAI22_X1 U2912 ( .A1(n290), .A2(n371), .B1(\unit_memory/DRAM/n2440 ), .B2(
        n374), .ZN(\unit_memory/DRAM/n2107 ) );
  OAI22_X1 U2913 ( .A1(n293), .A2(n371), .B1(\unit_memory/DRAM/n2441 ), .B2(
        n374), .ZN(\unit_memory/DRAM/n2106 ) );
  OAI22_X1 U2914 ( .A1(n296), .A2(n371), .B1(\unit_memory/DRAM/n2442 ), .B2(
        n374), .ZN(\unit_memory/DRAM/n2105 ) );
  OAI22_X1 U2915 ( .A1(n299), .A2(n371), .B1(\unit_memory/DRAM/n2443 ), .B2(
        n375), .ZN(\unit_memory/DRAM/n2104 ) );
  OAI22_X1 U2916 ( .A1(n302), .A2(n371), .B1(\unit_memory/DRAM/n2444 ), .B2(
        n375), .ZN(\unit_memory/DRAM/n2103 ) );
  OAI22_X1 U2917 ( .A1(n305), .A2(n371), .B1(\unit_memory/DRAM/n2445 ), .B2(
        n375), .ZN(\unit_memory/DRAM/n2102 ) );
  OAI22_X1 U2918 ( .A1(n308), .A2(n371), .B1(\unit_memory/DRAM/n2446 ), .B2(
        n375), .ZN(\unit_memory/DRAM/n2101 ) );
  OAI22_X1 U2919 ( .A1(n311), .A2(n371), .B1(\unit_memory/DRAM/n2447 ), .B2(
        n376), .ZN(\unit_memory/DRAM/n2100 ) );
  OAI22_X1 U2920 ( .A1(n335), .A2(n370), .B1(\unit_memory/DRAM/n2455 ), .B2(
        n378), .ZN(\unit_memory/DRAM/n2092 ) );
  OAI22_X1 U2921 ( .A1(n311), .A2(n382), .B1(\unit_memory/DRAM/n2479 ), .B2(
        n387), .ZN(\unit_memory/DRAM/n2068 ) );
  OAI22_X1 U2922 ( .A1(n335), .A2(n381), .B1(\unit_memory/DRAM/n2487 ), .B2(
        n389), .ZN(\unit_memory/DRAM/n2060 ) );
  OAI22_X1 U2923 ( .A1(n251), .A2(n392), .B1(\unit_memory/DRAM/n2495 ), .B2(
        n394), .ZN(\unit_memory/DRAM/n2052 ) );
  OAI22_X1 U2924 ( .A1(n266), .A2(n393), .B1(\unit_memory/DRAM/n2496 ), .B2(
        n394), .ZN(\unit_memory/DRAM/n2051 ) );
  OAI22_X1 U2925 ( .A1(n269), .A2(n392), .B1(\unit_memory/DRAM/n2497 ), .B2(
        n394), .ZN(\unit_memory/DRAM/n2050 ) );
  OAI22_X1 U2926 ( .A1(n272), .A2(n393), .B1(\unit_memory/DRAM/n2498 ), .B2(
        n394), .ZN(\unit_memory/DRAM/n2049 ) );
  OAI22_X1 U2927 ( .A1(n275), .A2(n392), .B1(\unit_memory/DRAM/n2499 ), .B2(
        n395), .ZN(\unit_memory/DRAM/n2048 ) );
  OAI22_X1 U2928 ( .A1(n278), .A2(n393), .B1(\unit_memory/DRAM/n2500 ), .B2(
        n395), .ZN(\unit_memory/DRAM/n2047 ) );
  OAI22_X1 U2929 ( .A1(n281), .A2(n392), .B1(\unit_memory/DRAM/n2501 ), .B2(
        n395), .ZN(\unit_memory/DRAM/n2046 ) );
  OAI22_X1 U2930 ( .A1(n284), .A2(n393), .B1(\unit_memory/DRAM/n2502 ), .B2(
        n395), .ZN(\unit_memory/DRAM/n2045 ) );
  OAI22_X1 U2931 ( .A1(n287), .A2(n393), .B1(\unit_memory/DRAM/n2503 ), .B2(
        n396), .ZN(\unit_memory/DRAM/n2044 ) );
  OAI22_X1 U2932 ( .A1(n290), .A2(n393), .B1(\unit_memory/DRAM/n2504 ), .B2(
        n396), .ZN(\unit_memory/DRAM/n2043 ) );
  OAI22_X1 U2933 ( .A1(n293), .A2(n393), .B1(\unit_memory/DRAM/n2505 ), .B2(
        n396), .ZN(\unit_memory/DRAM/n2042 ) );
  OAI22_X1 U2934 ( .A1(n296), .A2(n393), .B1(\unit_memory/DRAM/n2506 ), .B2(
        n396), .ZN(\unit_memory/DRAM/n2041 ) );
  OAI22_X1 U2935 ( .A1(n299), .A2(n393), .B1(\unit_memory/DRAM/n2507 ), .B2(
        n397), .ZN(\unit_memory/DRAM/n2040 ) );
  OAI22_X1 U2936 ( .A1(n302), .A2(n393), .B1(\unit_memory/DRAM/n2508 ), .B2(
        n397), .ZN(\unit_memory/DRAM/n2039 ) );
  OAI22_X1 U2937 ( .A1(n305), .A2(n393), .B1(\unit_memory/DRAM/n2509 ), .B2(
        n397), .ZN(\unit_memory/DRAM/n2038 ) );
  OAI22_X1 U2938 ( .A1(n308), .A2(n393), .B1(\unit_memory/DRAM/n2510 ), .B2(
        n397), .ZN(\unit_memory/DRAM/n2037 ) );
  OAI22_X1 U2939 ( .A1(n311), .A2(n393), .B1(\unit_memory/DRAM/n2511 ), .B2(
        n398), .ZN(\unit_memory/DRAM/n2036 ) );
  OAI22_X1 U2940 ( .A1(n335), .A2(n392), .B1(\unit_memory/DRAM/n2519 ), .B2(
        n400), .ZN(\unit_memory/DRAM/n2028 ) );
  OAI22_X1 U2941 ( .A1(n251), .A2(n414), .B1(\unit_memory/DRAM/n2559 ), .B2(
        n416), .ZN(\unit_memory/DRAM/n1988 ) );
  OAI22_X1 U2942 ( .A1(n266), .A2(n415), .B1(\unit_memory/DRAM/n2560 ), .B2(
        n416), .ZN(\unit_memory/DRAM/n1987 ) );
  OAI22_X1 U2943 ( .A1(n269), .A2(n414), .B1(\unit_memory/DRAM/n2561 ), .B2(
        n416), .ZN(\unit_memory/DRAM/n1986 ) );
  OAI22_X1 U2944 ( .A1(n272), .A2(n415), .B1(\unit_memory/DRAM/n2562 ), .B2(
        n416), .ZN(\unit_memory/DRAM/n1985 ) );
  OAI22_X1 U2945 ( .A1(n275), .A2(n414), .B1(\unit_memory/DRAM/n2563 ), .B2(
        n417), .ZN(\unit_memory/DRAM/n1984 ) );
  OAI22_X1 U2946 ( .A1(n278), .A2(n415), .B1(\unit_memory/DRAM/n2564 ), .B2(
        n417), .ZN(\unit_memory/DRAM/n1983 ) );
  OAI22_X1 U2947 ( .A1(n281), .A2(n414), .B1(\unit_memory/DRAM/n2565 ), .B2(
        n417), .ZN(\unit_memory/DRAM/n1982 ) );
  OAI22_X1 U2948 ( .A1(n284), .A2(n415), .B1(\unit_memory/DRAM/n2566 ), .B2(
        n417), .ZN(\unit_memory/DRAM/n1981 ) );
  OAI22_X1 U2949 ( .A1(n287), .A2(n415), .B1(\unit_memory/DRAM/n2567 ), .B2(
        n418), .ZN(\unit_memory/DRAM/n1980 ) );
  OAI22_X1 U2950 ( .A1(n290), .A2(n415), .B1(\unit_memory/DRAM/n2568 ), .B2(
        n418), .ZN(\unit_memory/DRAM/n1979 ) );
  OAI22_X1 U2951 ( .A1(n293), .A2(n415), .B1(\unit_memory/DRAM/n2569 ), .B2(
        n418), .ZN(\unit_memory/DRAM/n1978 ) );
  OAI22_X1 U2952 ( .A1(n296), .A2(n415), .B1(\unit_memory/DRAM/n2570 ), .B2(
        n418), .ZN(\unit_memory/DRAM/n1977 ) );
  OAI22_X1 U2953 ( .A1(n299), .A2(n415), .B1(\unit_memory/DRAM/n2571 ), .B2(
        n419), .ZN(\unit_memory/DRAM/n1976 ) );
  OAI22_X1 U2954 ( .A1(n302), .A2(n415), .B1(\unit_memory/DRAM/n2572 ), .B2(
        n419), .ZN(\unit_memory/DRAM/n1975 ) );
  OAI22_X1 U2955 ( .A1(n305), .A2(n415), .B1(\unit_memory/DRAM/n2573 ), .B2(
        n419), .ZN(\unit_memory/DRAM/n1974 ) );
  OAI22_X1 U2956 ( .A1(n308), .A2(n415), .B1(\unit_memory/DRAM/n2574 ), .B2(
        n419), .ZN(\unit_memory/DRAM/n1973 ) );
  OAI22_X1 U2957 ( .A1(n311), .A2(n415), .B1(\unit_memory/DRAM/n2575 ), .B2(
        n420), .ZN(\unit_memory/DRAM/n1972 ) );
  OAI22_X1 U2958 ( .A1(n335), .A2(n414), .B1(\unit_memory/DRAM/n2583 ), .B2(
        n422), .ZN(\unit_memory/DRAM/n1964 ) );
  OAI22_X1 U2959 ( .A1(n311), .A2(n426), .B1(\unit_memory/DRAM/n2607 ), .B2(
        n431), .ZN(\unit_memory/DRAM/n1940 ) );
  OAI22_X1 U2960 ( .A1(n335), .A2(n425), .B1(\unit_memory/DRAM/n2615 ), .B2(
        n433), .ZN(\unit_memory/DRAM/n1932 ) );
  OAI22_X1 U2961 ( .A1(n250), .A2(n525), .B1(\unit_memory/DRAM/n2879 ), .B2(
        n526), .ZN(\unit_memory/DRAM/n1668 ) );
  OAI22_X1 U2962 ( .A1(n267), .A2(n524), .B1(\unit_memory/DRAM/n2880 ), .B2(
        n526), .ZN(\unit_memory/DRAM/n1667 ) );
  OAI22_X1 U2963 ( .A1(n270), .A2(n525), .B1(\unit_memory/DRAM/n2881 ), .B2(
        n526), .ZN(\unit_memory/DRAM/n1666 ) );
  OAI22_X1 U2964 ( .A1(n273), .A2(n524), .B1(\unit_memory/DRAM/n2882 ), .B2(
        n526), .ZN(\unit_memory/DRAM/n1665 ) );
  OAI22_X1 U2965 ( .A1(n276), .A2(n525), .B1(\unit_memory/DRAM/n2883 ), .B2(
        n527), .ZN(\unit_memory/DRAM/n1664 ) );
  OAI22_X1 U2966 ( .A1(n279), .A2(n524), .B1(\unit_memory/DRAM/n2884 ), .B2(
        n527), .ZN(\unit_memory/DRAM/n1663 ) );
  OAI22_X1 U2967 ( .A1(n282), .A2(n525), .B1(\unit_memory/DRAM/n2885 ), .B2(
        n527), .ZN(\unit_memory/DRAM/n1662 ) );
  OAI22_X1 U2968 ( .A1(n285), .A2(n524), .B1(\unit_memory/DRAM/n2886 ), .B2(
        n527), .ZN(\unit_memory/DRAM/n1661 ) );
  OAI22_X1 U2969 ( .A1(n250), .A2(n536), .B1(\unit_memory/DRAM/n2911 ), .B2(
        n537), .ZN(\unit_memory/DRAM/n1636 ) );
  OAI22_X1 U2970 ( .A1(n267), .A2(n535), .B1(\unit_memory/DRAM/n2912 ), .B2(
        n537), .ZN(\unit_memory/DRAM/n1635 ) );
  OAI22_X1 U2971 ( .A1(n270), .A2(n536), .B1(\unit_memory/DRAM/n2913 ), .B2(
        n537), .ZN(\unit_memory/DRAM/n1634 ) );
  OAI22_X1 U2972 ( .A1(n273), .A2(n535), .B1(\unit_memory/DRAM/n2914 ), .B2(
        n537), .ZN(\unit_memory/DRAM/n1633 ) );
  OAI22_X1 U2973 ( .A1(n276), .A2(n536), .B1(\unit_memory/DRAM/n2915 ), .B2(
        n538), .ZN(\unit_memory/DRAM/n1632 ) );
  OAI22_X1 U2974 ( .A1(n279), .A2(n535), .B1(\unit_memory/DRAM/n2916 ), .B2(
        n538), .ZN(\unit_memory/DRAM/n1631 ) );
  OAI22_X1 U2975 ( .A1(n282), .A2(n536), .B1(\unit_memory/DRAM/n2917 ), .B2(
        n538), .ZN(\unit_memory/DRAM/n1630 ) );
  OAI22_X1 U2976 ( .A1(n285), .A2(n535), .B1(\unit_memory/DRAM/n2918 ), .B2(
        n538), .ZN(\unit_memory/DRAM/n1629 ) );
  OAI22_X1 U2977 ( .A1(n288), .A2(n536), .B1(\unit_memory/DRAM/n2919 ), .B2(
        n539), .ZN(\unit_memory/DRAM/n1628 ) );
  OAI22_X1 U2978 ( .A1(n291), .A2(n536), .B1(\unit_memory/DRAM/n2920 ), .B2(
        n539), .ZN(\unit_memory/DRAM/n1627 ) );
  OAI22_X1 U2979 ( .A1(n294), .A2(n536), .B1(\unit_memory/DRAM/n2921 ), .B2(
        n539), .ZN(\unit_memory/DRAM/n1626 ) );
  OAI22_X1 U2980 ( .A1(n297), .A2(n536), .B1(\unit_memory/DRAM/n2922 ), .B2(
        n539), .ZN(\unit_memory/DRAM/n1625 ) );
  OAI22_X1 U2981 ( .A1(n300), .A2(n536), .B1(\unit_memory/DRAM/n2923 ), .B2(
        n540), .ZN(\unit_memory/DRAM/n1624 ) );
  OAI22_X1 U2982 ( .A1(n303), .A2(n536), .B1(\unit_memory/DRAM/n2924 ), .B2(
        n540), .ZN(\unit_memory/DRAM/n1623 ) );
  OAI22_X1 U2983 ( .A1(n306), .A2(n536), .B1(\unit_memory/DRAM/n2925 ), .B2(
        n540), .ZN(\unit_memory/DRAM/n1622 ) );
  OAI22_X1 U2984 ( .A1(n309), .A2(n536), .B1(\unit_memory/DRAM/n2926 ), .B2(
        n540), .ZN(\unit_memory/DRAM/n1621 ) );
  OAI22_X1 U2985 ( .A1(n312), .A2(n536), .B1(\unit_memory/DRAM/n2927 ), .B2(
        n541), .ZN(\unit_memory/DRAM/n1620 ) );
  OAI22_X1 U2986 ( .A1(n315), .A2(n536), .B1(\unit_memory/DRAM/n2928 ), .B2(
        n541), .ZN(\unit_memory/DRAM/n1619 ) );
  OAI22_X1 U2987 ( .A1(n318), .A2(n536), .B1(\unit_memory/DRAM/n2929 ), .B2(
        n541), .ZN(\unit_memory/DRAM/n1618 ) );
  OAI22_X1 U2988 ( .A1(n321), .A2(n536), .B1(\unit_memory/DRAM/n2930 ), .B2(
        n541), .ZN(\unit_memory/DRAM/n1617 ) );
  OAI22_X1 U2989 ( .A1(n324), .A2(n535), .B1(\unit_memory/DRAM/n2931 ), .B2(
        n542), .ZN(\unit_memory/DRAM/n1616 ) );
  OAI22_X1 U2990 ( .A1(n327), .A2(n535), .B1(\unit_memory/DRAM/n2932 ), .B2(
        n542), .ZN(\unit_memory/DRAM/n1615 ) );
  OAI22_X1 U2991 ( .A1(n330), .A2(n535), .B1(\unit_memory/DRAM/n2933 ), .B2(
        n542), .ZN(\unit_memory/DRAM/n1614 ) );
  OAI22_X1 U2992 ( .A1(n333), .A2(n535), .B1(\unit_memory/DRAM/n2934 ), .B2(
        n542), .ZN(\unit_memory/DRAM/n1613 ) );
  OAI22_X1 U2993 ( .A1(n336), .A2(n535), .B1(\unit_memory/DRAM/n2935 ), .B2(
        n543), .ZN(\unit_memory/DRAM/n1612 ) );
  OAI22_X1 U2994 ( .A1(n339), .A2(n535), .B1(\unit_memory/DRAM/n2936 ), .B2(
        n543), .ZN(\unit_memory/DRAM/n1611 ) );
  OAI22_X1 U2995 ( .A1(n342), .A2(n535), .B1(\unit_memory/DRAM/n2937 ), .B2(
        n543), .ZN(\unit_memory/DRAM/n1610 ) );
  OAI22_X1 U2996 ( .A1(n345), .A2(n535), .B1(\unit_memory/DRAM/n2938 ), .B2(
        n543), .ZN(\unit_memory/DRAM/n1609 ) );
  OAI22_X1 U2997 ( .A1(n348), .A2(n535), .B1(\unit_memory/DRAM/n2939 ), .B2(
        n544), .ZN(\unit_memory/DRAM/n1608 ) );
  OAI22_X1 U2998 ( .A1(n351), .A2(n535), .B1(\unit_memory/DRAM/n2940 ), .B2(
        n544), .ZN(\unit_memory/DRAM/n1607 ) );
  OAI22_X1 U2999 ( .A1(n354), .A2(n535), .B1(\unit_memory/DRAM/n2941 ), .B2(
        n544), .ZN(\unit_memory/DRAM/n1606 ) );
  OAI22_X1 U3000 ( .A1(n357), .A2(n535), .B1(\unit_memory/DRAM/n2942 ), .B2(
        n544), .ZN(\unit_memory/DRAM/n1605 ) );
  OAI22_X1 U3001 ( .A1(n249), .A2(n569), .B1(\unit_memory/DRAM/n3007 ), .B2(
        n570), .ZN(\unit_memory/DRAM/n1540 ) );
  OAI22_X1 U3002 ( .A1(n267), .A2(n568), .B1(\unit_memory/DRAM/n3008 ), .B2(
        n570), .ZN(\unit_memory/DRAM/n1539 ) );
  OAI22_X1 U3003 ( .A1(n270), .A2(n569), .B1(\unit_memory/DRAM/n3009 ), .B2(
        n570), .ZN(\unit_memory/DRAM/n1538 ) );
  OAI22_X1 U3004 ( .A1(n273), .A2(n568), .B1(\unit_memory/DRAM/n3010 ), .B2(
        n570), .ZN(\unit_memory/DRAM/n1537 ) );
  OAI22_X1 U3005 ( .A1(n276), .A2(n569), .B1(\unit_memory/DRAM/n3011 ), .B2(
        n571), .ZN(\unit_memory/DRAM/n1536 ) );
  OAI22_X1 U3006 ( .A1(n279), .A2(n568), .B1(\unit_memory/DRAM/n3012 ), .B2(
        n571), .ZN(\unit_memory/DRAM/n1535 ) );
  OAI22_X1 U3007 ( .A1(n282), .A2(n569), .B1(\unit_memory/DRAM/n3013 ), .B2(
        n571), .ZN(\unit_memory/DRAM/n1534 ) );
  OAI22_X1 U3008 ( .A1(n285), .A2(n568), .B1(\unit_memory/DRAM/n3014 ), .B2(
        n571), .ZN(\unit_memory/DRAM/n1533 ) );
  OAI22_X1 U3009 ( .A1(n249), .A2(n580), .B1(\unit_memory/DRAM/n3039 ), .B2(
        n581), .ZN(\unit_memory/DRAM/n1508 ) );
  OAI22_X1 U3010 ( .A1(n267), .A2(n579), .B1(\unit_memory/DRAM/n3040 ), .B2(
        n581), .ZN(\unit_memory/DRAM/n1507 ) );
  OAI22_X1 U3011 ( .A1(n270), .A2(n580), .B1(\unit_memory/DRAM/n3041 ), .B2(
        n581), .ZN(\unit_memory/DRAM/n1506 ) );
  OAI22_X1 U3012 ( .A1(n273), .A2(n579), .B1(\unit_memory/DRAM/n3042 ), .B2(
        n581), .ZN(\unit_memory/DRAM/n1505 ) );
  OAI22_X1 U3013 ( .A1(n276), .A2(n580), .B1(\unit_memory/DRAM/n3043 ), .B2(
        n582), .ZN(\unit_memory/DRAM/n1504 ) );
  OAI22_X1 U3014 ( .A1(n279), .A2(n579), .B1(\unit_memory/DRAM/n3044 ), .B2(
        n582), .ZN(\unit_memory/DRAM/n1503 ) );
  OAI22_X1 U3015 ( .A1(n282), .A2(n580), .B1(\unit_memory/DRAM/n3045 ), .B2(
        n582), .ZN(\unit_memory/DRAM/n1502 ) );
  OAI22_X1 U3016 ( .A1(n285), .A2(n579), .B1(\unit_memory/DRAM/n3046 ), .B2(
        n582), .ZN(\unit_memory/DRAM/n1501 ) );
  OAI22_X1 U3017 ( .A1(n288), .A2(n580), .B1(\unit_memory/DRAM/n3047 ), .B2(
        n583), .ZN(\unit_memory/DRAM/n1500 ) );
  OAI22_X1 U3018 ( .A1(n291), .A2(n580), .B1(\unit_memory/DRAM/n3048 ), .B2(
        n583), .ZN(\unit_memory/DRAM/n1499 ) );
  OAI22_X1 U3019 ( .A1(n294), .A2(n580), .B1(\unit_memory/DRAM/n3049 ), .B2(
        n583), .ZN(\unit_memory/DRAM/n1498 ) );
  OAI22_X1 U3020 ( .A1(n297), .A2(n580), .B1(\unit_memory/DRAM/n3050 ), .B2(
        n583), .ZN(\unit_memory/DRAM/n1497 ) );
  OAI22_X1 U3021 ( .A1(n300), .A2(n580), .B1(\unit_memory/DRAM/n3051 ), .B2(
        n584), .ZN(\unit_memory/DRAM/n1496 ) );
  OAI22_X1 U3022 ( .A1(n303), .A2(n580), .B1(\unit_memory/DRAM/n3052 ), .B2(
        n584), .ZN(\unit_memory/DRAM/n1495 ) );
  OAI22_X1 U3023 ( .A1(n306), .A2(n580), .B1(\unit_memory/DRAM/n3053 ), .B2(
        n584), .ZN(\unit_memory/DRAM/n1494 ) );
  OAI22_X1 U3024 ( .A1(n309), .A2(n580), .B1(\unit_memory/DRAM/n3054 ), .B2(
        n584), .ZN(\unit_memory/DRAM/n1493 ) );
  OAI22_X1 U3025 ( .A1(n312), .A2(n580), .B1(\unit_memory/DRAM/n3055 ), .B2(
        n585), .ZN(\unit_memory/DRAM/n1492 ) );
  OAI22_X1 U3026 ( .A1(n315), .A2(n580), .B1(\unit_memory/DRAM/n3056 ), .B2(
        n585), .ZN(\unit_memory/DRAM/n1491 ) );
  OAI22_X1 U3027 ( .A1(n318), .A2(n580), .B1(\unit_memory/DRAM/n3057 ), .B2(
        n585), .ZN(\unit_memory/DRAM/n1490 ) );
  OAI22_X1 U3028 ( .A1(n321), .A2(n580), .B1(\unit_memory/DRAM/n3058 ), .B2(
        n585), .ZN(\unit_memory/DRAM/n1489 ) );
  OAI22_X1 U3029 ( .A1(n324), .A2(n579), .B1(\unit_memory/DRAM/n3059 ), .B2(
        n586), .ZN(\unit_memory/DRAM/n1488 ) );
  OAI22_X1 U3030 ( .A1(n327), .A2(n579), .B1(\unit_memory/DRAM/n3060 ), .B2(
        n586), .ZN(\unit_memory/DRAM/n1487 ) );
  OAI22_X1 U3031 ( .A1(n330), .A2(n579), .B1(\unit_memory/DRAM/n3061 ), .B2(
        n586), .ZN(\unit_memory/DRAM/n1486 ) );
  OAI22_X1 U3032 ( .A1(n333), .A2(n579), .B1(\unit_memory/DRAM/n3062 ), .B2(
        n586), .ZN(\unit_memory/DRAM/n1485 ) );
  OAI22_X1 U3033 ( .A1(n336), .A2(n579), .B1(\unit_memory/DRAM/n3063 ), .B2(
        n587), .ZN(\unit_memory/DRAM/n1484 ) );
  OAI22_X1 U3034 ( .A1(n339), .A2(n579), .B1(\unit_memory/DRAM/n3064 ), .B2(
        n587), .ZN(\unit_memory/DRAM/n1483 ) );
  OAI22_X1 U3035 ( .A1(n342), .A2(n579), .B1(\unit_memory/DRAM/n3065 ), .B2(
        n587), .ZN(\unit_memory/DRAM/n1482 ) );
  OAI22_X1 U3036 ( .A1(n345), .A2(n579), .B1(\unit_memory/DRAM/n3066 ), .B2(
        n587), .ZN(\unit_memory/DRAM/n1481 ) );
  OAI22_X1 U3037 ( .A1(n348), .A2(n579), .B1(\unit_memory/DRAM/n3067 ), .B2(
        n588), .ZN(\unit_memory/DRAM/n1480 ) );
  OAI22_X1 U3038 ( .A1(n351), .A2(n579), .B1(\unit_memory/DRAM/n3068 ), .B2(
        n588), .ZN(\unit_memory/DRAM/n1479 ) );
  OAI22_X1 U3039 ( .A1(n354), .A2(n579), .B1(\unit_memory/DRAM/n3069 ), .B2(
        n588), .ZN(\unit_memory/DRAM/n1478 ) );
  OAI22_X1 U3040 ( .A1(n357), .A2(n579), .B1(\unit_memory/DRAM/n3070 ), .B2(
        n588), .ZN(\unit_memory/DRAM/n1477 ) );
  OAI22_X1 U3041 ( .A1(n249), .A2(n612), .B1(\unit_memory/DRAM/n3135 ), .B2(
        n614), .ZN(\unit_memory/DRAM/n1412 ) );
  OAI22_X1 U3042 ( .A1(n268), .A2(n613), .B1(\unit_memory/DRAM/n3136 ), .B2(
        n614), .ZN(\unit_memory/DRAM/n1411 ) );
  OAI22_X1 U3043 ( .A1(n271), .A2(n613), .B1(\unit_memory/DRAM/n3137 ), .B2(
        n614), .ZN(\unit_memory/DRAM/n1410 ) );
  OAI22_X1 U3044 ( .A1(n274), .A2(n612), .B1(\unit_memory/DRAM/n3138 ), .B2(
        n614), .ZN(\unit_memory/DRAM/n1409 ) );
  OAI22_X1 U3045 ( .A1(n277), .A2(n613), .B1(\unit_memory/DRAM/n3139 ), .B2(
        n615), .ZN(\unit_memory/DRAM/n1408 ) );
  OAI22_X1 U3046 ( .A1(n280), .A2(n612), .B1(\unit_memory/DRAM/n3140 ), .B2(
        n615), .ZN(\unit_memory/DRAM/n1407 ) );
  OAI22_X1 U3047 ( .A1(n283), .A2(n613), .B1(\unit_memory/DRAM/n3141 ), .B2(
        n615), .ZN(\unit_memory/DRAM/n1406 ) );
  OAI22_X1 U3048 ( .A1(n286), .A2(n612), .B1(\unit_memory/DRAM/n3142 ), .B2(
        n615), .ZN(\unit_memory/DRAM/n1405 ) );
  OAI22_X1 U3049 ( .A1(n249), .A2(n623), .B1(\unit_memory/DRAM/n3167 ), .B2(
        n625), .ZN(\unit_memory/DRAM/n1380 ) );
  OAI22_X1 U3050 ( .A1(n268), .A2(n624), .B1(\unit_memory/DRAM/n3168 ), .B2(
        n625), .ZN(\unit_memory/DRAM/n1379 ) );
  OAI22_X1 U3051 ( .A1(n271), .A2(n624), .B1(\unit_memory/DRAM/n3169 ), .B2(
        n625), .ZN(\unit_memory/DRAM/n1378 ) );
  OAI22_X1 U3052 ( .A1(n274), .A2(n623), .B1(\unit_memory/DRAM/n3170 ), .B2(
        n625), .ZN(\unit_memory/DRAM/n1377 ) );
  OAI22_X1 U3053 ( .A1(n277), .A2(n624), .B1(\unit_memory/DRAM/n3171 ), .B2(
        n626), .ZN(\unit_memory/DRAM/n1376 ) );
  OAI22_X1 U3054 ( .A1(n280), .A2(n623), .B1(\unit_memory/DRAM/n3172 ), .B2(
        n626), .ZN(\unit_memory/DRAM/n1375 ) );
  OAI22_X1 U3055 ( .A1(n283), .A2(n624), .B1(\unit_memory/DRAM/n3173 ), .B2(
        n626), .ZN(\unit_memory/DRAM/n1374 ) );
  OAI22_X1 U3056 ( .A1(n286), .A2(n623), .B1(\unit_memory/DRAM/n3174 ), .B2(
        n626), .ZN(\unit_memory/DRAM/n1373 ) );
  OAI22_X1 U3057 ( .A1(n289), .A2(n624), .B1(\unit_memory/DRAM/n3175 ), .B2(
        n627), .ZN(\unit_memory/DRAM/n1372 ) );
  OAI22_X1 U3058 ( .A1(n292), .A2(n624), .B1(\unit_memory/DRAM/n3176 ), .B2(
        n627), .ZN(\unit_memory/DRAM/n1371 ) );
  OAI22_X1 U3059 ( .A1(n295), .A2(n624), .B1(\unit_memory/DRAM/n3177 ), .B2(
        n627), .ZN(\unit_memory/DRAM/n1370 ) );
  OAI22_X1 U3060 ( .A1(n298), .A2(n624), .B1(\unit_memory/DRAM/n3178 ), .B2(
        n627), .ZN(\unit_memory/DRAM/n1369 ) );
  OAI22_X1 U3061 ( .A1(n301), .A2(n624), .B1(\unit_memory/DRAM/n3179 ), .B2(
        n628), .ZN(\unit_memory/DRAM/n1368 ) );
  OAI22_X1 U3062 ( .A1(n304), .A2(n624), .B1(\unit_memory/DRAM/n3180 ), .B2(
        n628), .ZN(\unit_memory/DRAM/n1367 ) );
  OAI22_X1 U3063 ( .A1(n307), .A2(n624), .B1(\unit_memory/DRAM/n3181 ), .B2(
        n628), .ZN(\unit_memory/DRAM/n1366 ) );
  OAI22_X1 U3064 ( .A1(n310), .A2(n624), .B1(\unit_memory/DRAM/n3182 ), .B2(
        n628), .ZN(\unit_memory/DRAM/n1365 ) );
  OAI22_X1 U3065 ( .A1(n313), .A2(n624), .B1(\unit_memory/DRAM/n3183 ), .B2(
        n629), .ZN(\unit_memory/DRAM/n1364 ) );
  OAI22_X1 U3066 ( .A1(n316), .A2(n624), .B1(\unit_memory/DRAM/n3184 ), .B2(
        n629), .ZN(\unit_memory/DRAM/n1363 ) );
  OAI22_X1 U3067 ( .A1(n319), .A2(n624), .B1(\unit_memory/DRAM/n3185 ), .B2(
        n629), .ZN(\unit_memory/DRAM/n1362 ) );
  OAI22_X1 U3068 ( .A1(n322), .A2(n624), .B1(\unit_memory/DRAM/n3186 ), .B2(
        n629), .ZN(\unit_memory/DRAM/n1361 ) );
  OAI22_X1 U3069 ( .A1(n325), .A2(n623), .B1(\unit_memory/DRAM/n3187 ), .B2(
        n630), .ZN(\unit_memory/DRAM/n1360 ) );
  OAI22_X1 U3070 ( .A1(n328), .A2(n623), .B1(\unit_memory/DRAM/n3188 ), .B2(
        n630), .ZN(\unit_memory/DRAM/n1359 ) );
  OAI22_X1 U3071 ( .A1(n331), .A2(n623), .B1(\unit_memory/DRAM/n3189 ), .B2(
        n630), .ZN(\unit_memory/DRAM/n1358 ) );
  OAI22_X1 U3072 ( .A1(n334), .A2(n623), .B1(\unit_memory/DRAM/n3190 ), .B2(
        n630), .ZN(\unit_memory/DRAM/n1357 ) );
  OAI22_X1 U3073 ( .A1(n337), .A2(n623), .B1(\unit_memory/DRAM/n3191 ), .B2(
        n631), .ZN(\unit_memory/DRAM/n1356 ) );
  OAI22_X1 U3074 ( .A1(n340), .A2(n623), .B1(\unit_memory/DRAM/n3192 ), .B2(
        n631), .ZN(\unit_memory/DRAM/n1355 ) );
  OAI22_X1 U3075 ( .A1(n343), .A2(n623), .B1(\unit_memory/DRAM/n3193 ), .B2(
        n631), .ZN(\unit_memory/DRAM/n1354 ) );
  OAI22_X1 U3076 ( .A1(n346), .A2(n623), .B1(\unit_memory/DRAM/n3194 ), .B2(
        n631), .ZN(\unit_memory/DRAM/n1353 ) );
  OAI22_X1 U3077 ( .A1(n349), .A2(n623), .B1(\unit_memory/DRAM/n3195 ), .B2(
        n632), .ZN(\unit_memory/DRAM/n1352 ) );
  OAI22_X1 U3078 ( .A1(n352), .A2(n623), .B1(\unit_memory/DRAM/n3196 ), .B2(
        n632), .ZN(\unit_memory/DRAM/n1351 ) );
  OAI22_X1 U3079 ( .A1(n355), .A2(n623), .B1(\unit_memory/DRAM/n3197 ), .B2(
        n632), .ZN(\unit_memory/DRAM/n1350 ) );
  OAI22_X1 U3080 ( .A1(n357), .A2(n623), .B1(\unit_memory/DRAM/n3198 ), .B2(
        n632), .ZN(\unit_memory/DRAM/n1349 ) );
  OAI22_X1 U3081 ( .A1(n249), .A2(n657), .B1(\unit_memory/DRAM/n3263 ), .B2(
        n658), .ZN(\unit_memory/DRAM/n1284 ) );
  OAI22_X1 U3082 ( .A1(n268), .A2(n656), .B1(\unit_memory/DRAM/n3264 ), .B2(
        n658), .ZN(\unit_memory/DRAM/n1283 ) );
  OAI22_X1 U3083 ( .A1(n271), .A2(n657), .B1(\unit_memory/DRAM/n3265 ), .B2(
        n658), .ZN(\unit_memory/DRAM/n1282 ) );
  OAI22_X1 U3084 ( .A1(n274), .A2(n656), .B1(\unit_memory/DRAM/n3266 ), .B2(
        n658), .ZN(\unit_memory/DRAM/n1281 ) );
  OAI22_X1 U3085 ( .A1(n277), .A2(n657), .B1(\unit_memory/DRAM/n3267 ), .B2(
        n659), .ZN(\unit_memory/DRAM/n1280 ) );
  OAI22_X1 U3086 ( .A1(n280), .A2(n656), .B1(\unit_memory/DRAM/n3268 ), .B2(
        n659), .ZN(\unit_memory/DRAM/n1279 ) );
  OAI22_X1 U3087 ( .A1(n283), .A2(n657), .B1(\unit_memory/DRAM/n3269 ), .B2(
        n659), .ZN(\unit_memory/DRAM/n1278 ) );
  OAI22_X1 U3088 ( .A1(n286), .A2(n656), .B1(\unit_memory/DRAM/n3270 ), .B2(
        n659), .ZN(\unit_memory/DRAM/n1277 ) );
  OAI22_X1 U3089 ( .A1(n249), .A2(n668), .B1(\unit_memory/DRAM/n3295 ), .B2(
        n669), .ZN(\unit_memory/DRAM/n1252 ) );
  OAI22_X1 U3090 ( .A1(n268), .A2(n667), .B1(\unit_memory/DRAM/n3296 ), .B2(
        n669), .ZN(\unit_memory/DRAM/n1251 ) );
  OAI22_X1 U3091 ( .A1(n271), .A2(n668), .B1(\unit_memory/DRAM/n3297 ), .B2(
        n669), .ZN(\unit_memory/DRAM/n1250 ) );
  OAI22_X1 U3092 ( .A1(n274), .A2(n667), .B1(\unit_memory/DRAM/n3298 ), .B2(
        n669), .ZN(\unit_memory/DRAM/n1249 ) );
  OAI22_X1 U3093 ( .A1(n277), .A2(n668), .B1(\unit_memory/DRAM/n3299 ), .B2(
        n670), .ZN(\unit_memory/DRAM/n1248 ) );
  OAI22_X1 U3094 ( .A1(n280), .A2(n667), .B1(\unit_memory/DRAM/n3300 ), .B2(
        n670), .ZN(\unit_memory/DRAM/n1247 ) );
  OAI22_X1 U3095 ( .A1(n283), .A2(n668), .B1(\unit_memory/DRAM/n3301 ), .B2(
        n670), .ZN(\unit_memory/DRAM/n1246 ) );
  OAI22_X1 U3096 ( .A1(n286), .A2(n667), .B1(\unit_memory/DRAM/n3302 ), .B2(
        n670), .ZN(\unit_memory/DRAM/n1245 ) );
  OAI22_X1 U3097 ( .A1(n289), .A2(n668), .B1(\unit_memory/DRAM/n3303 ), .B2(
        n671), .ZN(\unit_memory/DRAM/n1244 ) );
  OAI22_X1 U3098 ( .A1(n292), .A2(n668), .B1(\unit_memory/DRAM/n3304 ), .B2(
        n671), .ZN(\unit_memory/DRAM/n1243 ) );
  OAI22_X1 U3099 ( .A1(n295), .A2(n668), .B1(\unit_memory/DRAM/n3305 ), .B2(
        n671), .ZN(\unit_memory/DRAM/n1242 ) );
  OAI22_X1 U3100 ( .A1(n298), .A2(n668), .B1(\unit_memory/DRAM/n3306 ), .B2(
        n671), .ZN(\unit_memory/DRAM/n1241 ) );
  OAI22_X1 U3101 ( .A1(n301), .A2(n668), .B1(\unit_memory/DRAM/n3307 ), .B2(
        n672), .ZN(\unit_memory/DRAM/n1240 ) );
  OAI22_X1 U3102 ( .A1(n304), .A2(n668), .B1(\unit_memory/DRAM/n3308 ), .B2(
        n672), .ZN(\unit_memory/DRAM/n1239 ) );
  OAI22_X1 U3103 ( .A1(n307), .A2(n668), .B1(\unit_memory/DRAM/n3309 ), .B2(
        n672), .ZN(\unit_memory/DRAM/n1238 ) );
  OAI22_X1 U3104 ( .A1(n310), .A2(n668), .B1(\unit_memory/DRAM/n3310 ), .B2(
        n672), .ZN(\unit_memory/DRAM/n1237 ) );
  OAI22_X1 U3105 ( .A1(n313), .A2(n668), .B1(\unit_memory/DRAM/n3311 ), .B2(
        n673), .ZN(\unit_memory/DRAM/n1236 ) );
  OAI22_X1 U3106 ( .A1(n316), .A2(n668), .B1(\unit_memory/DRAM/n3312 ), .B2(
        n673), .ZN(\unit_memory/DRAM/n1235 ) );
  OAI22_X1 U3107 ( .A1(n319), .A2(n668), .B1(\unit_memory/DRAM/n3313 ), .B2(
        n673), .ZN(\unit_memory/DRAM/n1234 ) );
  OAI22_X1 U3108 ( .A1(n322), .A2(n668), .B1(\unit_memory/DRAM/n3314 ), .B2(
        n673), .ZN(\unit_memory/DRAM/n1233 ) );
  OAI22_X1 U3109 ( .A1(n325), .A2(n667), .B1(\unit_memory/DRAM/n3315 ), .B2(
        n674), .ZN(\unit_memory/DRAM/n1232 ) );
  OAI22_X1 U3110 ( .A1(n328), .A2(n667), .B1(\unit_memory/DRAM/n3316 ), .B2(
        n674), .ZN(\unit_memory/DRAM/n1231 ) );
  OAI22_X1 U3111 ( .A1(n331), .A2(n667), .B1(\unit_memory/DRAM/n3317 ), .B2(
        n674), .ZN(\unit_memory/DRAM/n1230 ) );
  OAI22_X1 U3112 ( .A1(n334), .A2(n667), .B1(\unit_memory/DRAM/n3318 ), .B2(
        n674), .ZN(\unit_memory/DRAM/n1229 ) );
  OAI22_X1 U3113 ( .A1(n337), .A2(n667), .B1(\unit_memory/DRAM/n3319 ), .B2(
        n675), .ZN(\unit_memory/DRAM/n1228 ) );
  OAI22_X1 U3114 ( .A1(n340), .A2(n667), .B1(\unit_memory/DRAM/n3320 ), .B2(
        n675), .ZN(\unit_memory/DRAM/n1227 ) );
  OAI22_X1 U3115 ( .A1(n343), .A2(n667), .B1(\unit_memory/DRAM/n3321 ), .B2(
        n675), .ZN(\unit_memory/DRAM/n1226 ) );
  OAI22_X1 U3116 ( .A1(n346), .A2(n667), .B1(\unit_memory/DRAM/n3322 ), .B2(
        n675), .ZN(\unit_memory/DRAM/n1225 ) );
  OAI22_X1 U3117 ( .A1(n349), .A2(n667), .B1(\unit_memory/DRAM/n3323 ), .B2(
        n676), .ZN(\unit_memory/DRAM/n1224 ) );
  OAI22_X1 U3118 ( .A1(n352), .A2(n667), .B1(\unit_memory/DRAM/n3324 ), .B2(
        n676), .ZN(\unit_memory/DRAM/n1223 ) );
  OAI22_X1 U3119 ( .A1(n355), .A2(n667), .B1(\unit_memory/DRAM/n3325 ), .B2(
        n676), .ZN(\unit_memory/DRAM/n1222 ) );
  OAI22_X1 U3120 ( .A1(n358), .A2(n667), .B1(\unit_memory/DRAM/n3326 ), .B2(
        n676), .ZN(\unit_memory/DRAM/n1221 ) );
  OAI22_X1 U3121 ( .A1(n288), .A2(n525), .B1(\unit_memory/DRAM/n2887 ), .B2(
        n528), .ZN(\unit_memory/DRAM/n1660 ) );
  OAI22_X1 U3122 ( .A1(n291), .A2(n525), .B1(\unit_memory/DRAM/n2888 ), .B2(
        n528), .ZN(\unit_memory/DRAM/n1659 ) );
  OAI22_X1 U3123 ( .A1(n294), .A2(n525), .B1(\unit_memory/DRAM/n2889 ), .B2(
        n528), .ZN(\unit_memory/DRAM/n1658 ) );
  OAI22_X1 U3124 ( .A1(n297), .A2(n525), .B1(\unit_memory/DRAM/n2890 ), .B2(
        n528), .ZN(\unit_memory/DRAM/n1657 ) );
  OAI22_X1 U3125 ( .A1(n300), .A2(n525), .B1(\unit_memory/DRAM/n2891 ), .B2(
        n529), .ZN(\unit_memory/DRAM/n1656 ) );
  OAI22_X1 U3126 ( .A1(n303), .A2(n525), .B1(\unit_memory/DRAM/n2892 ), .B2(
        n529), .ZN(\unit_memory/DRAM/n1655 ) );
  OAI22_X1 U3127 ( .A1(n306), .A2(n525), .B1(\unit_memory/DRAM/n2893 ), .B2(
        n529), .ZN(\unit_memory/DRAM/n1654 ) );
  OAI22_X1 U3128 ( .A1(n309), .A2(n525), .B1(\unit_memory/DRAM/n2894 ), .B2(
        n529), .ZN(\unit_memory/DRAM/n1653 ) );
  OAI22_X1 U3129 ( .A1(n312), .A2(n525), .B1(\unit_memory/DRAM/n2895 ), .B2(
        n530), .ZN(\unit_memory/DRAM/n1652 ) );
  OAI22_X1 U3130 ( .A1(n315), .A2(n525), .B1(\unit_memory/DRAM/n2896 ), .B2(
        n530), .ZN(\unit_memory/DRAM/n1651 ) );
  OAI22_X1 U3131 ( .A1(n318), .A2(n525), .B1(\unit_memory/DRAM/n2897 ), .B2(
        n530), .ZN(\unit_memory/DRAM/n1650 ) );
  OAI22_X1 U3132 ( .A1(n321), .A2(n525), .B1(\unit_memory/DRAM/n2898 ), .B2(
        n530), .ZN(\unit_memory/DRAM/n1649 ) );
  OAI22_X1 U3133 ( .A1(n324), .A2(n524), .B1(\unit_memory/DRAM/n2899 ), .B2(
        n531), .ZN(\unit_memory/DRAM/n1648 ) );
  OAI22_X1 U3134 ( .A1(n327), .A2(n524), .B1(\unit_memory/DRAM/n2900 ), .B2(
        n531), .ZN(\unit_memory/DRAM/n1647 ) );
  OAI22_X1 U3135 ( .A1(n330), .A2(n524), .B1(\unit_memory/DRAM/n2901 ), .B2(
        n531), .ZN(\unit_memory/DRAM/n1646 ) );
  OAI22_X1 U3136 ( .A1(n333), .A2(n524), .B1(\unit_memory/DRAM/n2902 ), .B2(
        n531), .ZN(\unit_memory/DRAM/n1645 ) );
  OAI22_X1 U3137 ( .A1(n336), .A2(n524), .B1(\unit_memory/DRAM/n2903 ), .B2(
        n532), .ZN(\unit_memory/DRAM/n1644 ) );
  OAI22_X1 U3138 ( .A1(n339), .A2(n524), .B1(\unit_memory/DRAM/n2904 ), .B2(
        n532), .ZN(\unit_memory/DRAM/n1643 ) );
  OAI22_X1 U3139 ( .A1(n342), .A2(n524), .B1(\unit_memory/DRAM/n2905 ), .B2(
        n532), .ZN(\unit_memory/DRAM/n1642 ) );
  OAI22_X1 U3140 ( .A1(n345), .A2(n524), .B1(\unit_memory/DRAM/n2906 ), .B2(
        n532), .ZN(\unit_memory/DRAM/n1641 ) );
  OAI22_X1 U3141 ( .A1(n348), .A2(n524), .B1(\unit_memory/DRAM/n2907 ), .B2(
        n533), .ZN(\unit_memory/DRAM/n1640 ) );
  OAI22_X1 U3142 ( .A1(n351), .A2(n524), .B1(\unit_memory/DRAM/n2908 ), .B2(
        n533), .ZN(\unit_memory/DRAM/n1639 ) );
  OAI22_X1 U3143 ( .A1(n354), .A2(n524), .B1(\unit_memory/DRAM/n2909 ), .B2(
        n533), .ZN(\unit_memory/DRAM/n1638 ) );
  OAI22_X1 U3144 ( .A1(n357), .A2(n524), .B1(\unit_memory/DRAM/n2910 ), .B2(
        n533), .ZN(\unit_memory/DRAM/n1637 ) );
  OAI22_X1 U3145 ( .A1(n250), .A2(n547), .B1(\unit_memory/DRAM/n2943 ), .B2(
        n548), .ZN(\unit_memory/DRAM/n1604 ) );
  OAI22_X1 U3146 ( .A1(n267), .A2(n546), .B1(\unit_memory/DRAM/n2944 ), .B2(
        n548), .ZN(\unit_memory/DRAM/n1603 ) );
  OAI22_X1 U3147 ( .A1(n270), .A2(n547), .B1(\unit_memory/DRAM/n2945 ), .B2(
        n548), .ZN(\unit_memory/DRAM/n1602 ) );
  OAI22_X1 U3148 ( .A1(n273), .A2(n546), .B1(\unit_memory/DRAM/n2946 ), .B2(
        n548), .ZN(\unit_memory/DRAM/n1601 ) );
  OAI22_X1 U3149 ( .A1(n276), .A2(n547), .B1(\unit_memory/DRAM/n2947 ), .B2(
        n549), .ZN(\unit_memory/DRAM/n1600 ) );
  OAI22_X1 U3150 ( .A1(n279), .A2(n546), .B1(\unit_memory/DRAM/n2948 ), .B2(
        n549), .ZN(\unit_memory/DRAM/n1599 ) );
  OAI22_X1 U3151 ( .A1(n282), .A2(n547), .B1(\unit_memory/DRAM/n2949 ), .B2(
        n549), .ZN(\unit_memory/DRAM/n1598 ) );
  OAI22_X1 U3152 ( .A1(n285), .A2(n546), .B1(\unit_memory/DRAM/n2950 ), .B2(
        n549), .ZN(\unit_memory/DRAM/n1597 ) );
  OAI22_X1 U3153 ( .A1(n288), .A2(n547), .B1(\unit_memory/DRAM/n2951 ), .B2(
        n550), .ZN(\unit_memory/DRAM/n1596 ) );
  OAI22_X1 U3154 ( .A1(n291), .A2(n547), .B1(\unit_memory/DRAM/n2952 ), .B2(
        n550), .ZN(\unit_memory/DRAM/n1595 ) );
  OAI22_X1 U3155 ( .A1(n294), .A2(n547), .B1(\unit_memory/DRAM/n2953 ), .B2(
        n550), .ZN(\unit_memory/DRAM/n1594 ) );
  OAI22_X1 U3156 ( .A1(n297), .A2(n547), .B1(\unit_memory/DRAM/n2954 ), .B2(
        n550), .ZN(\unit_memory/DRAM/n1593 ) );
  OAI22_X1 U3157 ( .A1(n300), .A2(n547), .B1(\unit_memory/DRAM/n2955 ), .B2(
        n551), .ZN(\unit_memory/DRAM/n1592 ) );
  OAI22_X1 U3158 ( .A1(n303), .A2(n547), .B1(\unit_memory/DRAM/n2956 ), .B2(
        n551), .ZN(\unit_memory/DRAM/n1591 ) );
  OAI22_X1 U3159 ( .A1(n306), .A2(n547), .B1(\unit_memory/DRAM/n2957 ), .B2(
        n551), .ZN(\unit_memory/DRAM/n1590 ) );
  OAI22_X1 U3160 ( .A1(n309), .A2(n547), .B1(\unit_memory/DRAM/n2958 ), .B2(
        n551), .ZN(\unit_memory/DRAM/n1589 ) );
  OAI22_X1 U3161 ( .A1(n312), .A2(n547), .B1(\unit_memory/DRAM/n2959 ), .B2(
        n552), .ZN(\unit_memory/DRAM/n1588 ) );
  OAI22_X1 U3162 ( .A1(n315), .A2(n547), .B1(\unit_memory/DRAM/n2960 ), .B2(
        n552), .ZN(\unit_memory/DRAM/n1587 ) );
  OAI22_X1 U3163 ( .A1(n318), .A2(n547), .B1(\unit_memory/DRAM/n2961 ), .B2(
        n552), .ZN(\unit_memory/DRAM/n1586 ) );
  OAI22_X1 U3164 ( .A1(n321), .A2(n547), .B1(\unit_memory/DRAM/n2962 ), .B2(
        n552), .ZN(\unit_memory/DRAM/n1585 ) );
  OAI22_X1 U3165 ( .A1(n324), .A2(n546), .B1(\unit_memory/DRAM/n2963 ), .B2(
        n553), .ZN(\unit_memory/DRAM/n1584 ) );
  OAI22_X1 U3166 ( .A1(n327), .A2(n546), .B1(\unit_memory/DRAM/n2964 ), .B2(
        n553), .ZN(\unit_memory/DRAM/n1583 ) );
  OAI22_X1 U3167 ( .A1(n330), .A2(n546), .B1(\unit_memory/DRAM/n2965 ), .B2(
        n553), .ZN(\unit_memory/DRAM/n1582 ) );
  OAI22_X1 U3168 ( .A1(n333), .A2(n546), .B1(\unit_memory/DRAM/n2966 ), .B2(
        n553), .ZN(\unit_memory/DRAM/n1581 ) );
  OAI22_X1 U3169 ( .A1(n336), .A2(n546), .B1(\unit_memory/DRAM/n2967 ), .B2(
        n554), .ZN(\unit_memory/DRAM/n1580 ) );
  OAI22_X1 U3170 ( .A1(n339), .A2(n546), .B1(\unit_memory/DRAM/n2968 ), .B2(
        n554), .ZN(\unit_memory/DRAM/n1579 ) );
  OAI22_X1 U3171 ( .A1(n342), .A2(n546), .B1(\unit_memory/DRAM/n2969 ), .B2(
        n554), .ZN(\unit_memory/DRAM/n1578 ) );
  OAI22_X1 U3172 ( .A1(n345), .A2(n546), .B1(\unit_memory/DRAM/n2970 ), .B2(
        n554), .ZN(\unit_memory/DRAM/n1577 ) );
  OAI22_X1 U3173 ( .A1(n348), .A2(n546), .B1(\unit_memory/DRAM/n2971 ), .B2(
        n555), .ZN(\unit_memory/DRAM/n1576 ) );
  OAI22_X1 U3174 ( .A1(n351), .A2(n546), .B1(\unit_memory/DRAM/n2972 ), .B2(
        n555), .ZN(\unit_memory/DRAM/n1575 ) );
  OAI22_X1 U3175 ( .A1(n354), .A2(n546), .B1(\unit_memory/DRAM/n2973 ), .B2(
        n555), .ZN(\unit_memory/DRAM/n1574 ) );
  OAI22_X1 U3176 ( .A1(n357), .A2(n546), .B1(\unit_memory/DRAM/n2974 ), .B2(
        n555), .ZN(\unit_memory/DRAM/n1573 ) );
  OAI22_X1 U3177 ( .A1(n250), .A2(n558), .B1(\unit_memory/DRAM/n2975 ), .B2(
        n559), .ZN(\unit_memory/DRAM/n1572 ) );
  OAI22_X1 U3178 ( .A1(n267), .A2(n557), .B1(\unit_memory/DRAM/n2976 ), .B2(
        n559), .ZN(\unit_memory/DRAM/n1571 ) );
  OAI22_X1 U3179 ( .A1(n270), .A2(n558), .B1(\unit_memory/DRAM/n2977 ), .B2(
        n559), .ZN(\unit_memory/DRAM/n1570 ) );
  OAI22_X1 U3180 ( .A1(n273), .A2(n557), .B1(\unit_memory/DRAM/n2978 ), .B2(
        n559), .ZN(\unit_memory/DRAM/n1569 ) );
  OAI22_X1 U3181 ( .A1(n276), .A2(n558), .B1(\unit_memory/DRAM/n2979 ), .B2(
        n560), .ZN(\unit_memory/DRAM/n1568 ) );
  OAI22_X1 U3182 ( .A1(n279), .A2(n557), .B1(\unit_memory/DRAM/n2980 ), .B2(
        n560), .ZN(\unit_memory/DRAM/n1567 ) );
  OAI22_X1 U3183 ( .A1(n282), .A2(n558), .B1(\unit_memory/DRAM/n2981 ), .B2(
        n560), .ZN(\unit_memory/DRAM/n1566 ) );
  OAI22_X1 U3184 ( .A1(n285), .A2(n557), .B1(\unit_memory/DRAM/n2982 ), .B2(
        n560), .ZN(\unit_memory/DRAM/n1565 ) );
  OAI22_X1 U3185 ( .A1(n288), .A2(n558), .B1(\unit_memory/DRAM/n2983 ), .B2(
        n561), .ZN(\unit_memory/DRAM/n1564 ) );
  OAI22_X1 U3186 ( .A1(n291), .A2(n558), .B1(\unit_memory/DRAM/n2984 ), .B2(
        n561), .ZN(\unit_memory/DRAM/n1563 ) );
  OAI22_X1 U3187 ( .A1(n294), .A2(n558), .B1(\unit_memory/DRAM/n2985 ), .B2(
        n561), .ZN(\unit_memory/DRAM/n1562 ) );
  OAI22_X1 U3188 ( .A1(n297), .A2(n558), .B1(\unit_memory/DRAM/n2986 ), .B2(
        n561), .ZN(\unit_memory/DRAM/n1561 ) );
  OAI22_X1 U3189 ( .A1(n300), .A2(n558), .B1(\unit_memory/DRAM/n2987 ), .B2(
        n562), .ZN(\unit_memory/DRAM/n1560 ) );
  OAI22_X1 U3190 ( .A1(n303), .A2(n558), .B1(\unit_memory/DRAM/n2988 ), .B2(
        n562), .ZN(\unit_memory/DRAM/n1559 ) );
  OAI22_X1 U3191 ( .A1(n306), .A2(n558), .B1(\unit_memory/DRAM/n2989 ), .B2(
        n562), .ZN(\unit_memory/DRAM/n1558 ) );
  OAI22_X1 U3192 ( .A1(n309), .A2(n558), .B1(\unit_memory/DRAM/n2990 ), .B2(
        n562), .ZN(\unit_memory/DRAM/n1557 ) );
  OAI22_X1 U3193 ( .A1(n312), .A2(n558), .B1(\unit_memory/DRAM/n2991 ), .B2(
        n563), .ZN(\unit_memory/DRAM/n1556 ) );
  OAI22_X1 U3194 ( .A1(n315), .A2(n558), .B1(\unit_memory/DRAM/n2992 ), .B2(
        n563), .ZN(\unit_memory/DRAM/n1555 ) );
  OAI22_X1 U3195 ( .A1(n318), .A2(n558), .B1(\unit_memory/DRAM/n2993 ), .B2(
        n563), .ZN(\unit_memory/DRAM/n1554 ) );
  OAI22_X1 U3196 ( .A1(n321), .A2(n558), .B1(\unit_memory/DRAM/n2994 ), .B2(
        n563), .ZN(\unit_memory/DRAM/n1553 ) );
  OAI22_X1 U3197 ( .A1(n324), .A2(n557), .B1(\unit_memory/DRAM/n2995 ), .B2(
        n564), .ZN(\unit_memory/DRAM/n1552 ) );
  OAI22_X1 U3198 ( .A1(n327), .A2(n557), .B1(\unit_memory/DRAM/n2996 ), .B2(
        n564), .ZN(\unit_memory/DRAM/n1551 ) );
  OAI22_X1 U3199 ( .A1(n330), .A2(n557), .B1(\unit_memory/DRAM/n2997 ), .B2(
        n564), .ZN(\unit_memory/DRAM/n1550 ) );
  OAI22_X1 U3200 ( .A1(n333), .A2(n557), .B1(\unit_memory/DRAM/n2998 ), .B2(
        n564), .ZN(\unit_memory/DRAM/n1549 ) );
  OAI22_X1 U3201 ( .A1(n336), .A2(n557), .B1(\unit_memory/DRAM/n2999 ), .B2(
        n565), .ZN(\unit_memory/DRAM/n1548 ) );
  OAI22_X1 U3202 ( .A1(n339), .A2(n557), .B1(\unit_memory/DRAM/n3000 ), .B2(
        n565), .ZN(\unit_memory/DRAM/n1547 ) );
  OAI22_X1 U3203 ( .A1(n342), .A2(n557), .B1(\unit_memory/DRAM/n3001 ), .B2(
        n565), .ZN(\unit_memory/DRAM/n1546 ) );
  OAI22_X1 U3204 ( .A1(n345), .A2(n557), .B1(\unit_memory/DRAM/n3002 ), .B2(
        n565), .ZN(\unit_memory/DRAM/n1545 ) );
  OAI22_X1 U3205 ( .A1(n348), .A2(n557), .B1(\unit_memory/DRAM/n3003 ), .B2(
        n566), .ZN(\unit_memory/DRAM/n1544 ) );
  OAI22_X1 U3206 ( .A1(n351), .A2(n557), .B1(\unit_memory/DRAM/n3004 ), .B2(
        n566), .ZN(\unit_memory/DRAM/n1543 ) );
  OAI22_X1 U3207 ( .A1(n354), .A2(n557), .B1(\unit_memory/DRAM/n3005 ), .B2(
        n566), .ZN(\unit_memory/DRAM/n1542 ) );
  OAI22_X1 U3208 ( .A1(n357), .A2(n557), .B1(\unit_memory/DRAM/n3006 ), .B2(
        n566), .ZN(\unit_memory/DRAM/n1541 ) );
  OAI22_X1 U3209 ( .A1(n288), .A2(n569), .B1(\unit_memory/DRAM/n3015 ), .B2(
        n572), .ZN(\unit_memory/DRAM/n1532 ) );
  OAI22_X1 U3210 ( .A1(n291), .A2(n569), .B1(\unit_memory/DRAM/n3016 ), .B2(
        n572), .ZN(\unit_memory/DRAM/n1531 ) );
  OAI22_X1 U3211 ( .A1(n294), .A2(n569), .B1(\unit_memory/DRAM/n3017 ), .B2(
        n572), .ZN(\unit_memory/DRAM/n1530 ) );
  OAI22_X1 U3212 ( .A1(n297), .A2(n569), .B1(\unit_memory/DRAM/n3018 ), .B2(
        n572), .ZN(\unit_memory/DRAM/n1529 ) );
  OAI22_X1 U3213 ( .A1(n300), .A2(n569), .B1(\unit_memory/DRAM/n3019 ), .B2(
        n573), .ZN(\unit_memory/DRAM/n1528 ) );
  OAI22_X1 U3214 ( .A1(n303), .A2(n569), .B1(\unit_memory/DRAM/n3020 ), .B2(
        n573), .ZN(\unit_memory/DRAM/n1527 ) );
  OAI22_X1 U3215 ( .A1(n306), .A2(n569), .B1(\unit_memory/DRAM/n3021 ), .B2(
        n573), .ZN(\unit_memory/DRAM/n1526 ) );
  OAI22_X1 U3216 ( .A1(n309), .A2(n569), .B1(\unit_memory/DRAM/n3022 ), .B2(
        n573), .ZN(\unit_memory/DRAM/n1525 ) );
  OAI22_X1 U3217 ( .A1(n312), .A2(n569), .B1(\unit_memory/DRAM/n3023 ), .B2(
        n574), .ZN(\unit_memory/DRAM/n1524 ) );
  OAI22_X1 U3218 ( .A1(n315), .A2(n569), .B1(\unit_memory/DRAM/n3024 ), .B2(
        n574), .ZN(\unit_memory/DRAM/n1523 ) );
  OAI22_X1 U3219 ( .A1(n318), .A2(n569), .B1(\unit_memory/DRAM/n3025 ), .B2(
        n574), .ZN(\unit_memory/DRAM/n1522 ) );
  OAI22_X1 U3220 ( .A1(n321), .A2(n569), .B1(\unit_memory/DRAM/n3026 ), .B2(
        n574), .ZN(\unit_memory/DRAM/n1521 ) );
  OAI22_X1 U3221 ( .A1(n324), .A2(n568), .B1(\unit_memory/DRAM/n3027 ), .B2(
        n575), .ZN(\unit_memory/DRAM/n1520 ) );
  OAI22_X1 U3222 ( .A1(n327), .A2(n568), .B1(\unit_memory/DRAM/n3028 ), .B2(
        n575), .ZN(\unit_memory/DRAM/n1519 ) );
  OAI22_X1 U3223 ( .A1(n330), .A2(n568), .B1(\unit_memory/DRAM/n3029 ), .B2(
        n575), .ZN(\unit_memory/DRAM/n1518 ) );
  OAI22_X1 U3224 ( .A1(n333), .A2(n568), .B1(\unit_memory/DRAM/n3030 ), .B2(
        n575), .ZN(\unit_memory/DRAM/n1517 ) );
  OAI22_X1 U3225 ( .A1(n336), .A2(n568), .B1(\unit_memory/DRAM/n3031 ), .B2(
        n576), .ZN(\unit_memory/DRAM/n1516 ) );
  OAI22_X1 U3226 ( .A1(n339), .A2(n568), .B1(\unit_memory/DRAM/n3032 ), .B2(
        n576), .ZN(\unit_memory/DRAM/n1515 ) );
  OAI22_X1 U3227 ( .A1(n342), .A2(n568), .B1(\unit_memory/DRAM/n3033 ), .B2(
        n576), .ZN(\unit_memory/DRAM/n1514 ) );
  OAI22_X1 U3228 ( .A1(n345), .A2(n568), .B1(\unit_memory/DRAM/n3034 ), .B2(
        n576), .ZN(\unit_memory/DRAM/n1513 ) );
  OAI22_X1 U3229 ( .A1(n348), .A2(n568), .B1(\unit_memory/DRAM/n3035 ), .B2(
        n577), .ZN(\unit_memory/DRAM/n1512 ) );
  OAI22_X1 U3230 ( .A1(n351), .A2(n568), .B1(\unit_memory/DRAM/n3036 ), .B2(
        n577), .ZN(\unit_memory/DRAM/n1511 ) );
  OAI22_X1 U3231 ( .A1(n354), .A2(n568), .B1(\unit_memory/DRAM/n3037 ), .B2(
        n577), .ZN(\unit_memory/DRAM/n1510 ) );
  OAI22_X1 U3232 ( .A1(n357), .A2(n568), .B1(\unit_memory/DRAM/n3038 ), .B2(
        n577), .ZN(\unit_memory/DRAM/n1509 ) );
  OAI22_X1 U3233 ( .A1(n249), .A2(n591), .B1(\unit_memory/DRAM/n3071 ), .B2(
        n592), .ZN(\unit_memory/DRAM/n1476 ) );
  OAI22_X1 U3234 ( .A1(n267), .A2(n590), .B1(\unit_memory/DRAM/n3072 ), .B2(
        n592), .ZN(\unit_memory/DRAM/n1475 ) );
  OAI22_X1 U3235 ( .A1(n270), .A2(n591), .B1(\unit_memory/DRAM/n3073 ), .B2(
        n592), .ZN(\unit_memory/DRAM/n1474 ) );
  OAI22_X1 U3236 ( .A1(n273), .A2(n590), .B1(\unit_memory/DRAM/n3074 ), .B2(
        n592), .ZN(\unit_memory/DRAM/n1473 ) );
  OAI22_X1 U3237 ( .A1(n276), .A2(n591), .B1(\unit_memory/DRAM/n3075 ), .B2(
        n593), .ZN(\unit_memory/DRAM/n1472 ) );
  OAI22_X1 U3238 ( .A1(n279), .A2(n590), .B1(\unit_memory/DRAM/n3076 ), .B2(
        n593), .ZN(\unit_memory/DRAM/n1471 ) );
  OAI22_X1 U3239 ( .A1(n282), .A2(n591), .B1(\unit_memory/DRAM/n3077 ), .B2(
        n593), .ZN(\unit_memory/DRAM/n1470 ) );
  OAI22_X1 U3240 ( .A1(n285), .A2(n590), .B1(\unit_memory/DRAM/n3078 ), .B2(
        n593), .ZN(\unit_memory/DRAM/n1469 ) );
  OAI22_X1 U3241 ( .A1(n288), .A2(n591), .B1(\unit_memory/DRAM/n3079 ), .B2(
        n594), .ZN(\unit_memory/DRAM/n1468 ) );
  OAI22_X1 U3242 ( .A1(n291), .A2(n591), .B1(\unit_memory/DRAM/n3080 ), .B2(
        n594), .ZN(\unit_memory/DRAM/n1467 ) );
  OAI22_X1 U3243 ( .A1(n294), .A2(n591), .B1(\unit_memory/DRAM/n3081 ), .B2(
        n594), .ZN(\unit_memory/DRAM/n1466 ) );
  OAI22_X1 U3244 ( .A1(n297), .A2(n591), .B1(\unit_memory/DRAM/n3082 ), .B2(
        n594), .ZN(\unit_memory/DRAM/n1465 ) );
  OAI22_X1 U3245 ( .A1(n300), .A2(n591), .B1(\unit_memory/DRAM/n3083 ), .B2(
        n595), .ZN(\unit_memory/DRAM/n1464 ) );
  OAI22_X1 U3246 ( .A1(n303), .A2(n591), .B1(\unit_memory/DRAM/n3084 ), .B2(
        n595), .ZN(\unit_memory/DRAM/n1463 ) );
  OAI22_X1 U3247 ( .A1(n306), .A2(n591), .B1(\unit_memory/DRAM/n3085 ), .B2(
        n595), .ZN(\unit_memory/DRAM/n1462 ) );
  OAI22_X1 U3248 ( .A1(n309), .A2(n591), .B1(\unit_memory/DRAM/n3086 ), .B2(
        n595), .ZN(\unit_memory/DRAM/n1461 ) );
  OAI22_X1 U3249 ( .A1(n312), .A2(n591), .B1(\unit_memory/DRAM/n3087 ), .B2(
        n596), .ZN(\unit_memory/DRAM/n1460 ) );
  OAI22_X1 U3250 ( .A1(n315), .A2(n591), .B1(\unit_memory/DRAM/n3088 ), .B2(
        n596), .ZN(\unit_memory/DRAM/n1459 ) );
  OAI22_X1 U3251 ( .A1(n318), .A2(n591), .B1(\unit_memory/DRAM/n3089 ), .B2(
        n596), .ZN(\unit_memory/DRAM/n1458 ) );
  OAI22_X1 U3252 ( .A1(n321), .A2(n591), .B1(\unit_memory/DRAM/n3090 ), .B2(
        n596), .ZN(\unit_memory/DRAM/n1457 ) );
  OAI22_X1 U3253 ( .A1(n324), .A2(n590), .B1(\unit_memory/DRAM/n3091 ), .B2(
        n597), .ZN(\unit_memory/DRAM/n1456 ) );
  OAI22_X1 U3254 ( .A1(n327), .A2(n590), .B1(\unit_memory/DRAM/n3092 ), .B2(
        n597), .ZN(\unit_memory/DRAM/n1455 ) );
  OAI22_X1 U3255 ( .A1(n330), .A2(n590), .B1(\unit_memory/DRAM/n3093 ), .B2(
        n597), .ZN(\unit_memory/DRAM/n1454 ) );
  OAI22_X1 U3256 ( .A1(n333), .A2(n590), .B1(\unit_memory/DRAM/n3094 ), .B2(
        n597), .ZN(\unit_memory/DRAM/n1453 ) );
  OAI22_X1 U3257 ( .A1(n336), .A2(n590), .B1(\unit_memory/DRAM/n3095 ), .B2(
        n598), .ZN(\unit_memory/DRAM/n1452 ) );
  OAI22_X1 U3258 ( .A1(n339), .A2(n590), .B1(\unit_memory/DRAM/n3096 ), .B2(
        n598), .ZN(\unit_memory/DRAM/n1451 ) );
  OAI22_X1 U3259 ( .A1(n342), .A2(n590), .B1(\unit_memory/DRAM/n3097 ), .B2(
        n598), .ZN(\unit_memory/DRAM/n1450 ) );
  OAI22_X1 U3260 ( .A1(n345), .A2(n590), .B1(\unit_memory/DRAM/n3098 ), .B2(
        n598), .ZN(\unit_memory/DRAM/n1449 ) );
  OAI22_X1 U3261 ( .A1(n348), .A2(n590), .B1(\unit_memory/DRAM/n3099 ), .B2(
        n599), .ZN(\unit_memory/DRAM/n1448 ) );
  OAI22_X1 U3262 ( .A1(n351), .A2(n590), .B1(\unit_memory/DRAM/n3100 ), .B2(
        n599), .ZN(\unit_memory/DRAM/n1447 ) );
  OAI22_X1 U3263 ( .A1(n354), .A2(n590), .B1(\unit_memory/DRAM/n3101 ), .B2(
        n599), .ZN(\unit_memory/DRAM/n1446 ) );
  OAI22_X1 U3264 ( .A1(n357), .A2(n590), .B1(\unit_memory/DRAM/n3102 ), .B2(
        n599), .ZN(\unit_memory/DRAM/n1445 ) );
  OAI22_X1 U3265 ( .A1(n249), .A2(n602), .B1(\unit_memory/DRAM/n3103 ), .B2(
        n603), .ZN(\unit_memory/DRAM/n1444 ) );
  OAI22_X1 U3266 ( .A1(n267), .A2(n601), .B1(\unit_memory/DRAM/n3104 ), .B2(
        n603), .ZN(\unit_memory/DRAM/n1443 ) );
  OAI22_X1 U3267 ( .A1(n270), .A2(n602), .B1(\unit_memory/DRAM/n3105 ), .B2(
        n603), .ZN(\unit_memory/DRAM/n1442 ) );
  OAI22_X1 U3268 ( .A1(n273), .A2(n601), .B1(\unit_memory/DRAM/n3106 ), .B2(
        n603), .ZN(\unit_memory/DRAM/n1441 ) );
  OAI22_X1 U3269 ( .A1(n276), .A2(n602), .B1(\unit_memory/DRAM/n3107 ), .B2(
        n604), .ZN(\unit_memory/DRAM/n1440 ) );
  OAI22_X1 U3270 ( .A1(n279), .A2(n601), .B1(\unit_memory/DRAM/n3108 ), .B2(
        n604), .ZN(\unit_memory/DRAM/n1439 ) );
  OAI22_X1 U3271 ( .A1(n282), .A2(n602), .B1(\unit_memory/DRAM/n3109 ), .B2(
        n604), .ZN(\unit_memory/DRAM/n1438 ) );
  OAI22_X1 U3272 ( .A1(n285), .A2(n601), .B1(\unit_memory/DRAM/n3110 ), .B2(
        n604), .ZN(\unit_memory/DRAM/n1437 ) );
  OAI22_X1 U3273 ( .A1(n288), .A2(n602), .B1(\unit_memory/DRAM/n3111 ), .B2(
        n605), .ZN(\unit_memory/DRAM/n1436 ) );
  OAI22_X1 U3274 ( .A1(n291), .A2(n602), .B1(\unit_memory/DRAM/n3112 ), .B2(
        n605), .ZN(\unit_memory/DRAM/n1435 ) );
  OAI22_X1 U3275 ( .A1(n294), .A2(n602), .B1(\unit_memory/DRAM/n3113 ), .B2(
        n605), .ZN(\unit_memory/DRAM/n1434 ) );
  OAI22_X1 U3276 ( .A1(n297), .A2(n602), .B1(\unit_memory/DRAM/n3114 ), .B2(
        n605), .ZN(\unit_memory/DRAM/n1433 ) );
  OAI22_X1 U3277 ( .A1(n300), .A2(n602), .B1(\unit_memory/DRAM/n3115 ), .B2(
        n606), .ZN(\unit_memory/DRAM/n1432 ) );
  OAI22_X1 U3278 ( .A1(n303), .A2(n602), .B1(\unit_memory/DRAM/n3116 ), .B2(
        n606), .ZN(\unit_memory/DRAM/n1431 ) );
  OAI22_X1 U3279 ( .A1(n306), .A2(n602), .B1(\unit_memory/DRAM/n3117 ), .B2(
        n606), .ZN(\unit_memory/DRAM/n1430 ) );
  OAI22_X1 U3280 ( .A1(n309), .A2(n602), .B1(\unit_memory/DRAM/n3118 ), .B2(
        n606), .ZN(\unit_memory/DRAM/n1429 ) );
  OAI22_X1 U3281 ( .A1(n312), .A2(n602), .B1(\unit_memory/DRAM/n3119 ), .B2(
        n607), .ZN(\unit_memory/DRAM/n1428 ) );
  OAI22_X1 U3282 ( .A1(n315), .A2(n602), .B1(\unit_memory/DRAM/n3120 ), .B2(
        n607), .ZN(\unit_memory/DRAM/n1427 ) );
  OAI22_X1 U3283 ( .A1(n318), .A2(n602), .B1(\unit_memory/DRAM/n3121 ), .B2(
        n607), .ZN(\unit_memory/DRAM/n1426 ) );
  OAI22_X1 U3284 ( .A1(n321), .A2(n602), .B1(\unit_memory/DRAM/n3122 ), .B2(
        n607), .ZN(\unit_memory/DRAM/n1425 ) );
  OAI22_X1 U3285 ( .A1(n324), .A2(n601), .B1(\unit_memory/DRAM/n3123 ), .B2(
        n608), .ZN(\unit_memory/DRAM/n1424 ) );
  OAI22_X1 U3286 ( .A1(n327), .A2(n601), .B1(\unit_memory/DRAM/n3124 ), .B2(
        n608), .ZN(\unit_memory/DRAM/n1423 ) );
  OAI22_X1 U3287 ( .A1(n330), .A2(n601), .B1(\unit_memory/DRAM/n3125 ), .B2(
        n608), .ZN(\unit_memory/DRAM/n1422 ) );
  OAI22_X1 U3288 ( .A1(n333), .A2(n601), .B1(\unit_memory/DRAM/n3126 ), .B2(
        n608), .ZN(\unit_memory/DRAM/n1421 ) );
  OAI22_X1 U3289 ( .A1(n336), .A2(n601), .B1(\unit_memory/DRAM/n3127 ), .B2(
        n609), .ZN(\unit_memory/DRAM/n1420 ) );
  OAI22_X1 U3290 ( .A1(n339), .A2(n601), .B1(\unit_memory/DRAM/n3128 ), .B2(
        n609), .ZN(\unit_memory/DRAM/n1419 ) );
  OAI22_X1 U3291 ( .A1(n342), .A2(n601), .B1(\unit_memory/DRAM/n3129 ), .B2(
        n609), .ZN(\unit_memory/DRAM/n1418 ) );
  OAI22_X1 U3292 ( .A1(n345), .A2(n601), .B1(\unit_memory/DRAM/n3130 ), .B2(
        n609), .ZN(\unit_memory/DRAM/n1417 ) );
  OAI22_X1 U3293 ( .A1(n348), .A2(n601), .B1(\unit_memory/DRAM/n3131 ), .B2(
        n610), .ZN(\unit_memory/DRAM/n1416 ) );
  OAI22_X1 U3294 ( .A1(n351), .A2(n601), .B1(\unit_memory/DRAM/n3132 ), .B2(
        n610), .ZN(\unit_memory/DRAM/n1415 ) );
  OAI22_X1 U3295 ( .A1(n354), .A2(n601), .B1(\unit_memory/DRAM/n3133 ), .B2(
        n610), .ZN(\unit_memory/DRAM/n1414 ) );
  OAI22_X1 U3296 ( .A1(n357), .A2(n601), .B1(\unit_memory/DRAM/n3134 ), .B2(
        n610), .ZN(\unit_memory/DRAM/n1413 ) );
  OAI22_X1 U3297 ( .A1(n289), .A2(n613), .B1(\unit_memory/DRAM/n3143 ), .B2(
        n616), .ZN(\unit_memory/DRAM/n1404 ) );
  OAI22_X1 U3298 ( .A1(n292), .A2(n613), .B1(\unit_memory/DRAM/n3144 ), .B2(
        n616), .ZN(\unit_memory/DRAM/n1403 ) );
  OAI22_X1 U3299 ( .A1(n295), .A2(n613), .B1(\unit_memory/DRAM/n3145 ), .B2(
        n616), .ZN(\unit_memory/DRAM/n1402 ) );
  OAI22_X1 U3300 ( .A1(n298), .A2(n613), .B1(\unit_memory/DRAM/n3146 ), .B2(
        n616), .ZN(\unit_memory/DRAM/n1401 ) );
  OAI22_X1 U3301 ( .A1(n301), .A2(n613), .B1(\unit_memory/DRAM/n3147 ), .B2(
        n617), .ZN(\unit_memory/DRAM/n1400 ) );
  OAI22_X1 U3302 ( .A1(n304), .A2(n613), .B1(\unit_memory/DRAM/n3148 ), .B2(
        n617), .ZN(\unit_memory/DRAM/n1399 ) );
  OAI22_X1 U3303 ( .A1(n307), .A2(n613), .B1(\unit_memory/DRAM/n3149 ), .B2(
        n617), .ZN(\unit_memory/DRAM/n1398 ) );
  OAI22_X1 U3304 ( .A1(n310), .A2(n613), .B1(\unit_memory/DRAM/n3150 ), .B2(
        n617), .ZN(\unit_memory/DRAM/n1397 ) );
  OAI22_X1 U3305 ( .A1(n313), .A2(n613), .B1(\unit_memory/DRAM/n3151 ), .B2(
        n618), .ZN(\unit_memory/DRAM/n1396 ) );
  OAI22_X1 U3306 ( .A1(n316), .A2(n613), .B1(\unit_memory/DRAM/n3152 ), .B2(
        n618), .ZN(\unit_memory/DRAM/n1395 ) );
  OAI22_X1 U3307 ( .A1(n319), .A2(n613), .B1(\unit_memory/DRAM/n3153 ), .B2(
        n618), .ZN(\unit_memory/DRAM/n1394 ) );
  OAI22_X1 U3308 ( .A1(n322), .A2(n613), .B1(\unit_memory/DRAM/n3154 ), .B2(
        n618), .ZN(\unit_memory/DRAM/n1393 ) );
  OAI22_X1 U3309 ( .A1(n325), .A2(n612), .B1(\unit_memory/DRAM/n3155 ), .B2(
        n619), .ZN(\unit_memory/DRAM/n1392 ) );
  OAI22_X1 U3310 ( .A1(n328), .A2(n612), .B1(\unit_memory/DRAM/n3156 ), .B2(
        n619), .ZN(\unit_memory/DRAM/n1391 ) );
  OAI22_X1 U3311 ( .A1(n331), .A2(n612), .B1(\unit_memory/DRAM/n3157 ), .B2(
        n619), .ZN(\unit_memory/DRAM/n1390 ) );
  OAI22_X1 U3312 ( .A1(n334), .A2(n612), .B1(\unit_memory/DRAM/n3158 ), .B2(
        n619), .ZN(\unit_memory/DRAM/n1389 ) );
  OAI22_X1 U3313 ( .A1(n337), .A2(n612), .B1(\unit_memory/DRAM/n3159 ), .B2(
        n620), .ZN(\unit_memory/DRAM/n1388 ) );
  OAI22_X1 U3314 ( .A1(n340), .A2(n612), .B1(\unit_memory/DRAM/n3160 ), .B2(
        n620), .ZN(\unit_memory/DRAM/n1387 ) );
  OAI22_X1 U3315 ( .A1(n343), .A2(n612), .B1(\unit_memory/DRAM/n3161 ), .B2(
        n620), .ZN(\unit_memory/DRAM/n1386 ) );
  OAI22_X1 U3316 ( .A1(n346), .A2(n612), .B1(\unit_memory/DRAM/n3162 ), .B2(
        n620), .ZN(\unit_memory/DRAM/n1385 ) );
  OAI22_X1 U3317 ( .A1(n349), .A2(n612), .B1(\unit_memory/DRAM/n3163 ), .B2(
        n621), .ZN(\unit_memory/DRAM/n1384 ) );
  OAI22_X1 U3318 ( .A1(n352), .A2(n612), .B1(\unit_memory/DRAM/n3164 ), .B2(
        n621), .ZN(\unit_memory/DRAM/n1383 ) );
  OAI22_X1 U3319 ( .A1(n355), .A2(n612), .B1(\unit_memory/DRAM/n3165 ), .B2(
        n621), .ZN(\unit_memory/DRAM/n1382 ) );
  OAI22_X1 U3320 ( .A1(n357), .A2(n612), .B1(\unit_memory/DRAM/n3166 ), .B2(
        n621), .ZN(\unit_memory/DRAM/n1381 ) );
  OAI22_X1 U3321 ( .A1(n249), .A2(n635), .B1(\unit_memory/DRAM/n3199 ), .B2(
        n636), .ZN(\unit_memory/DRAM/n1348 ) );
  OAI22_X1 U3322 ( .A1(n268), .A2(n634), .B1(\unit_memory/DRAM/n3200 ), .B2(
        n636), .ZN(\unit_memory/DRAM/n1347 ) );
  OAI22_X1 U3323 ( .A1(n271), .A2(n635), .B1(\unit_memory/DRAM/n3201 ), .B2(
        n636), .ZN(\unit_memory/DRAM/n1346 ) );
  OAI22_X1 U3324 ( .A1(n274), .A2(n634), .B1(\unit_memory/DRAM/n3202 ), .B2(
        n636), .ZN(\unit_memory/DRAM/n1345 ) );
  OAI22_X1 U3325 ( .A1(n277), .A2(n635), .B1(\unit_memory/DRAM/n3203 ), .B2(
        n637), .ZN(\unit_memory/DRAM/n1344 ) );
  OAI22_X1 U3326 ( .A1(n280), .A2(n634), .B1(\unit_memory/DRAM/n3204 ), .B2(
        n637), .ZN(\unit_memory/DRAM/n1343 ) );
  OAI22_X1 U3327 ( .A1(n283), .A2(n635), .B1(\unit_memory/DRAM/n3205 ), .B2(
        n637), .ZN(\unit_memory/DRAM/n1342 ) );
  OAI22_X1 U3328 ( .A1(n286), .A2(n634), .B1(\unit_memory/DRAM/n3206 ), .B2(
        n637), .ZN(\unit_memory/DRAM/n1341 ) );
  OAI22_X1 U3329 ( .A1(n289), .A2(n635), .B1(\unit_memory/DRAM/n3207 ), .B2(
        n638), .ZN(\unit_memory/DRAM/n1340 ) );
  OAI22_X1 U3330 ( .A1(n292), .A2(n635), .B1(\unit_memory/DRAM/n3208 ), .B2(
        n638), .ZN(\unit_memory/DRAM/n1339 ) );
  OAI22_X1 U3331 ( .A1(n295), .A2(n635), .B1(\unit_memory/DRAM/n3209 ), .B2(
        n638), .ZN(\unit_memory/DRAM/n1338 ) );
  OAI22_X1 U3332 ( .A1(n298), .A2(n635), .B1(\unit_memory/DRAM/n3210 ), .B2(
        n638), .ZN(\unit_memory/DRAM/n1337 ) );
  OAI22_X1 U3333 ( .A1(n301), .A2(n635), .B1(\unit_memory/DRAM/n3211 ), .B2(
        n639), .ZN(\unit_memory/DRAM/n1336 ) );
  OAI22_X1 U3334 ( .A1(n304), .A2(n635), .B1(\unit_memory/DRAM/n3212 ), .B2(
        n639), .ZN(\unit_memory/DRAM/n1335 ) );
  OAI22_X1 U3335 ( .A1(n307), .A2(n635), .B1(\unit_memory/DRAM/n3213 ), .B2(
        n639), .ZN(\unit_memory/DRAM/n1334 ) );
  OAI22_X1 U3336 ( .A1(n310), .A2(n635), .B1(\unit_memory/DRAM/n3214 ), .B2(
        n639), .ZN(\unit_memory/DRAM/n1333 ) );
  OAI22_X1 U3337 ( .A1(n313), .A2(n635), .B1(\unit_memory/DRAM/n3215 ), .B2(
        n640), .ZN(\unit_memory/DRAM/n1332 ) );
  OAI22_X1 U3338 ( .A1(n316), .A2(n635), .B1(\unit_memory/DRAM/n3216 ), .B2(
        n640), .ZN(\unit_memory/DRAM/n1331 ) );
  OAI22_X1 U3339 ( .A1(n319), .A2(n635), .B1(\unit_memory/DRAM/n3217 ), .B2(
        n640), .ZN(\unit_memory/DRAM/n1330 ) );
  OAI22_X1 U3340 ( .A1(n322), .A2(n635), .B1(\unit_memory/DRAM/n3218 ), .B2(
        n640), .ZN(\unit_memory/DRAM/n1329 ) );
  OAI22_X1 U3341 ( .A1(n325), .A2(n634), .B1(\unit_memory/DRAM/n3219 ), .B2(
        n641), .ZN(\unit_memory/DRAM/n1328 ) );
  OAI22_X1 U3342 ( .A1(n328), .A2(n634), .B1(\unit_memory/DRAM/n3220 ), .B2(
        n641), .ZN(\unit_memory/DRAM/n1327 ) );
  OAI22_X1 U3343 ( .A1(n331), .A2(n634), .B1(\unit_memory/DRAM/n3221 ), .B2(
        n641), .ZN(\unit_memory/DRAM/n1326 ) );
  OAI22_X1 U3344 ( .A1(n334), .A2(n634), .B1(\unit_memory/DRAM/n3222 ), .B2(
        n641), .ZN(\unit_memory/DRAM/n1325 ) );
  OAI22_X1 U3345 ( .A1(n337), .A2(n634), .B1(\unit_memory/DRAM/n3223 ), .B2(
        n642), .ZN(\unit_memory/DRAM/n1324 ) );
  OAI22_X1 U3346 ( .A1(n340), .A2(n634), .B1(\unit_memory/DRAM/n3224 ), .B2(
        n642), .ZN(\unit_memory/DRAM/n1323 ) );
  OAI22_X1 U3347 ( .A1(n343), .A2(n634), .B1(\unit_memory/DRAM/n3225 ), .B2(
        n642), .ZN(\unit_memory/DRAM/n1322 ) );
  OAI22_X1 U3348 ( .A1(n346), .A2(n634), .B1(\unit_memory/DRAM/n3226 ), .B2(
        n642), .ZN(\unit_memory/DRAM/n1321 ) );
  OAI22_X1 U3349 ( .A1(n349), .A2(n634), .B1(\unit_memory/DRAM/n3227 ), .B2(
        n643), .ZN(\unit_memory/DRAM/n1320 ) );
  OAI22_X1 U3350 ( .A1(n352), .A2(n634), .B1(\unit_memory/DRAM/n3228 ), .B2(
        n643), .ZN(\unit_memory/DRAM/n1319 ) );
  OAI22_X1 U3351 ( .A1(n355), .A2(n634), .B1(\unit_memory/DRAM/n3229 ), .B2(
        n643), .ZN(\unit_memory/DRAM/n1318 ) );
  OAI22_X1 U3352 ( .A1(n358), .A2(n634), .B1(\unit_memory/DRAM/n3230 ), .B2(
        n643), .ZN(\unit_memory/DRAM/n1317 ) );
  OAI22_X1 U3353 ( .A1(n249), .A2(n646), .B1(\unit_memory/DRAM/n3231 ), .B2(
        n647), .ZN(\unit_memory/DRAM/n1316 ) );
  OAI22_X1 U3354 ( .A1(n268), .A2(n645), .B1(\unit_memory/DRAM/n3232 ), .B2(
        n647), .ZN(\unit_memory/DRAM/n1315 ) );
  OAI22_X1 U3355 ( .A1(n271), .A2(n646), .B1(\unit_memory/DRAM/n3233 ), .B2(
        n647), .ZN(\unit_memory/DRAM/n1314 ) );
  OAI22_X1 U3356 ( .A1(n274), .A2(n645), .B1(\unit_memory/DRAM/n3234 ), .B2(
        n647), .ZN(\unit_memory/DRAM/n1313 ) );
  OAI22_X1 U3357 ( .A1(n277), .A2(n646), .B1(\unit_memory/DRAM/n3235 ), .B2(
        n648), .ZN(\unit_memory/DRAM/n1312 ) );
  OAI22_X1 U3358 ( .A1(n280), .A2(n645), .B1(\unit_memory/DRAM/n3236 ), .B2(
        n648), .ZN(\unit_memory/DRAM/n1311 ) );
  OAI22_X1 U3359 ( .A1(n283), .A2(n646), .B1(\unit_memory/DRAM/n3237 ), .B2(
        n648), .ZN(\unit_memory/DRAM/n1310 ) );
  OAI22_X1 U3360 ( .A1(n286), .A2(n645), .B1(\unit_memory/DRAM/n3238 ), .B2(
        n648), .ZN(\unit_memory/DRAM/n1309 ) );
  OAI22_X1 U3361 ( .A1(n289), .A2(n646), .B1(\unit_memory/DRAM/n3239 ), .B2(
        n649), .ZN(\unit_memory/DRAM/n1308 ) );
  OAI22_X1 U3362 ( .A1(n292), .A2(n646), .B1(\unit_memory/DRAM/n3240 ), .B2(
        n649), .ZN(\unit_memory/DRAM/n1307 ) );
  OAI22_X1 U3363 ( .A1(n295), .A2(n646), .B1(\unit_memory/DRAM/n3241 ), .B2(
        n649), .ZN(\unit_memory/DRAM/n1306 ) );
  OAI22_X1 U3364 ( .A1(n298), .A2(n646), .B1(\unit_memory/DRAM/n3242 ), .B2(
        n649), .ZN(\unit_memory/DRAM/n1305 ) );
  OAI22_X1 U3365 ( .A1(n301), .A2(n646), .B1(\unit_memory/DRAM/n3243 ), .B2(
        n650), .ZN(\unit_memory/DRAM/n1304 ) );
  OAI22_X1 U3366 ( .A1(n304), .A2(n646), .B1(\unit_memory/DRAM/n3244 ), .B2(
        n650), .ZN(\unit_memory/DRAM/n1303 ) );
  OAI22_X1 U3367 ( .A1(n307), .A2(n646), .B1(\unit_memory/DRAM/n3245 ), .B2(
        n650), .ZN(\unit_memory/DRAM/n1302 ) );
  OAI22_X1 U3368 ( .A1(n310), .A2(n646), .B1(\unit_memory/DRAM/n3246 ), .B2(
        n650), .ZN(\unit_memory/DRAM/n1301 ) );
  OAI22_X1 U3369 ( .A1(n313), .A2(n646), .B1(\unit_memory/DRAM/n3247 ), .B2(
        n651), .ZN(\unit_memory/DRAM/n1300 ) );
  OAI22_X1 U3370 ( .A1(n316), .A2(n646), .B1(\unit_memory/DRAM/n3248 ), .B2(
        n651), .ZN(\unit_memory/DRAM/n1299 ) );
  OAI22_X1 U3371 ( .A1(n319), .A2(n646), .B1(\unit_memory/DRAM/n3249 ), .B2(
        n651), .ZN(\unit_memory/DRAM/n1298 ) );
  OAI22_X1 U3372 ( .A1(n322), .A2(n646), .B1(\unit_memory/DRAM/n3250 ), .B2(
        n651), .ZN(\unit_memory/DRAM/n1297 ) );
  OAI22_X1 U3373 ( .A1(n325), .A2(n645), .B1(\unit_memory/DRAM/n3251 ), .B2(
        n652), .ZN(\unit_memory/DRAM/n1296 ) );
  OAI22_X1 U3374 ( .A1(n328), .A2(n645), .B1(\unit_memory/DRAM/n3252 ), .B2(
        n652), .ZN(\unit_memory/DRAM/n1295 ) );
  OAI22_X1 U3375 ( .A1(n331), .A2(n645), .B1(\unit_memory/DRAM/n3253 ), .B2(
        n652), .ZN(\unit_memory/DRAM/n1294 ) );
  OAI22_X1 U3376 ( .A1(n334), .A2(n645), .B1(\unit_memory/DRAM/n3254 ), .B2(
        n652), .ZN(\unit_memory/DRAM/n1293 ) );
  OAI22_X1 U3377 ( .A1(n337), .A2(n645), .B1(\unit_memory/DRAM/n3255 ), .B2(
        n653), .ZN(\unit_memory/DRAM/n1292 ) );
  OAI22_X1 U3378 ( .A1(n340), .A2(n645), .B1(\unit_memory/DRAM/n3256 ), .B2(
        n653), .ZN(\unit_memory/DRAM/n1291 ) );
  OAI22_X1 U3379 ( .A1(n343), .A2(n645), .B1(\unit_memory/DRAM/n3257 ), .B2(
        n653), .ZN(\unit_memory/DRAM/n1290 ) );
  OAI22_X1 U3380 ( .A1(n346), .A2(n645), .B1(\unit_memory/DRAM/n3258 ), .B2(
        n653), .ZN(\unit_memory/DRAM/n1289 ) );
  OAI22_X1 U3381 ( .A1(n349), .A2(n645), .B1(\unit_memory/DRAM/n3259 ), .B2(
        n654), .ZN(\unit_memory/DRAM/n1288 ) );
  OAI22_X1 U3382 ( .A1(n352), .A2(n645), .B1(\unit_memory/DRAM/n3260 ), .B2(
        n654), .ZN(\unit_memory/DRAM/n1287 ) );
  OAI22_X1 U3383 ( .A1(n355), .A2(n645), .B1(\unit_memory/DRAM/n3261 ), .B2(
        n654), .ZN(\unit_memory/DRAM/n1286 ) );
  OAI22_X1 U3384 ( .A1(n358), .A2(n645), .B1(\unit_memory/DRAM/n3262 ), .B2(
        n654), .ZN(\unit_memory/DRAM/n1285 ) );
  OAI22_X1 U3385 ( .A1(n289), .A2(n657), .B1(\unit_memory/DRAM/n3271 ), .B2(
        n660), .ZN(\unit_memory/DRAM/n1276 ) );
  OAI22_X1 U3386 ( .A1(n292), .A2(n657), .B1(\unit_memory/DRAM/n3272 ), .B2(
        n660), .ZN(\unit_memory/DRAM/n1275 ) );
  OAI22_X1 U3387 ( .A1(n295), .A2(n657), .B1(\unit_memory/DRAM/n3273 ), .B2(
        n660), .ZN(\unit_memory/DRAM/n1274 ) );
  OAI22_X1 U3388 ( .A1(n298), .A2(n657), .B1(\unit_memory/DRAM/n3274 ), .B2(
        n660), .ZN(\unit_memory/DRAM/n1273 ) );
  OAI22_X1 U3389 ( .A1(n301), .A2(n657), .B1(\unit_memory/DRAM/n3275 ), .B2(
        n661), .ZN(\unit_memory/DRAM/n1272 ) );
  OAI22_X1 U3390 ( .A1(n304), .A2(n657), .B1(\unit_memory/DRAM/n3276 ), .B2(
        n661), .ZN(\unit_memory/DRAM/n1271 ) );
  OAI22_X1 U3391 ( .A1(n307), .A2(n657), .B1(\unit_memory/DRAM/n3277 ), .B2(
        n661), .ZN(\unit_memory/DRAM/n1270 ) );
  OAI22_X1 U3392 ( .A1(n310), .A2(n657), .B1(\unit_memory/DRAM/n3278 ), .B2(
        n661), .ZN(\unit_memory/DRAM/n1269 ) );
  OAI22_X1 U3393 ( .A1(n313), .A2(n657), .B1(\unit_memory/DRAM/n3279 ), .B2(
        n662), .ZN(\unit_memory/DRAM/n1268 ) );
  OAI22_X1 U3394 ( .A1(n316), .A2(n657), .B1(\unit_memory/DRAM/n3280 ), .B2(
        n662), .ZN(\unit_memory/DRAM/n1267 ) );
  OAI22_X1 U3395 ( .A1(n319), .A2(n657), .B1(\unit_memory/DRAM/n3281 ), .B2(
        n662), .ZN(\unit_memory/DRAM/n1266 ) );
  OAI22_X1 U3396 ( .A1(n322), .A2(n657), .B1(\unit_memory/DRAM/n3282 ), .B2(
        n662), .ZN(\unit_memory/DRAM/n1265 ) );
  OAI22_X1 U3397 ( .A1(n325), .A2(n656), .B1(\unit_memory/DRAM/n3283 ), .B2(
        n663), .ZN(\unit_memory/DRAM/n1264 ) );
  OAI22_X1 U3398 ( .A1(n328), .A2(n656), .B1(\unit_memory/DRAM/n3284 ), .B2(
        n663), .ZN(\unit_memory/DRAM/n1263 ) );
  OAI22_X1 U3399 ( .A1(n331), .A2(n656), .B1(\unit_memory/DRAM/n3285 ), .B2(
        n663), .ZN(\unit_memory/DRAM/n1262 ) );
  OAI22_X1 U3400 ( .A1(n334), .A2(n656), .B1(\unit_memory/DRAM/n3286 ), .B2(
        n663), .ZN(\unit_memory/DRAM/n1261 ) );
  OAI22_X1 U3401 ( .A1(n337), .A2(n656), .B1(\unit_memory/DRAM/n3287 ), .B2(
        n664), .ZN(\unit_memory/DRAM/n1260 ) );
  OAI22_X1 U3402 ( .A1(n340), .A2(n656), .B1(\unit_memory/DRAM/n3288 ), .B2(
        n664), .ZN(\unit_memory/DRAM/n1259 ) );
  OAI22_X1 U3403 ( .A1(n343), .A2(n656), .B1(\unit_memory/DRAM/n3289 ), .B2(
        n664), .ZN(\unit_memory/DRAM/n1258 ) );
  OAI22_X1 U3404 ( .A1(n346), .A2(n656), .B1(\unit_memory/DRAM/n3290 ), .B2(
        n664), .ZN(\unit_memory/DRAM/n1257 ) );
  OAI22_X1 U3405 ( .A1(n349), .A2(n656), .B1(\unit_memory/DRAM/n3291 ), .B2(
        n665), .ZN(\unit_memory/DRAM/n1256 ) );
  OAI22_X1 U3406 ( .A1(n352), .A2(n656), .B1(\unit_memory/DRAM/n3292 ), .B2(
        n665), .ZN(\unit_memory/DRAM/n1255 ) );
  OAI22_X1 U3407 ( .A1(n355), .A2(n656), .B1(\unit_memory/DRAM/n3293 ), .B2(
        n665), .ZN(\unit_memory/DRAM/n1254 ) );
  OAI22_X1 U3408 ( .A1(n358), .A2(n656), .B1(\unit_memory/DRAM/n3294 ), .B2(
        n665), .ZN(\unit_memory/DRAM/n1253 ) );
  OAI22_X1 U3409 ( .A1(n249), .A2(n679), .B1(\unit_memory/DRAM/n3327 ), .B2(
        n680), .ZN(\unit_memory/DRAM/n1220 ) );
  OAI22_X1 U3410 ( .A1(n266), .A2(n678), .B1(\unit_memory/DRAM/n3328 ), .B2(
        n680), .ZN(\unit_memory/DRAM/n1219 ) );
  OAI22_X1 U3411 ( .A1(n269), .A2(n679), .B1(\unit_memory/DRAM/n3329 ), .B2(
        n680), .ZN(\unit_memory/DRAM/n1218 ) );
  OAI22_X1 U3412 ( .A1(n272), .A2(n678), .B1(\unit_memory/DRAM/n3330 ), .B2(
        n680), .ZN(\unit_memory/DRAM/n1217 ) );
  OAI22_X1 U3413 ( .A1(n275), .A2(n679), .B1(\unit_memory/DRAM/n3331 ), .B2(
        n681), .ZN(\unit_memory/DRAM/n1216 ) );
  OAI22_X1 U3414 ( .A1(n278), .A2(n678), .B1(\unit_memory/DRAM/n3332 ), .B2(
        n681), .ZN(\unit_memory/DRAM/n1215 ) );
  OAI22_X1 U3415 ( .A1(n281), .A2(n679), .B1(\unit_memory/DRAM/n3333 ), .B2(
        n681), .ZN(\unit_memory/DRAM/n1214 ) );
  OAI22_X1 U3416 ( .A1(n284), .A2(n678), .B1(\unit_memory/DRAM/n3334 ), .B2(
        n681), .ZN(\unit_memory/DRAM/n1213 ) );
  OAI22_X1 U3417 ( .A1(n287), .A2(n679), .B1(\unit_memory/DRAM/n3335 ), .B2(
        n682), .ZN(\unit_memory/DRAM/n1212 ) );
  OAI22_X1 U3418 ( .A1(n290), .A2(n679), .B1(\unit_memory/DRAM/n3336 ), .B2(
        n682), .ZN(\unit_memory/DRAM/n1211 ) );
  OAI22_X1 U3419 ( .A1(n293), .A2(n679), .B1(\unit_memory/DRAM/n3337 ), .B2(
        n682), .ZN(\unit_memory/DRAM/n1210 ) );
  OAI22_X1 U3420 ( .A1(n296), .A2(n679), .B1(\unit_memory/DRAM/n3338 ), .B2(
        n682), .ZN(\unit_memory/DRAM/n1209 ) );
  OAI22_X1 U3421 ( .A1(n299), .A2(n679), .B1(\unit_memory/DRAM/n3339 ), .B2(
        n683), .ZN(\unit_memory/DRAM/n1208 ) );
  OAI22_X1 U3422 ( .A1(n302), .A2(n679), .B1(\unit_memory/DRAM/n3340 ), .B2(
        n683), .ZN(\unit_memory/DRAM/n1207 ) );
  OAI22_X1 U3423 ( .A1(n305), .A2(n679), .B1(\unit_memory/DRAM/n3341 ), .B2(
        n683), .ZN(\unit_memory/DRAM/n1206 ) );
  OAI22_X1 U3424 ( .A1(n308), .A2(n679), .B1(\unit_memory/DRAM/n3342 ), .B2(
        n683), .ZN(\unit_memory/DRAM/n1205 ) );
  OAI22_X1 U3425 ( .A1(n311), .A2(n679), .B1(\unit_memory/DRAM/n3343 ), .B2(
        n684), .ZN(\unit_memory/DRAM/n1204 ) );
  OAI22_X1 U3426 ( .A1(n314), .A2(n679), .B1(\unit_memory/DRAM/n3344 ), .B2(
        n684), .ZN(\unit_memory/DRAM/n1203 ) );
  OAI22_X1 U3427 ( .A1(n317), .A2(n679), .B1(\unit_memory/DRAM/n3345 ), .B2(
        n684), .ZN(\unit_memory/DRAM/n1202 ) );
  OAI22_X1 U3428 ( .A1(n320), .A2(n679), .B1(\unit_memory/DRAM/n3346 ), .B2(
        n684), .ZN(\unit_memory/DRAM/n1201 ) );
  OAI22_X1 U3429 ( .A1(n323), .A2(n678), .B1(\unit_memory/DRAM/n3347 ), .B2(
        n685), .ZN(\unit_memory/DRAM/n1200 ) );
  OAI22_X1 U3430 ( .A1(n326), .A2(n678), .B1(\unit_memory/DRAM/n3348 ), .B2(
        n685), .ZN(\unit_memory/DRAM/n1199 ) );
  OAI22_X1 U3431 ( .A1(n329), .A2(n678), .B1(\unit_memory/DRAM/n3349 ), .B2(
        n685), .ZN(\unit_memory/DRAM/n1198 ) );
  OAI22_X1 U3432 ( .A1(n332), .A2(n678), .B1(\unit_memory/DRAM/n3350 ), .B2(
        n685), .ZN(\unit_memory/DRAM/n1197 ) );
  OAI22_X1 U3433 ( .A1(n335), .A2(n678), .B1(\unit_memory/DRAM/n3351 ), .B2(
        n686), .ZN(\unit_memory/DRAM/n1196 ) );
  OAI22_X1 U3434 ( .A1(n338), .A2(n678), .B1(\unit_memory/DRAM/n3352 ), .B2(
        n686), .ZN(\unit_memory/DRAM/n1195 ) );
  OAI22_X1 U3435 ( .A1(n341), .A2(n678), .B1(\unit_memory/DRAM/n3353 ), .B2(
        n686), .ZN(\unit_memory/DRAM/n1194 ) );
  OAI22_X1 U3436 ( .A1(n344), .A2(n678), .B1(\unit_memory/DRAM/n3354 ), .B2(
        n686), .ZN(\unit_memory/DRAM/n1193 ) );
  OAI22_X1 U3437 ( .A1(n347), .A2(n678), .B1(\unit_memory/DRAM/n3355 ), .B2(
        n687), .ZN(\unit_memory/DRAM/n1192 ) );
  OAI22_X1 U3438 ( .A1(n350), .A2(n678), .B1(\unit_memory/DRAM/n3356 ), .B2(
        n687), .ZN(\unit_memory/DRAM/n1191 ) );
  OAI22_X1 U3439 ( .A1(n353), .A2(n678), .B1(\unit_memory/DRAM/n3357 ), .B2(
        n687), .ZN(\unit_memory/DRAM/n1190 ) );
  OAI22_X1 U3440 ( .A1(n358), .A2(n678), .B1(\unit_memory/DRAM/n3358 ), .B2(
        n687), .ZN(\unit_memory/DRAM/n1189 ) );
  OAI22_X1 U3441 ( .A1(n314), .A2(n360), .B1(\unit_memory/DRAM/n2416 ), .B2(
        n365), .ZN(\unit_memory/DRAM/n2131 ) );
  OAI22_X1 U3442 ( .A1(n317), .A2(n360), .B1(\unit_memory/DRAM/n2417 ), .B2(
        n365), .ZN(\unit_memory/DRAM/n2130 ) );
  OAI22_X1 U3443 ( .A1(n320), .A2(n360), .B1(\unit_memory/DRAM/n2418 ), .B2(
        n365), .ZN(\unit_memory/DRAM/n2129 ) );
  OAI22_X1 U3444 ( .A1(n323), .A2(n359), .B1(\unit_memory/DRAM/n2419 ), .B2(
        n366), .ZN(\unit_memory/DRAM/n2128 ) );
  OAI22_X1 U3445 ( .A1(n326), .A2(n359), .B1(\unit_memory/DRAM/n2420 ), .B2(
        n366), .ZN(\unit_memory/DRAM/n2127 ) );
  OAI22_X1 U3446 ( .A1(n329), .A2(n359), .B1(\unit_memory/DRAM/n2421 ), .B2(
        n366), .ZN(\unit_memory/DRAM/n2126 ) );
  OAI22_X1 U3447 ( .A1(n332), .A2(n359), .B1(\unit_memory/DRAM/n2422 ), .B2(
        n366), .ZN(\unit_memory/DRAM/n2125 ) );
  OAI22_X1 U3448 ( .A1(n338), .A2(n359), .B1(\unit_memory/DRAM/n2424 ), .B2(
        n367), .ZN(\unit_memory/DRAM/n2123 ) );
  OAI22_X1 U3449 ( .A1(n341), .A2(n359), .B1(\unit_memory/DRAM/n2425 ), .B2(
        n367), .ZN(\unit_memory/DRAM/n2122 ) );
  OAI22_X1 U3450 ( .A1(n344), .A2(n359), .B1(\unit_memory/DRAM/n2426 ), .B2(
        n367), .ZN(\unit_memory/DRAM/n2121 ) );
  OAI22_X1 U3451 ( .A1(n347), .A2(n359), .B1(\unit_memory/DRAM/n2427 ), .B2(
        n368), .ZN(\unit_memory/DRAM/n2120 ) );
  OAI22_X1 U3452 ( .A1(n350), .A2(n359), .B1(\unit_memory/DRAM/n2428 ), .B2(
        n368), .ZN(\unit_memory/DRAM/n2119 ) );
  OAI22_X1 U3453 ( .A1(n353), .A2(n359), .B1(\unit_memory/DRAM/n2429 ), .B2(
        n368), .ZN(\unit_memory/DRAM/n2118 ) );
  OAI22_X1 U3454 ( .A1(n356), .A2(n359), .B1(\unit_memory/DRAM/n2430 ), .B2(
        n368), .ZN(\unit_memory/DRAM/n2117 ) );
  OAI22_X1 U3455 ( .A1(n314), .A2(n404), .B1(\unit_memory/DRAM/n2544 ), .B2(
        n409), .ZN(\unit_memory/DRAM/n2003 ) );
  OAI22_X1 U3456 ( .A1(n317), .A2(n404), .B1(\unit_memory/DRAM/n2545 ), .B2(
        n409), .ZN(\unit_memory/DRAM/n2002 ) );
  OAI22_X1 U3457 ( .A1(n320), .A2(n404), .B1(\unit_memory/DRAM/n2546 ), .B2(
        n409), .ZN(\unit_memory/DRAM/n2001 ) );
  OAI22_X1 U3458 ( .A1(n323), .A2(n403), .B1(\unit_memory/DRAM/n2547 ), .B2(
        n410), .ZN(\unit_memory/DRAM/n2000 ) );
  OAI22_X1 U3459 ( .A1(n326), .A2(n403), .B1(\unit_memory/DRAM/n2548 ), .B2(
        n410), .ZN(\unit_memory/DRAM/n1999 ) );
  OAI22_X1 U3460 ( .A1(n329), .A2(n403), .B1(\unit_memory/DRAM/n2549 ), .B2(
        n410), .ZN(\unit_memory/DRAM/n1998 ) );
  OAI22_X1 U3461 ( .A1(n332), .A2(n403), .B1(\unit_memory/DRAM/n2550 ), .B2(
        n410), .ZN(\unit_memory/DRAM/n1997 ) );
  OAI22_X1 U3462 ( .A1(n338), .A2(n403), .B1(\unit_memory/DRAM/n2552 ), .B2(
        n411), .ZN(\unit_memory/DRAM/n1995 ) );
  OAI22_X1 U3463 ( .A1(n341), .A2(n403), .B1(\unit_memory/DRAM/n2553 ), .B2(
        n411), .ZN(\unit_memory/DRAM/n1994 ) );
  OAI22_X1 U3464 ( .A1(n344), .A2(n403), .B1(\unit_memory/DRAM/n2554 ), .B2(
        n411), .ZN(\unit_memory/DRAM/n1993 ) );
  OAI22_X1 U3465 ( .A1(n347), .A2(n403), .B1(\unit_memory/DRAM/n2555 ), .B2(
        n412), .ZN(\unit_memory/DRAM/n1992 ) );
  OAI22_X1 U3466 ( .A1(n350), .A2(n403), .B1(\unit_memory/DRAM/n2556 ), .B2(
        n412), .ZN(\unit_memory/DRAM/n1991 ) );
  OAI22_X1 U3467 ( .A1(n353), .A2(n403), .B1(\unit_memory/DRAM/n2557 ), .B2(
        n412), .ZN(\unit_memory/DRAM/n1990 ) );
  OAI22_X1 U3468 ( .A1(n356), .A2(n403), .B1(\unit_memory/DRAM/n2558 ), .B2(
        n412), .ZN(\unit_memory/DRAM/n1989 ) );
  OAI22_X1 U3469 ( .A1(n261), .A2(n314), .B1(\unit_memory/DRAM/n2384 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2163 ) );
  OAI22_X1 U3470 ( .A1(n261), .A2(n317), .B1(\unit_memory/DRAM/n2385 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2162 ) );
  OAI22_X1 U3471 ( .A1(n261), .A2(n320), .B1(\unit_memory/DRAM/n2386 ), .B2(
        n256), .ZN(\unit_memory/DRAM/n2161 ) );
  OAI22_X1 U3472 ( .A1(n262), .A2(n323), .B1(\unit_memory/DRAM/n2387 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2160 ) );
  OAI22_X1 U3473 ( .A1(n262), .A2(n326), .B1(\unit_memory/DRAM/n2388 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2159 ) );
  OAI22_X1 U3474 ( .A1(n262), .A2(n329), .B1(\unit_memory/DRAM/n2389 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2158 ) );
  OAI22_X1 U3475 ( .A1(n262), .A2(n332), .B1(\unit_memory/DRAM/n2390 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2157 ) );
  OAI22_X1 U3476 ( .A1(n263), .A2(n338), .B1(\unit_memory/DRAM/n2392 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2155 ) );
  OAI22_X1 U3477 ( .A1(n263), .A2(n341), .B1(\unit_memory/DRAM/n2393 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2154 ) );
  OAI22_X1 U3478 ( .A1(n263), .A2(n344), .B1(\unit_memory/DRAM/n2394 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2153 ) );
  OAI22_X1 U3479 ( .A1(n264), .A2(n347), .B1(\unit_memory/DRAM/n2395 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2152 ) );
  OAI22_X1 U3480 ( .A1(n264), .A2(n350), .B1(\unit_memory/DRAM/n2396 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2151 ) );
  OAI22_X1 U3481 ( .A1(n264), .A2(n353), .B1(\unit_memory/DRAM/n2397 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2150 ) );
  OAI22_X1 U3482 ( .A1(n264), .A2(n356), .B1(\unit_memory/DRAM/n2398 ), .B2(
        n255), .ZN(\unit_memory/DRAM/n2149 ) );
  OAI22_X1 U3483 ( .A1(n314), .A2(n371), .B1(\unit_memory/DRAM/n2448 ), .B2(
        n376), .ZN(\unit_memory/DRAM/n2099 ) );
  OAI22_X1 U3484 ( .A1(n317), .A2(n371), .B1(\unit_memory/DRAM/n2449 ), .B2(
        n376), .ZN(\unit_memory/DRAM/n2098 ) );
  OAI22_X1 U3485 ( .A1(n320), .A2(n371), .B1(\unit_memory/DRAM/n2450 ), .B2(
        n376), .ZN(\unit_memory/DRAM/n2097 ) );
  OAI22_X1 U3486 ( .A1(n323), .A2(n370), .B1(\unit_memory/DRAM/n2451 ), .B2(
        n377), .ZN(\unit_memory/DRAM/n2096 ) );
  OAI22_X1 U3487 ( .A1(n326), .A2(n370), .B1(\unit_memory/DRAM/n2452 ), .B2(
        n377), .ZN(\unit_memory/DRAM/n2095 ) );
  OAI22_X1 U3488 ( .A1(n329), .A2(n370), .B1(\unit_memory/DRAM/n2453 ), .B2(
        n377), .ZN(\unit_memory/DRAM/n2094 ) );
  OAI22_X1 U3489 ( .A1(n332), .A2(n370), .B1(\unit_memory/DRAM/n2454 ), .B2(
        n377), .ZN(\unit_memory/DRAM/n2093 ) );
  OAI22_X1 U3490 ( .A1(n338), .A2(n370), .B1(\unit_memory/DRAM/n2456 ), .B2(
        n378), .ZN(\unit_memory/DRAM/n2091 ) );
  OAI22_X1 U3491 ( .A1(n341), .A2(n370), .B1(\unit_memory/DRAM/n2457 ), .B2(
        n378), .ZN(\unit_memory/DRAM/n2090 ) );
  OAI22_X1 U3492 ( .A1(n344), .A2(n370), .B1(\unit_memory/DRAM/n2458 ), .B2(
        n378), .ZN(\unit_memory/DRAM/n2089 ) );
  OAI22_X1 U3493 ( .A1(n347), .A2(n370), .B1(\unit_memory/DRAM/n2459 ), .B2(
        n379), .ZN(\unit_memory/DRAM/n2088 ) );
  OAI22_X1 U3494 ( .A1(n350), .A2(n370), .B1(\unit_memory/DRAM/n2460 ), .B2(
        n379), .ZN(\unit_memory/DRAM/n2087 ) );
  OAI22_X1 U3495 ( .A1(n353), .A2(n370), .B1(\unit_memory/DRAM/n2461 ), .B2(
        n379), .ZN(\unit_memory/DRAM/n2086 ) );
  OAI22_X1 U3496 ( .A1(n356), .A2(n370), .B1(\unit_memory/DRAM/n2462 ), .B2(
        n379), .ZN(\unit_memory/DRAM/n2085 ) );
  OAI22_X1 U3497 ( .A1(n251), .A2(n381), .B1(\unit_memory/DRAM/n2463 ), .B2(
        n383), .ZN(\unit_memory/DRAM/n2084 ) );
  OAI22_X1 U3498 ( .A1(n266), .A2(n382), .B1(\unit_memory/DRAM/n2464 ), .B2(
        n383), .ZN(\unit_memory/DRAM/n2083 ) );
  OAI22_X1 U3499 ( .A1(n269), .A2(n381), .B1(\unit_memory/DRAM/n2465 ), .B2(
        n383), .ZN(\unit_memory/DRAM/n2082 ) );
  OAI22_X1 U3500 ( .A1(n272), .A2(n382), .B1(\unit_memory/DRAM/n2466 ), .B2(
        n383), .ZN(\unit_memory/DRAM/n2081 ) );
  OAI22_X1 U3501 ( .A1(n275), .A2(n381), .B1(\unit_memory/DRAM/n2467 ), .B2(
        n384), .ZN(\unit_memory/DRAM/n2080 ) );
  OAI22_X1 U3502 ( .A1(n278), .A2(n382), .B1(\unit_memory/DRAM/n2468 ), .B2(
        n384), .ZN(\unit_memory/DRAM/n2079 ) );
  OAI22_X1 U3503 ( .A1(n281), .A2(n381), .B1(\unit_memory/DRAM/n2469 ), .B2(
        n384), .ZN(\unit_memory/DRAM/n2078 ) );
  OAI22_X1 U3504 ( .A1(n284), .A2(n382), .B1(\unit_memory/DRAM/n2470 ), .B2(
        n384), .ZN(\unit_memory/DRAM/n2077 ) );
  OAI22_X1 U3505 ( .A1(n287), .A2(n382), .B1(\unit_memory/DRAM/n2471 ), .B2(
        n385), .ZN(\unit_memory/DRAM/n2076 ) );
  OAI22_X1 U3506 ( .A1(n290), .A2(n382), .B1(\unit_memory/DRAM/n2472 ), .B2(
        n385), .ZN(\unit_memory/DRAM/n2075 ) );
  OAI22_X1 U3507 ( .A1(n293), .A2(n382), .B1(\unit_memory/DRAM/n2473 ), .B2(
        n385), .ZN(\unit_memory/DRAM/n2074 ) );
  OAI22_X1 U3508 ( .A1(n296), .A2(n382), .B1(\unit_memory/DRAM/n2474 ), .B2(
        n385), .ZN(\unit_memory/DRAM/n2073 ) );
  OAI22_X1 U3509 ( .A1(n299), .A2(n382), .B1(\unit_memory/DRAM/n2475 ), .B2(
        n386), .ZN(\unit_memory/DRAM/n2072 ) );
  OAI22_X1 U3510 ( .A1(n302), .A2(n382), .B1(\unit_memory/DRAM/n2476 ), .B2(
        n386), .ZN(\unit_memory/DRAM/n2071 ) );
  OAI22_X1 U3511 ( .A1(n305), .A2(n382), .B1(\unit_memory/DRAM/n2477 ), .B2(
        n386), .ZN(\unit_memory/DRAM/n2070 ) );
  OAI22_X1 U3512 ( .A1(n308), .A2(n382), .B1(\unit_memory/DRAM/n2478 ), .B2(
        n386), .ZN(\unit_memory/DRAM/n2069 ) );
  OAI22_X1 U3513 ( .A1(n314), .A2(n382), .B1(\unit_memory/DRAM/n2480 ), .B2(
        n387), .ZN(\unit_memory/DRAM/n2067 ) );
  OAI22_X1 U3514 ( .A1(n317), .A2(n382), .B1(\unit_memory/DRAM/n2481 ), .B2(
        n387), .ZN(\unit_memory/DRAM/n2066 ) );
  OAI22_X1 U3515 ( .A1(n320), .A2(n382), .B1(\unit_memory/DRAM/n2482 ), .B2(
        n387), .ZN(\unit_memory/DRAM/n2065 ) );
  OAI22_X1 U3516 ( .A1(n323), .A2(n381), .B1(\unit_memory/DRAM/n2483 ), .B2(
        n388), .ZN(\unit_memory/DRAM/n2064 ) );
  OAI22_X1 U3517 ( .A1(n326), .A2(n381), .B1(\unit_memory/DRAM/n2484 ), .B2(
        n388), .ZN(\unit_memory/DRAM/n2063 ) );
  OAI22_X1 U3518 ( .A1(n329), .A2(n381), .B1(\unit_memory/DRAM/n2485 ), .B2(
        n388), .ZN(\unit_memory/DRAM/n2062 ) );
  OAI22_X1 U3519 ( .A1(n332), .A2(n381), .B1(\unit_memory/DRAM/n2486 ), .B2(
        n388), .ZN(\unit_memory/DRAM/n2061 ) );
  OAI22_X1 U3520 ( .A1(n338), .A2(n381), .B1(\unit_memory/DRAM/n2488 ), .B2(
        n389), .ZN(\unit_memory/DRAM/n2059 ) );
  OAI22_X1 U3521 ( .A1(n341), .A2(n381), .B1(\unit_memory/DRAM/n2489 ), .B2(
        n389), .ZN(\unit_memory/DRAM/n2058 ) );
  OAI22_X1 U3522 ( .A1(n344), .A2(n381), .B1(\unit_memory/DRAM/n2490 ), .B2(
        n389), .ZN(\unit_memory/DRAM/n2057 ) );
  OAI22_X1 U3523 ( .A1(n347), .A2(n381), .B1(\unit_memory/DRAM/n2491 ), .B2(
        n390), .ZN(\unit_memory/DRAM/n2056 ) );
  OAI22_X1 U3524 ( .A1(n350), .A2(n381), .B1(\unit_memory/DRAM/n2492 ), .B2(
        n390), .ZN(\unit_memory/DRAM/n2055 ) );
  OAI22_X1 U3525 ( .A1(n353), .A2(n381), .B1(\unit_memory/DRAM/n2493 ), .B2(
        n390), .ZN(\unit_memory/DRAM/n2054 ) );
  OAI22_X1 U3526 ( .A1(n356), .A2(n381), .B1(\unit_memory/DRAM/n2494 ), .B2(
        n390), .ZN(\unit_memory/DRAM/n2053 ) );
  OAI22_X1 U3527 ( .A1(n314), .A2(n393), .B1(\unit_memory/DRAM/n2512 ), .B2(
        n398), .ZN(\unit_memory/DRAM/n2035 ) );
  OAI22_X1 U3528 ( .A1(n317), .A2(n393), .B1(\unit_memory/DRAM/n2513 ), .B2(
        n398), .ZN(\unit_memory/DRAM/n2034 ) );
  OAI22_X1 U3529 ( .A1(n320), .A2(n393), .B1(\unit_memory/DRAM/n2514 ), .B2(
        n398), .ZN(\unit_memory/DRAM/n2033 ) );
  OAI22_X1 U3530 ( .A1(n323), .A2(n392), .B1(\unit_memory/DRAM/n2515 ), .B2(
        n399), .ZN(\unit_memory/DRAM/n2032 ) );
  OAI22_X1 U3531 ( .A1(n326), .A2(n392), .B1(\unit_memory/DRAM/n2516 ), .B2(
        n399), .ZN(\unit_memory/DRAM/n2031 ) );
  OAI22_X1 U3532 ( .A1(n329), .A2(n392), .B1(\unit_memory/DRAM/n2517 ), .B2(
        n399), .ZN(\unit_memory/DRAM/n2030 ) );
  OAI22_X1 U3533 ( .A1(n332), .A2(n392), .B1(\unit_memory/DRAM/n2518 ), .B2(
        n399), .ZN(\unit_memory/DRAM/n2029 ) );
  OAI22_X1 U3534 ( .A1(n338), .A2(n392), .B1(\unit_memory/DRAM/n2520 ), .B2(
        n400), .ZN(\unit_memory/DRAM/n2027 ) );
  OAI22_X1 U3535 ( .A1(n341), .A2(n392), .B1(\unit_memory/DRAM/n2521 ), .B2(
        n400), .ZN(\unit_memory/DRAM/n2026 ) );
  OAI22_X1 U3536 ( .A1(n344), .A2(n392), .B1(\unit_memory/DRAM/n2522 ), .B2(
        n400), .ZN(\unit_memory/DRAM/n2025 ) );
  OAI22_X1 U3537 ( .A1(n347), .A2(n392), .B1(\unit_memory/DRAM/n2523 ), .B2(
        n401), .ZN(\unit_memory/DRAM/n2024 ) );
  OAI22_X1 U3538 ( .A1(n350), .A2(n392), .B1(\unit_memory/DRAM/n2524 ), .B2(
        n401), .ZN(\unit_memory/DRAM/n2023 ) );
  OAI22_X1 U3539 ( .A1(n353), .A2(n392), .B1(\unit_memory/DRAM/n2525 ), .B2(
        n401), .ZN(\unit_memory/DRAM/n2022 ) );
  OAI22_X1 U3540 ( .A1(n356), .A2(n392), .B1(\unit_memory/DRAM/n2526 ), .B2(
        n401), .ZN(\unit_memory/DRAM/n2021 ) );
  OAI22_X1 U3541 ( .A1(n314), .A2(n415), .B1(\unit_memory/DRAM/n2576 ), .B2(
        n420), .ZN(\unit_memory/DRAM/n1971 ) );
  OAI22_X1 U3542 ( .A1(n317), .A2(n415), .B1(\unit_memory/DRAM/n2577 ), .B2(
        n420), .ZN(\unit_memory/DRAM/n1970 ) );
  OAI22_X1 U3543 ( .A1(n320), .A2(n415), .B1(\unit_memory/DRAM/n2578 ), .B2(
        n420), .ZN(\unit_memory/DRAM/n1969 ) );
  OAI22_X1 U3544 ( .A1(n323), .A2(n414), .B1(\unit_memory/DRAM/n2579 ), .B2(
        n421), .ZN(\unit_memory/DRAM/n1968 ) );
  OAI22_X1 U3545 ( .A1(n326), .A2(n414), .B1(\unit_memory/DRAM/n2580 ), .B2(
        n421), .ZN(\unit_memory/DRAM/n1967 ) );
  OAI22_X1 U3546 ( .A1(n329), .A2(n414), .B1(\unit_memory/DRAM/n2581 ), .B2(
        n421), .ZN(\unit_memory/DRAM/n1966 ) );
  OAI22_X1 U3547 ( .A1(n332), .A2(n414), .B1(\unit_memory/DRAM/n2582 ), .B2(
        n421), .ZN(\unit_memory/DRAM/n1965 ) );
  OAI22_X1 U3548 ( .A1(n338), .A2(n414), .B1(\unit_memory/DRAM/n2584 ), .B2(
        n422), .ZN(\unit_memory/DRAM/n1963 ) );
  OAI22_X1 U3549 ( .A1(n341), .A2(n414), .B1(\unit_memory/DRAM/n2585 ), .B2(
        n422), .ZN(\unit_memory/DRAM/n1962 ) );
  OAI22_X1 U3550 ( .A1(n344), .A2(n414), .B1(\unit_memory/DRAM/n2586 ), .B2(
        n422), .ZN(\unit_memory/DRAM/n1961 ) );
  OAI22_X1 U3551 ( .A1(n347), .A2(n414), .B1(\unit_memory/DRAM/n2587 ), .B2(
        n423), .ZN(\unit_memory/DRAM/n1960 ) );
  OAI22_X1 U3552 ( .A1(n350), .A2(n414), .B1(\unit_memory/DRAM/n2588 ), .B2(
        n423), .ZN(\unit_memory/DRAM/n1959 ) );
  OAI22_X1 U3553 ( .A1(n353), .A2(n414), .B1(\unit_memory/DRAM/n2589 ), .B2(
        n423), .ZN(\unit_memory/DRAM/n1958 ) );
  OAI22_X1 U3554 ( .A1(n356), .A2(n414), .B1(\unit_memory/DRAM/n2590 ), .B2(
        n423), .ZN(\unit_memory/DRAM/n1957 ) );
  OAI22_X1 U3555 ( .A1(n251), .A2(n425), .B1(\unit_memory/DRAM/n2591 ), .B2(
        n427), .ZN(\unit_memory/DRAM/n1956 ) );
  OAI22_X1 U3556 ( .A1(n266), .A2(n426), .B1(\unit_memory/DRAM/n2592 ), .B2(
        n427), .ZN(\unit_memory/DRAM/n1955 ) );
  OAI22_X1 U3557 ( .A1(n269), .A2(n425), .B1(\unit_memory/DRAM/n2593 ), .B2(
        n427), .ZN(\unit_memory/DRAM/n1954 ) );
  OAI22_X1 U3558 ( .A1(n272), .A2(n426), .B1(\unit_memory/DRAM/n2594 ), .B2(
        n427), .ZN(\unit_memory/DRAM/n1953 ) );
  OAI22_X1 U3559 ( .A1(n275), .A2(n425), .B1(\unit_memory/DRAM/n2595 ), .B2(
        n428), .ZN(\unit_memory/DRAM/n1952 ) );
  OAI22_X1 U3560 ( .A1(n278), .A2(n426), .B1(\unit_memory/DRAM/n2596 ), .B2(
        n428), .ZN(\unit_memory/DRAM/n1951 ) );
  OAI22_X1 U3561 ( .A1(n281), .A2(n425), .B1(\unit_memory/DRAM/n2597 ), .B2(
        n428), .ZN(\unit_memory/DRAM/n1950 ) );
  OAI22_X1 U3562 ( .A1(n284), .A2(n426), .B1(\unit_memory/DRAM/n2598 ), .B2(
        n428), .ZN(\unit_memory/DRAM/n1949 ) );
  OAI22_X1 U3563 ( .A1(n287), .A2(n426), .B1(\unit_memory/DRAM/n2599 ), .B2(
        n429), .ZN(\unit_memory/DRAM/n1948 ) );
  OAI22_X1 U3564 ( .A1(n290), .A2(n426), .B1(\unit_memory/DRAM/n2600 ), .B2(
        n429), .ZN(\unit_memory/DRAM/n1947 ) );
  OAI22_X1 U3565 ( .A1(n293), .A2(n426), .B1(\unit_memory/DRAM/n2601 ), .B2(
        n429), .ZN(\unit_memory/DRAM/n1946 ) );
  OAI22_X1 U3566 ( .A1(n296), .A2(n426), .B1(\unit_memory/DRAM/n2602 ), .B2(
        n429), .ZN(\unit_memory/DRAM/n1945 ) );
  OAI22_X1 U3567 ( .A1(n299), .A2(n426), .B1(\unit_memory/DRAM/n2603 ), .B2(
        n430), .ZN(\unit_memory/DRAM/n1944 ) );
  OAI22_X1 U3568 ( .A1(n302), .A2(n426), .B1(\unit_memory/DRAM/n2604 ), .B2(
        n430), .ZN(\unit_memory/DRAM/n1943 ) );
  OAI22_X1 U3569 ( .A1(n305), .A2(n426), .B1(\unit_memory/DRAM/n2605 ), .B2(
        n430), .ZN(\unit_memory/DRAM/n1942 ) );
  OAI22_X1 U3570 ( .A1(n308), .A2(n426), .B1(\unit_memory/DRAM/n2606 ), .B2(
        n430), .ZN(\unit_memory/DRAM/n1941 ) );
  OAI22_X1 U3571 ( .A1(n314), .A2(n426), .B1(\unit_memory/DRAM/n2608 ), .B2(
        n431), .ZN(\unit_memory/DRAM/n1939 ) );
  OAI22_X1 U3572 ( .A1(n317), .A2(n426), .B1(\unit_memory/DRAM/n2609 ), .B2(
        n431), .ZN(\unit_memory/DRAM/n1938 ) );
  OAI22_X1 U3573 ( .A1(n320), .A2(n426), .B1(\unit_memory/DRAM/n2610 ), .B2(
        n431), .ZN(\unit_memory/DRAM/n1937 ) );
  OAI22_X1 U3574 ( .A1(n323), .A2(n425), .B1(\unit_memory/DRAM/n2611 ), .B2(
        n432), .ZN(\unit_memory/DRAM/n1936 ) );
  OAI22_X1 U3575 ( .A1(n326), .A2(n425), .B1(\unit_memory/DRAM/n2612 ), .B2(
        n432), .ZN(\unit_memory/DRAM/n1935 ) );
  OAI22_X1 U3576 ( .A1(n329), .A2(n425), .B1(\unit_memory/DRAM/n2613 ), .B2(
        n432), .ZN(\unit_memory/DRAM/n1934 ) );
  OAI22_X1 U3577 ( .A1(n332), .A2(n425), .B1(\unit_memory/DRAM/n2614 ), .B2(
        n432), .ZN(\unit_memory/DRAM/n1933 ) );
  OAI22_X1 U3578 ( .A1(n338), .A2(n425), .B1(\unit_memory/DRAM/n2616 ), .B2(
        n433), .ZN(\unit_memory/DRAM/n1931 ) );
  OAI22_X1 U3579 ( .A1(n341), .A2(n425), .B1(\unit_memory/DRAM/n2617 ), .B2(
        n433), .ZN(\unit_memory/DRAM/n1930 ) );
  OAI22_X1 U3580 ( .A1(n344), .A2(n425), .B1(\unit_memory/DRAM/n2618 ), .B2(
        n433), .ZN(\unit_memory/DRAM/n1929 ) );
  OAI22_X1 U3581 ( .A1(n347), .A2(n425), .B1(\unit_memory/DRAM/n2619 ), .B2(
        n434), .ZN(\unit_memory/DRAM/n1928 ) );
  OAI22_X1 U3582 ( .A1(n350), .A2(n425), .B1(\unit_memory/DRAM/n2620 ), .B2(
        n434), .ZN(\unit_memory/DRAM/n1927 ) );
  OAI22_X1 U3583 ( .A1(n353), .A2(n425), .B1(\unit_memory/DRAM/n2621 ), .B2(
        n434), .ZN(\unit_memory/DRAM/n1926 ) );
  OAI22_X1 U3584 ( .A1(n356), .A2(n425), .B1(\unit_memory/DRAM/n2622 ), .B2(
        n434), .ZN(\unit_memory/DRAM/n1925 ) );
  OAI22_X1 U3585 ( .A1(n314), .A2(n448), .B1(\unit_memory/DRAM/n2672 ), .B2(
        n453), .ZN(\unit_memory/DRAM/n1875 ) );
  OAI22_X1 U3586 ( .A1(n317), .A2(n448), .B1(\unit_memory/DRAM/n2673 ), .B2(
        n453), .ZN(\unit_memory/DRAM/n1874 ) );
  OAI22_X1 U3587 ( .A1(n320), .A2(n448), .B1(\unit_memory/DRAM/n2674 ), .B2(
        n453), .ZN(\unit_memory/DRAM/n1873 ) );
  OAI22_X1 U3588 ( .A1(n323), .A2(n447), .B1(\unit_memory/DRAM/n2675 ), .B2(
        n454), .ZN(\unit_memory/DRAM/n1872 ) );
  OAI22_X1 U3589 ( .A1(n326), .A2(n447), .B1(\unit_memory/DRAM/n2676 ), .B2(
        n454), .ZN(\unit_memory/DRAM/n1871 ) );
  OAI22_X1 U3590 ( .A1(n329), .A2(n447), .B1(\unit_memory/DRAM/n2677 ), .B2(
        n454), .ZN(\unit_memory/DRAM/n1870 ) );
  OAI22_X1 U3591 ( .A1(n332), .A2(n447), .B1(\unit_memory/DRAM/n2678 ), .B2(
        n454), .ZN(\unit_memory/DRAM/n1869 ) );
  OAI22_X1 U3592 ( .A1(n338), .A2(n447), .B1(\unit_memory/DRAM/n2680 ), .B2(
        n455), .ZN(\unit_memory/DRAM/n1867 ) );
  OAI22_X1 U3593 ( .A1(n341), .A2(n447), .B1(\unit_memory/DRAM/n2681 ), .B2(
        n455), .ZN(\unit_memory/DRAM/n1866 ) );
  OAI22_X1 U3594 ( .A1(n344), .A2(n447), .B1(\unit_memory/DRAM/n2682 ), .B2(
        n455), .ZN(\unit_memory/DRAM/n1865 ) );
  OAI22_X1 U3595 ( .A1(n347), .A2(n447), .B1(\unit_memory/DRAM/n2683 ), .B2(
        n456), .ZN(\unit_memory/DRAM/n1864 ) );
  OAI22_X1 U3596 ( .A1(n350), .A2(n447), .B1(\unit_memory/DRAM/n2684 ), .B2(
        n456), .ZN(\unit_memory/DRAM/n1863 ) );
  OAI22_X1 U3597 ( .A1(n353), .A2(n447), .B1(\unit_memory/DRAM/n2685 ), .B2(
        n456), .ZN(\unit_memory/DRAM/n1862 ) );
  OAI22_X1 U3598 ( .A1(n356), .A2(n447), .B1(\unit_memory/DRAM/n2686 ), .B2(
        n456), .ZN(\unit_memory/DRAM/n1861 ) );
  OAI22_X1 U3599 ( .A1(n315), .A2(n492), .B1(\unit_memory/DRAM/n2800 ), .B2(
        n497), .ZN(\unit_memory/DRAM/n1747 ) );
  OAI22_X1 U3600 ( .A1(n318), .A2(n492), .B1(\unit_memory/DRAM/n2801 ), .B2(
        n497), .ZN(\unit_memory/DRAM/n1746 ) );
  OAI22_X1 U3601 ( .A1(n321), .A2(n492), .B1(\unit_memory/DRAM/n2802 ), .B2(
        n497), .ZN(\unit_memory/DRAM/n1745 ) );
  OAI22_X1 U3602 ( .A1(n324), .A2(n491), .B1(\unit_memory/DRAM/n2803 ), .B2(
        n498), .ZN(\unit_memory/DRAM/n1744 ) );
  OAI22_X1 U3603 ( .A1(n327), .A2(n491), .B1(\unit_memory/DRAM/n2804 ), .B2(
        n498), .ZN(\unit_memory/DRAM/n1743 ) );
  OAI22_X1 U3604 ( .A1(n330), .A2(n491), .B1(\unit_memory/DRAM/n2805 ), .B2(
        n498), .ZN(\unit_memory/DRAM/n1742 ) );
  OAI22_X1 U3605 ( .A1(n333), .A2(n491), .B1(\unit_memory/DRAM/n2806 ), .B2(
        n498), .ZN(\unit_memory/DRAM/n1741 ) );
  OAI22_X1 U3606 ( .A1(n339), .A2(n491), .B1(\unit_memory/DRAM/n2808 ), .B2(
        n499), .ZN(\unit_memory/DRAM/n1739 ) );
  OAI22_X1 U3607 ( .A1(n342), .A2(n491), .B1(\unit_memory/DRAM/n2809 ), .B2(
        n499), .ZN(\unit_memory/DRAM/n1738 ) );
  OAI22_X1 U3608 ( .A1(n345), .A2(n491), .B1(\unit_memory/DRAM/n2810 ), .B2(
        n499), .ZN(\unit_memory/DRAM/n1737 ) );
  OAI22_X1 U3609 ( .A1(n348), .A2(n491), .B1(\unit_memory/DRAM/n2811 ), .B2(
        n500), .ZN(\unit_memory/DRAM/n1736 ) );
  OAI22_X1 U3610 ( .A1(n351), .A2(n491), .B1(\unit_memory/DRAM/n2812 ), .B2(
        n500), .ZN(\unit_memory/DRAM/n1735 ) );
  OAI22_X1 U3611 ( .A1(n354), .A2(n491), .B1(\unit_memory/DRAM/n2813 ), .B2(
        n500), .ZN(\unit_memory/DRAM/n1734 ) );
  OAI22_X1 U3612 ( .A1(n357), .A2(n491), .B1(\unit_memory/DRAM/n2814 ), .B2(
        n500), .ZN(\unit_memory/DRAM/n1733 ) );
  OAI22_X1 U3613 ( .A1(n315), .A2(n437), .B1(\unit_memory/DRAM/n2640 ), .B2(
        n442), .ZN(\unit_memory/DRAM/n1907 ) );
  OAI22_X1 U3614 ( .A1(n318), .A2(n437), .B1(\unit_memory/DRAM/n2641 ), .B2(
        n442), .ZN(\unit_memory/DRAM/n1906 ) );
  OAI22_X1 U3615 ( .A1(n321), .A2(n437), .B1(\unit_memory/DRAM/n2642 ), .B2(
        n442), .ZN(\unit_memory/DRAM/n1905 ) );
  OAI22_X1 U3616 ( .A1(n324), .A2(n436), .B1(\unit_memory/DRAM/n2643 ), .B2(
        n443), .ZN(\unit_memory/DRAM/n1904 ) );
  OAI22_X1 U3617 ( .A1(n327), .A2(n436), .B1(\unit_memory/DRAM/n2644 ), .B2(
        n443), .ZN(\unit_memory/DRAM/n1903 ) );
  OAI22_X1 U3618 ( .A1(n330), .A2(n436), .B1(\unit_memory/DRAM/n2645 ), .B2(
        n443), .ZN(\unit_memory/DRAM/n1902 ) );
  OAI22_X1 U3619 ( .A1(n333), .A2(n436), .B1(\unit_memory/DRAM/n2646 ), .B2(
        n443), .ZN(\unit_memory/DRAM/n1901 ) );
  OAI22_X1 U3620 ( .A1(n339), .A2(n436), .B1(\unit_memory/DRAM/n2648 ), .B2(
        n444), .ZN(\unit_memory/DRAM/n1899 ) );
  OAI22_X1 U3621 ( .A1(n342), .A2(n436), .B1(\unit_memory/DRAM/n2649 ), .B2(
        n444), .ZN(\unit_memory/DRAM/n1898 ) );
  OAI22_X1 U3622 ( .A1(n345), .A2(n436), .B1(\unit_memory/DRAM/n2650 ), .B2(
        n444), .ZN(\unit_memory/DRAM/n1897 ) );
  OAI22_X1 U3623 ( .A1(n348), .A2(n436), .B1(\unit_memory/DRAM/n2651 ), .B2(
        n445), .ZN(\unit_memory/DRAM/n1896 ) );
  OAI22_X1 U3624 ( .A1(n351), .A2(n436), .B1(\unit_memory/DRAM/n2652 ), .B2(
        n445), .ZN(\unit_memory/DRAM/n1895 ) );
  OAI22_X1 U3625 ( .A1(n354), .A2(n436), .B1(\unit_memory/DRAM/n2653 ), .B2(
        n445), .ZN(\unit_memory/DRAM/n1894 ) );
  OAI22_X1 U3626 ( .A1(n356), .A2(n436), .B1(\unit_memory/DRAM/n2654 ), .B2(
        n445), .ZN(\unit_memory/DRAM/n1893 ) );
  OAI22_X1 U3627 ( .A1(n314), .A2(n459), .B1(\unit_memory/DRAM/n2704 ), .B2(
        n464), .ZN(\unit_memory/DRAM/n1843 ) );
  OAI22_X1 U3628 ( .A1(n317), .A2(n459), .B1(\unit_memory/DRAM/n2705 ), .B2(
        n464), .ZN(\unit_memory/DRAM/n1842 ) );
  OAI22_X1 U3629 ( .A1(n320), .A2(n459), .B1(\unit_memory/DRAM/n2706 ), .B2(
        n464), .ZN(\unit_memory/DRAM/n1841 ) );
  OAI22_X1 U3630 ( .A1(n323), .A2(n458), .B1(\unit_memory/DRAM/n2707 ), .B2(
        n465), .ZN(\unit_memory/DRAM/n1840 ) );
  OAI22_X1 U3631 ( .A1(n326), .A2(n458), .B1(\unit_memory/DRAM/n2708 ), .B2(
        n465), .ZN(\unit_memory/DRAM/n1839 ) );
  OAI22_X1 U3632 ( .A1(n329), .A2(n458), .B1(\unit_memory/DRAM/n2709 ), .B2(
        n465), .ZN(\unit_memory/DRAM/n1838 ) );
  OAI22_X1 U3633 ( .A1(n332), .A2(n458), .B1(\unit_memory/DRAM/n2710 ), .B2(
        n465), .ZN(\unit_memory/DRAM/n1837 ) );
  OAI22_X1 U3634 ( .A1(n338), .A2(n458), .B1(\unit_memory/DRAM/n2712 ), .B2(
        n466), .ZN(\unit_memory/DRAM/n1835 ) );
  OAI22_X1 U3635 ( .A1(n341), .A2(n458), .B1(\unit_memory/DRAM/n2713 ), .B2(
        n466), .ZN(\unit_memory/DRAM/n1834 ) );
  OAI22_X1 U3636 ( .A1(n344), .A2(n458), .B1(\unit_memory/DRAM/n2714 ), .B2(
        n466), .ZN(\unit_memory/DRAM/n1833 ) );
  OAI22_X1 U3637 ( .A1(n347), .A2(n458), .B1(\unit_memory/DRAM/n2715 ), .B2(
        n467), .ZN(\unit_memory/DRAM/n1832 ) );
  OAI22_X1 U3638 ( .A1(n350), .A2(n458), .B1(\unit_memory/DRAM/n2716 ), .B2(
        n467), .ZN(\unit_memory/DRAM/n1831 ) );
  OAI22_X1 U3639 ( .A1(n353), .A2(n458), .B1(\unit_memory/DRAM/n2717 ), .B2(
        n467), .ZN(\unit_memory/DRAM/n1830 ) );
  OAI22_X1 U3640 ( .A1(n356), .A2(n458), .B1(\unit_memory/DRAM/n2718 ), .B2(
        n467), .ZN(\unit_memory/DRAM/n1829 ) );
  OAI22_X1 U3641 ( .A1(n250), .A2(n469), .B1(\unit_memory/DRAM/n2719 ), .B2(
        n471), .ZN(\unit_memory/DRAM/n1828 ) );
  OAI22_X1 U3642 ( .A1(n266), .A2(n470), .B1(\unit_memory/DRAM/n2720 ), .B2(
        n471), .ZN(\unit_memory/DRAM/n1827 ) );
  OAI22_X1 U3643 ( .A1(n269), .A2(n469), .B1(\unit_memory/DRAM/n2721 ), .B2(
        n471), .ZN(\unit_memory/DRAM/n1826 ) );
  OAI22_X1 U3644 ( .A1(n272), .A2(n470), .B1(\unit_memory/DRAM/n2722 ), .B2(
        n471), .ZN(\unit_memory/DRAM/n1825 ) );
  OAI22_X1 U3645 ( .A1(n275), .A2(n469), .B1(\unit_memory/DRAM/n2723 ), .B2(
        n472), .ZN(\unit_memory/DRAM/n1824 ) );
  OAI22_X1 U3646 ( .A1(n278), .A2(n470), .B1(\unit_memory/DRAM/n2724 ), .B2(
        n472), .ZN(\unit_memory/DRAM/n1823 ) );
  OAI22_X1 U3647 ( .A1(n281), .A2(n469), .B1(\unit_memory/DRAM/n2725 ), .B2(
        n472), .ZN(\unit_memory/DRAM/n1822 ) );
  OAI22_X1 U3648 ( .A1(n284), .A2(n470), .B1(\unit_memory/DRAM/n2726 ), .B2(
        n472), .ZN(\unit_memory/DRAM/n1821 ) );
  OAI22_X1 U3649 ( .A1(n287), .A2(n470), .B1(\unit_memory/DRAM/n2727 ), .B2(
        n473), .ZN(\unit_memory/DRAM/n1820 ) );
  OAI22_X1 U3650 ( .A1(n290), .A2(n470), .B1(\unit_memory/DRAM/n2728 ), .B2(
        n473), .ZN(\unit_memory/DRAM/n1819 ) );
  OAI22_X1 U3651 ( .A1(n293), .A2(n470), .B1(\unit_memory/DRAM/n2729 ), .B2(
        n473), .ZN(\unit_memory/DRAM/n1818 ) );
  OAI22_X1 U3652 ( .A1(n296), .A2(n470), .B1(\unit_memory/DRAM/n2730 ), .B2(
        n473), .ZN(\unit_memory/DRAM/n1817 ) );
  OAI22_X1 U3653 ( .A1(n299), .A2(n470), .B1(\unit_memory/DRAM/n2731 ), .B2(
        n474), .ZN(\unit_memory/DRAM/n1816 ) );
  OAI22_X1 U3654 ( .A1(n302), .A2(n470), .B1(\unit_memory/DRAM/n2732 ), .B2(
        n474), .ZN(\unit_memory/DRAM/n1815 ) );
  OAI22_X1 U3655 ( .A1(n305), .A2(n470), .B1(\unit_memory/DRAM/n2733 ), .B2(
        n474), .ZN(\unit_memory/DRAM/n1814 ) );
  OAI22_X1 U3656 ( .A1(n308), .A2(n470), .B1(\unit_memory/DRAM/n2734 ), .B2(
        n474), .ZN(\unit_memory/DRAM/n1813 ) );
  OAI22_X1 U3657 ( .A1(n314), .A2(n470), .B1(\unit_memory/DRAM/n2736 ), .B2(
        n475), .ZN(\unit_memory/DRAM/n1811 ) );
  OAI22_X1 U3658 ( .A1(n317), .A2(n470), .B1(\unit_memory/DRAM/n2737 ), .B2(
        n475), .ZN(\unit_memory/DRAM/n1810 ) );
  OAI22_X1 U3659 ( .A1(n320), .A2(n470), .B1(\unit_memory/DRAM/n2738 ), .B2(
        n475), .ZN(\unit_memory/DRAM/n1809 ) );
  OAI22_X1 U3660 ( .A1(n323), .A2(n469), .B1(\unit_memory/DRAM/n2739 ), .B2(
        n476), .ZN(\unit_memory/DRAM/n1808 ) );
  OAI22_X1 U3661 ( .A1(n326), .A2(n469), .B1(\unit_memory/DRAM/n2740 ), .B2(
        n476), .ZN(\unit_memory/DRAM/n1807 ) );
  OAI22_X1 U3662 ( .A1(n329), .A2(n469), .B1(\unit_memory/DRAM/n2741 ), .B2(
        n476), .ZN(\unit_memory/DRAM/n1806 ) );
  OAI22_X1 U3663 ( .A1(n332), .A2(n469), .B1(\unit_memory/DRAM/n2742 ), .B2(
        n476), .ZN(\unit_memory/DRAM/n1805 ) );
  OAI22_X1 U3664 ( .A1(n338), .A2(n469), .B1(\unit_memory/DRAM/n2744 ), .B2(
        n477), .ZN(\unit_memory/DRAM/n1803 ) );
  OAI22_X1 U3665 ( .A1(n341), .A2(n469), .B1(\unit_memory/DRAM/n2745 ), .B2(
        n477), .ZN(\unit_memory/DRAM/n1802 ) );
  OAI22_X1 U3666 ( .A1(n344), .A2(n469), .B1(\unit_memory/DRAM/n2746 ), .B2(
        n477), .ZN(\unit_memory/DRAM/n1801 ) );
  OAI22_X1 U3667 ( .A1(n347), .A2(n469), .B1(\unit_memory/DRAM/n2747 ), .B2(
        n478), .ZN(\unit_memory/DRAM/n1800 ) );
  OAI22_X1 U3668 ( .A1(n350), .A2(n469), .B1(\unit_memory/DRAM/n2748 ), .B2(
        n478), .ZN(\unit_memory/DRAM/n1799 ) );
  OAI22_X1 U3669 ( .A1(n353), .A2(n469), .B1(\unit_memory/DRAM/n2749 ), .B2(
        n478), .ZN(\unit_memory/DRAM/n1798 ) );
  OAI22_X1 U3670 ( .A1(n356), .A2(n469), .B1(\unit_memory/DRAM/n2750 ), .B2(
        n478), .ZN(\unit_memory/DRAM/n1797 ) );
  OAI22_X1 U3671 ( .A1(n315), .A2(n481), .B1(\unit_memory/DRAM/n2768 ), .B2(
        n486), .ZN(\unit_memory/DRAM/n1779 ) );
  OAI22_X1 U3672 ( .A1(n318), .A2(n481), .B1(\unit_memory/DRAM/n2769 ), .B2(
        n486), .ZN(\unit_memory/DRAM/n1778 ) );
  OAI22_X1 U3673 ( .A1(n321), .A2(n481), .B1(\unit_memory/DRAM/n2770 ), .B2(
        n486), .ZN(\unit_memory/DRAM/n1777 ) );
  OAI22_X1 U3674 ( .A1(n324), .A2(n480), .B1(\unit_memory/DRAM/n2771 ), .B2(
        n487), .ZN(\unit_memory/DRAM/n1776 ) );
  OAI22_X1 U3675 ( .A1(n327), .A2(n480), .B1(\unit_memory/DRAM/n2772 ), .B2(
        n487), .ZN(\unit_memory/DRAM/n1775 ) );
  OAI22_X1 U3676 ( .A1(n330), .A2(n480), .B1(\unit_memory/DRAM/n2773 ), .B2(
        n487), .ZN(\unit_memory/DRAM/n1774 ) );
  OAI22_X1 U3677 ( .A1(n333), .A2(n480), .B1(\unit_memory/DRAM/n2774 ), .B2(
        n487), .ZN(\unit_memory/DRAM/n1773 ) );
  OAI22_X1 U3678 ( .A1(n339), .A2(n480), .B1(\unit_memory/DRAM/n2776 ), .B2(
        n488), .ZN(\unit_memory/DRAM/n1771 ) );
  OAI22_X1 U3679 ( .A1(n342), .A2(n480), .B1(\unit_memory/DRAM/n2777 ), .B2(
        n488), .ZN(\unit_memory/DRAM/n1770 ) );
  OAI22_X1 U3680 ( .A1(n345), .A2(n480), .B1(\unit_memory/DRAM/n2778 ), .B2(
        n488), .ZN(\unit_memory/DRAM/n1769 ) );
  OAI22_X1 U3681 ( .A1(n348), .A2(n480), .B1(\unit_memory/DRAM/n2779 ), .B2(
        n489), .ZN(\unit_memory/DRAM/n1768 ) );
  OAI22_X1 U3682 ( .A1(n351), .A2(n480), .B1(\unit_memory/DRAM/n2780 ), .B2(
        n489), .ZN(\unit_memory/DRAM/n1767 ) );
  OAI22_X1 U3683 ( .A1(n354), .A2(n480), .B1(\unit_memory/DRAM/n2781 ), .B2(
        n489), .ZN(\unit_memory/DRAM/n1766 ) );
  OAI22_X1 U3684 ( .A1(n356), .A2(n480), .B1(\unit_memory/DRAM/n2782 ), .B2(
        n489), .ZN(\unit_memory/DRAM/n1765 ) );
  OAI22_X1 U3685 ( .A1(n315), .A2(n503), .B1(\unit_memory/DRAM/n2832 ), .B2(
        n508), .ZN(\unit_memory/DRAM/n1715 ) );
  OAI22_X1 U3686 ( .A1(n318), .A2(n503), .B1(\unit_memory/DRAM/n2833 ), .B2(
        n508), .ZN(\unit_memory/DRAM/n1714 ) );
  OAI22_X1 U3687 ( .A1(n321), .A2(n503), .B1(\unit_memory/DRAM/n2834 ), .B2(
        n508), .ZN(\unit_memory/DRAM/n1713 ) );
  OAI22_X1 U3688 ( .A1(n324), .A2(n502), .B1(\unit_memory/DRAM/n2835 ), .B2(
        n509), .ZN(\unit_memory/DRAM/n1712 ) );
  OAI22_X1 U3689 ( .A1(n327), .A2(n502), .B1(\unit_memory/DRAM/n2836 ), .B2(
        n509), .ZN(\unit_memory/DRAM/n1711 ) );
  OAI22_X1 U3690 ( .A1(n330), .A2(n502), .B1(\unit_memory/DRAM/n2837 ), .B2(
        n509), .ZN(\unit_memory/DRAM/n1710 ) );
  OAI22_X1 U3691 ( .A1(n333), .A2(n502), .B1(\unit_memory/DRAM/n2838 ), .B2(
        n509), .ZN(\unit_memory/DRAM/n1709 ) );
  OAI22_X1 U3692 ( .A1(n339), .A2(n502), .B1(\unit_memory/DRAM/n2840 ), .B2(
        n510), .ZN(\unit_memory/DRAM/n1707 ) );
  OAI22_X1 U3693 ( .A1(n342), .A2(n502), .B1(\unit_memory/DRAM/n2841 ), .B2(
        n510), .ZN(\unit_memory/DRAM/n1706 ) );
  OAI22_X1 U3694 ( .A1(n345), .A2(n502), .B1(\unit_memory/DRAM/n2842 ), .B2(
        n510), .ZN(\unit_memory/DRAM/n1705 ) );
  OAI22_X1 U3695 ( .A1(n348), .A2(n502), .B1(\unit_memory/DRAM/n2843 ), .B2(
        n511), .ZN(\unit_memory/DRAM/n1704 ) );
  OAI22_X1 U3696 ( .A1(n351), .A2(n502), .B1(\unit_memory/DRAM/n2844 ), .B2(
        n511), .ZN(\unit_memory/DRAM/n1703 ) );
  OAI22_X1 U3697 ( .A1(n354), .A2(n502), .B1(\unit_memory/DRAM/n2845 ), .B2(
        n511), .ZN(\unit_memory/DRAM/n1702 ) );
  OAI22_X1 U3698 ( .A1(n357), .A2(n502), .B1(\unit_memory/DRAM/n2846 ), .B2(
        n511), .ZN(\unit_memory/DRAM/n1701 ) );
  OAI22_X1 U3699 ( .A1(n250), .A2(n514), .B1(\unit_memory/DRAM/n2847 ), .B2(
        n515), .ZN(\unit_memory/DRAM/n1700 ) );
  OAI22_X1 U3700 ( .A1(n267), .A2(n513), .B1(\unit_memory/DRAM/n2848 ), .B2(
        n515), .ZN(\unit_memory/DRAM/n1699 ) );
  OAI22_X1 U3701 ( .A1(n270), .A2(n514), .B1(\unit_memory/DRAM/n2849 ), .B2(
        n515), .ZN(\unit_memory/DRAM/n1698 ) );
  OAI22_X1 U3702 ( .A1(n273), .A2(n513), .B1(\unit_memory/DRAM/n2850 ), .B2(
        n515), .ZN(\unit_memory/DRAM/n1697 ) );
  OAI22_X1 U3703 ( .A1(n276), .A2(n514), .B1(\unit_memory/DRAM/n2851 ), .B2(
        n516), .ZN(\unit_memory/DRAM/n1696 ) );
  OAI22_X1 U3704 ( .A1(n279), .A2(n513), .B1(\unit_memory/DRAM/n2852 ), .B2(
        n516), .ZN(\unit_memory/DRAM/n1695 ) );
  OAI22_X1 U3705 ( .A1(n282), .A2(n514), .B1(\unit_memory/DRAM/n2853 ), .B2(
        n516), .ZN(\unit_memory/DRAM/n1694 ) );
  OAI22_X1 U3706 ( .A1(n285), .A2(n513), .B1(\unit_memory/DRAM/n2854 ), .B2(
        n516), .ZN(\unit_memory/DRAM/n1693 ) );
  OAI22_X1 U3707 ( .A1(n288), .A2(n514), .B1(\unit_memory/DRAM/n2855 ), .B2(
        n517), .ZN(\unit_memory/DRAM/n1692 ) );
  OAI22_X1 U3708 ( .A1(n291), .A2(n514), .B1(\unit_memory/DRAM/n2856 ), .B2(
        n517), .ZN(\unit_memory/DRAM/n1691 ) );
  OAI22_X1 U3709 ( .A1(n294), .A2(n514), .B1(\unit_memory/DRAM/n2857 ), .B2(
        n517), .ZN(\unit_memory/DRAM/n1690 ) );
  OAI22_X1 U3710 ( .A1(n297), .A2(n514), .B1(\unit_memory/DRAM/n2858 ), .B2(
        n517), .ZN(\unit_memory/DRAM/n1689 ) );
  OAI22_X1 U3711 ( .A1(n300), .A2(n514), .B1(\unit_memory/DRAM/n2859 ), .B2(
        n518), .ZN(\unit_memory/DRAM/n1688 ) );
  OAI22_X1 U3712 ( .A1(n303), .A2(n514), .B1(\unit_memory/DRAM/n2860 ), .B2(
        n518), .ZN(\unit_memory/DRAM/n1687 ) );
  OAI22_X1 U3713 ( .A1(n306), .A2(n514), .B1(\unit_memory/DRAM/n2861 ), .B2(
        n518), .ZN(\unit_memory/DRAM/n1686 ) );
  OAI22_X1 U3714 ( .A1(n309), .A2(n514), .B1(\unit_memory/DRAM/n2862 ), .B2(
        n518), .ZN(\unit_memory/DRAM/n1685 ) );
  OAI22_X1 U3715 ( .A1(n315), .A2(n514), .B1(\unit_memory/DRAM/n2864 ), .B2(
        n519), .ZN(\unit_memory/DRAM/n1683 ) );
  OAI22_X1 U3716 ( .A1(n318), .A2(n514), .B1(\unit_memory/DRAM/n2865 ), .B2(
        n519), .ZN(\unit_memory/DRAM/n1682 ) );
  OAI22_X1 U3717 ( .A1(n321), .A2(n514), .B1(\unit_memory/DRAM/n2866 ), .B2(
        n519), .ZN(\unit_memory/DRAM/n1681 ) );
  OAI22_X1 U3718 ( .A1(n324), .A2(n513), .B1(\unit_memory/DRAM/n2867 ), .B2(
        n520), .ZN(\unit_memory/DRAM/n1680 ) );
  OAI22_X1 U3719 ( .A1(n327), .A2(n513), .B1(\unit_memory/DRAM/n2868 ), .B2(
        n520), .ZN(\unit_memory/DRAM/n1679 ) );
  OAI22_X1 U3720 ( .A1(n330), .A2(n513), .B1(\unit_memory/DRAM/n2869 ), .B2(
        n520), .ZN(\unit_memory/DRAM/n1678 ) );
  OAI22_X1 U3721 ( .A1(n333), .A2(n513), .B1(\unit_memory/DRAM/n2870 ), .B2(
        n520), .ZN(\unit_memory/DRAM/n1677 ) );
  OAI22_X1 U3722 ( .A1(n339), .A2(n513), .B1(\unit_memory/DRAM/n2872 ), .B2(
        n521), .ZN(\unit_memory/DRAM/n1675 ) );
  OAI22_X1 U3723 ( .A1(n342), .A2(n513), .B1(\unit_memory/DRAM/n2873 ), .B2(
        n521), .ZN(\unit_memory/DRAM/n1674 ) );
  OAI22_X1 U3724 ( .A1(n345), .A2(n513), .B1(\unit_memory/DRAM/n2874 ), .B2(
        n521), .ZN(\unit_memory/DRAM/n1673 ) );
  OAI22_X1 U3725 ( .A1(n348), .A2(n513), .B1(\unit_memory/DRAM/n2875 ), .B2(
        n522), .ZN(\unit_memory/DRAM/n1672 ) );
  OAI22_X1 U3726 ( .A1(n351), .A2(n513), .B1(\unit_memory/DRAM/n2876 ), .B2(
        n522), .ZN(\unit_memory/DRAM/n1671 ) );
  OAI22_X1 U3727 ( .A1(n354), .A2(n513), .B1(\unit_memory/DRAM/n2877 ), .B2(
        n522), .ZN(\unit_memory/DRAM/n1670 ) );
  OAI22_X1 U3728 ( .A1(n357), .A2(n513), .B1(\unit_memory/DRAM/n2878 ), .B2(
        n522), .ZN(\unit_memory/DRAM/n1669 ) );
  OAI22_X1 U3729 ( .A1(n250), .A2(n437), .B1(\unit_memory/DRAM/n2623 ), .B2(
        n438), .ZN(\unit_memory/DRAM/n1924 ) );
  OAI22_X1 U3730 ( .A1(n267), .A2(n436), .B1(\unit_memory/DRAM/n2624 ), .B2(
        n438), .ZN(\unit_memory/DRAM/n1923 ) );
  OAI22_X1 U3731 ( .A1(n270), .A2(n437), .B1(\unit_memory/DRAM/n2625 ), .B2(
        n438), .ZN(\unit_memory/DRAM/n1922 ) );
  OAI22_X1 U3732 ( .A1(n273), .A2(n436), .B1(\unit_memory/DRAM/n2626 ), .B2(
        n438), .ZN(\unit_memory/DRAM/n1921 ) );
  OAI22_X1 U3733 ( .A1(n276), .A2(n437), .B1(\unit_memory/DRAM/n2627 ), .B2(
        n439), .ZN(\unit_memory/DRAM/n1920 ) );
  OAI22_X1 U3734 ( .A1(n279), .A2(n436), .B1(\unit_memory/DRAM/n2628 ), .B2(
        n439), .ZN(\unit_memory/DRAM/n1919 ) );
  OAI22_X1 U3735 ( .A1(n282), .A2(n437), .B1(\unit_memory/DRAM/n2629 ), .B2(
        n439), .ZN(\unit_memory/DRAM/n1918 ) );
  OAI22_X1 U3736 ( .A1(n285), .A2(n436), .B1(\unit_memory/DRAM/n2630 ), .B2(
        n439), .ZN(\unit_memory/DRAM/n1917 ) );
  OAI22_X1 U3737 ( .A1(n250), .A2(n447), .B1(\unit_memory/DRAM/n2655 ), .B2(
        n449), .ZN(\unit_memory/DRAM/n1892 ) );
  OAI22_X1 U3738 ( .A1(n266), .A2(n448), .B1(\unit_memory/DRAM/n2656 ), .B2(
        n449), .ZN(\unit_memory/DRAM/n1891 ) );
  OAI22_X1 U3739 ( .A1(n269), .A2(n447), .B1(\unit_memory/DRAM/n2657 ), .B2(
        n449), .ZN(\unit_memory/DRAM/n1890 ) );
  OAI22_X1 U3740 ( .A1(n272), .A2(n448), .B1(\unit_memory/DRAM/n2658 ), .B2(
        n449), .ZN(\unit_memory/DRAM/n1889 ) );
  OAI22_X1 U3741 ( .A1(n275), .A2(n447), .B1(\unit_memory/DRAM/n2659 ), .B2(
        n450), .ZN(\unit_memory/DRAM/n1888 ) );
  OAI22_X1 U3742 ( .A1(n278), .A2(n448), .B1(\unit_memory/DRAM/n2660 ), .B2(
        n450), .ZN(\unit_memory/DRAM/n1887 ) );
  OAI22_X1 U3743 ( .A1(n281), .A2(n447), .B1(\unit_memory/DRAM/n2661 ), .B2(
        n450), .ZN(\unit_memory/DRAM/n1886 ) );
  OAI22_X1 U3744 ( .A1(n284), .A2(n448), .B1(\unit_memory/DRAM/n2662 ), .B2(
        n450), .ZN(\unit_memory/DRAM/n1885 ) );
  OAI22_X1 U3745 ( .A1(n287), .A2(n448), .B1(\unit_memory/DRAM/n2663 ), .B2(
        n451), .ZN(\unit_memory/DRAM/n1884 ) );
  OAI22_X1 U3746 ( .A1(n290), .A2(n448), .B1(\unit_memory/DRAM/n2664 ), .B2(
        n451), .ZN(\unit_memory/DRAM/n1883 ) );
  OAI22_X1 U3747 ( .A1(n293), .A2(n448), .B1(\unit_memory/DRAM/n2665 ), .B2(
        n451), .ZN(\unit_memory/DRAM/n1882 ) );
  OAI22_X1 U3748 ( .A1(n296), .A2(n448), .B1(\unit_memory/DRAM/n2666 ), .B2(
        n451), .ZN(\unit_memory/DRAM/n1881 ) );
  OAI22_X1 U3749 ( .A1(n299), .A2(n448), .B1(\unit_memory/DRAM/n2667 ), .B2(
        n452), .ZN(\unit_memory/DRAM/n1880 ) );
  OAI22_X1 U3750 ( .A1(n302), .A2(n448), .B1(\unit_memory/DRAM/n2668 ), .B2(
        n452), .ZN(\unit_memory/DRAM/n1879 ) );
  OAI22_X1 U3751 ( .A1(n305), .A2(n448), .B1(\unit_memory/DRAM/n2669 ), .B2(
        n452), .ZN(\unit_memory/DRAM/n1878 ) );
  OAI22_X1 U3752 ( .A1(n308), .A2(n448), .B1(\unit_memory/DRAM/n2670 ), .B2(
        n452), .ZN(\unit_memory/DRAM/n1877 ) );
  OAI22_X1 U3753 ( .A1(n311), .A2(n448), .B1(\unit_memory/DRAM/n2671 ), .B2(
        n453), .ZN(\unit_memory/DRAM/n1876 ) );
  OAI22_X1 U3754 ( .A1(n335), .A2(n447), .B1(\unit_memory/DRAM/n2679 ), .B2(
        n455), .ZN(\unit_memory/DRAM/n1868 ) );
  OAI22_X1 U3755 ( .A1(n250), .A2(n481), .B1(\unit_memory/DRAM/n2751 ), .B2(
        n482), .ZN(\unit_memory/DRAM/n1796 ) );
  OAI22_X1 U3756 ( .A1(n267), .A2(n480), .B1(\unit_memory/DRAM/n2752 ), .B2(
        n482), .ZN(\unit_memory/DRAM/n1795 ) );
  OAI22_X1 U3757 ( .A1(n270), .A2(n481), .B1(\unit_memory/DRAM/n2753 ), .B2(
        n482), .ZN(\unit_memory/DRAM/n1794 ) );
  OAI22_X1 U3758 ( .A1(n273), .A2(n480), .B1(\unit_memory/DRAM/n2754 ), .B2(
        n482), .ZN(\unit_memory/DRAM/n1793 ) );
  OAI22_X1 U3759 ( .A1(n276), .A2(n481), .B1(\unit_memory/DRAM/n2755 ), .B2(
        n483), .ZN(\unit_memory/DRAM/n1792 ) );
  OAI22_X1 U3760 ( .A1(n279), .A2(n480), .B1(\unit_memory/DRAM/n2756 ), .B2(
        n483), .ZN(\unit_memory/DRAM/n1791 ) );
  OAI22_X1 U3761 ( .A1(n282), .A2(n481), .B1(\unit_memory/DRAM/n2757 ), .B2(
        n483), .ZN(\unit_memory/DRAM/n1790 ) );
  OAI22_X1 U3762 ( .A1(n285), .A2(n480), .B1(\unit_memory/DRAM/n2758 ), .B2(
        n483), .ZN(\unit_memory/DRAM/n1789 ) );
  OAI22_X1 U3763 ( .A1(n250), .A2(n492), .B1(\unit_memory/DRAM/n2783 ), .B2(
        n493), .ZN(\unit_memory/DRAM/n1764 ) );
  OAI22_X1 U3764 ( .A1(n267), .A2(n491), .B1(\unit_memory/DRAM/n2784 ), .B2(
        n493), .ZN(\unit_memory/DRAM/n1763 ) );
  OAI22_X1 U3765 ( .A1(n270), .A2(n492), .B1(\unit_memory/DRAM/n2785 ), .B2(
        n493), .ZN(\unit_memory/DRAM/n1762 ) );
  OAI22_X1 U3766 ( .A1(n273), .A2(n491), .B1(\unit_memory/DRAM/n2786 ), .B2(
        n493), .ZN(\unit_memory/DRAM/n1761 ) );
  OAI22_X1 U3767 ( .A1(n276), .A2(n492), .B1(\unit_memory/DRAM/n2787 ), .B2(
        n494), .ZN(\unit_memory/DRAM/n1760 ) );
  OAI22_X1 U3768 ( .A1(n279), .A2(n491), .B1(\unit_memory/DRAM/n2788 ), .B2(
        n494), .ZN(\unit_memory/DRAM/n1759 ) );
  OAI22_X1 U3769 ( .A1(n282), .A2(n492), .B1(\unit_memory/DRAM/n2789 ), .B2(
        n494), .ZN(\unit_memory/DRAM/n1758 ) );
  OAI22_X1 U3770 ( .A1(n285), .A2(n491), .B1(\unit_memory/DRAM/n2790 ), .B2(
        n494), .ZN(\unit_memory/DRAM/n1757 ) );
  OAI22_X1 U3771 ( .A1(n288), .A2(n492), .B1(\unit_memory/DRAM/n2791 ), .B2(
        n495), .ZN(\unit_memory/DRAM/n1756 ) );
  OAI22_X1 U3772 ( .A1(n291), .A2(n492), .B1(\unit_memory/DRAM/n2792 ), .B2(
        n495), .ZN(\unit_memory/DRAM/n1755 ) );
  OAI22_X1 U3773 ( .A1(n294), .A2(n492), .B1(\unit_memory/DRAM/n2793 ), .B2(
        n495), .ZN(\unit_memory/DRAM/n1754 ) );
  OAI22_X1 U3774 ( .A1(n297), .A2(n492), .B1(\unit_memory/DRAM/n2794 ), .B2(
        n495), .ZN(\unit_memory/DRAM/n1753 ) );
  OAI22_X1 U3775 ( .A1(n300), .A2(n492), .B1(\unit_memory/DRAM/n2795 ), .B2(
        n496), .ZN(\unit_memory/DRAM/n1752 ) );
  OAI22_X1 U3776 ( .A1(n303), .A2(n492), .B1(\unit_memory/DRAM/n2796 ), .B2(
        n496), .ZN(\unit_memory/DRAM/n1751 ) );
  OAI22_X1 U3777 ( .A1(n306), .A2(n492), .B1(\unit_memory/DRAM/n2797 ), .B2(
        n496), .ZN(\unit_memory/DRAM/n1750 ) );
  OAI22_X1 U3778 ( .A1(n309), .A2(n492), .B1(\unit_memory/DRAM/n2798 ), .B2(
        n496), .ZN(\unit_memory/DRAM/n1749 ) );
  OAI22_X1 U3779 ( .A1(n312), .A2(n492), .B1(\unit_memory/DRAM/n2799 ), .B2(
        n497), .ZN(\unit_memory/DRAM/n1748 ) );
  OAI22_X1 U3780 ( .A1(n336), .A2(n491), .B1(\unit_memory/DRAM/n2807 ), .B2(
        n499), .ZN(\unit_memory/DRAM/n1740 ) );
  OAI22_X1 U3781 ( .A1(n288), .A2(n437), .B1(\unit_memory/DRAM/n2631 ), .B2(
        n440), .ZN(\unit_memory/DRAM/n1916 ) );
  OAI22_X1 U3782 ( .A1(n291), .A2(n437), .B1(\unit_memory/DRAM/n2632 ), .B2(
        n440), .ZN(\unit_memory/DRAM/n1915 ) );
  OAI22_X1 U3783 ( .A1(n294), .A2(n437), .B1(\unit_memory/DRAM/n2633 ), .B2(
        n440), .ZN(\unit_memory/DRAM/n1914 ) );
  OAI22_X1 U3784 ( .A1(n297), .A2(n437), .B1(\unit_memory/DRAM/n2634 ), .B2(
        n440), .ZN(\unit_memory/DRAM/n1913 ) );
  OAI22_X1 U3785 ( .A1(n300), .A2(n437), .B1(\unit_memory/DRAM/n2635 ), .B2(
        n441), .ZN(\unit_memory/DRAM/n1912 ) );
  OAI22_X1 U3786 ( .A1(n303), .A2(n437), .B1(\unit_memory/DRAM/n2636 ), .B2(
        n441), .ZN(\unit_memory/DRAM/n1911 ) );
  OAI22_X1 U3787 ( .A1(n306), .A2(n437), .B1(\unit_memory/DRAM/n2637 ), .B2(
        n441), .ZN(\unit_memory/DRAM/n1910 ) );
  OAI22_X1 U3788 ( .A1(n309), .A2(n437), .B1(\unit_memory/DRAM/n2638 ), .B2(
        n441), .ZN(\unit_memory/DRAM/n1909 ) );
  OAI22_X1 U3789 ( .A1(n312), .A2(n437), .B1(\unit_memory/DRAM/n2639 ), .B2(
        n442), .ZN(\unit_memory/DRAM/n1908 ) );
  OAI22_X1 U3790 ( .A1(n336), .A2(n436), .B1(\unit_memory/DRAM/n2647 ), .B2(
        n444), .ZN(\unit_memory/DRAM/n1900 ) );
  OAI22_X1 U3791 ( .A1(n250), .A2(n458), .B1(\unit_memory/DRAM/n2687 ), .B2(
        n460), .ZN(\unit_memory/DRAM/n1860 ) );
  OAI22_X1 U3792 ( .A1(n266), .A2(n459), .B1(\unit_memory/DRAM/n2688 ), .B2(
        n460), .ZN(\unit_memory/DRAM/n1859 ) );
  OAI22_X1 U3793 ( .A1(n269), .A2(n458), .B1(\unit_memory/DRAM/n2689 ), .B2(
        n460), .ZN(\unit_memory/DRAM/n1858 ) );
  OAI22_X1 U3794 ( .A1(n272), .A2(n459), .B1(\unit_memory/DRAM/n2690 ), .B2(
        n460), .ZN(\unit_memory/DRAM/n1857 ) );
  OAI22_X1 U3795 ( .A1(n275), .A2(n458), .B1(\unit_memory/DRAM/n2691 ), .B2(
        n461), .ZN(\unit_memory/DRAM/n1856 ) );
  OAI22_X1 U3796 ( .A1(n278), .A2(n459), .B1(\unit_memory/DRAM/n2692 ), .B2(
        n461), .ZN(\unit_memory/DRAM/n1855 ) );
  OAI22_X1 U3797 ( .A1(n281), .A2(n458), .B1(\unit_memory/DRAM/n2693 ), .B2(
        n461), .ZN(\unit_memory/DRAM/n1854 ) );
  OAI22_X1 U3798 ( .A1(n284), .A2(n459), .B1(\unit_memory/DRAM/n2694 ), .B2(
        n461), .ZN(\unit_memory/DRAM/n1853 ) );
  OAI22_X1 U3799 ( .A1(n287), .A2(n459), .B1(\unit_memory/DRAM/n2695 ), .B2(
        n462), .ZN(\unit_memory/DRAM/n1852 ) );
  OAI22_X1 U3800 ( .A1(n290), .A2(n459), .B1(\unit_memory/DRAM/n2696 ), .B2(
        n462), .ZN(\unit_memory/DRAM/n1851 ) );
  OAI22_X1 U3801 ( .A1(n293), .A2(n459), .B1(\unit_memory/DRAM/n2697 ), .B2(
        n462), .ZN(\unit_memory/DRAM/n1850 ) );
  OAI22_X1 U3802 ( .A1(n296), .A2(n459), .B1(\unit_memory/DRAM/n2698 ), .B2(
        n462), .ZN(\unit_memory/DRAM/n1849 ) );
  OAI22_X1 U3803 ( .A1(n299), .A2(n459), .B1(\unit_memory/DRAM/n2699 ), .B2(
        n463), .ZN(\unit_memory/DRAM/n1848 ) );
  OAI22_X1 U3804 ( .A1(n302), .A2(n459), .B1(\unit_memory/DRAM/n2700 ), .B2(
        n463), .ZN(\unit_memory/DRAM/n1847 ) );
  OAI22_X1 U3805 ( .A1(n305), .A2(n459), .B1(\unit_memory/DRAM/n2701 ), .B2(
        n463), .ZN(\unit_memory/DRAM/n1846 ) );
  OAI22_X1 U3806 ( .A1(n308), .A2(n459), .B1(\unit_memory/DRAM/n2702 ), .B2(
        n463), .ZN(\unit_memory/DRAM/n1845 ) );
  OAI22_X1 U3807 ( .A1(n311), .A2(n459), .B1(\unit_memory/DRAM/n2703 ), .B2(
        n464), .ZN(\unit_memory/DRAM/n1844 ) );
  OAI22_X1 U3808 ( .A1(n335), .A2(n458), .B1(\unit_memory/DRAM/n2711 ), .B2(
        n466), .ZN(\unit_memory/DRAM/n1836 ) );
  OAI22_X1 U3809 ( .A1(n311), .A2(n470), .B1(\unit_memory/DRAM/n2735 ), .B2(
        n475), .ZN(\unit_memory/DRAM/n1812 ) );
  OAI22_X1 U3810 ( .A1(n335), .A2(n469), .B1(\unit_memory/DRAM/n2743 ), .B2(
        n477), .ZN(\unit_memory/DRAM/n1804 ) );
  OAI22_X1 U3811 ( .A1(n288), .A2(n481), .B1(\unit_memory/DRAM/n2759 ), .B2(
        n484), .ZN(\unit_memory/DRAM/n1788 ) );
  OAI22_X1 U3812 ( .A1(n291), .A2(n481), .B1(\unit_memory/DRAM/n2760 ), .B2(
        n484), .ZN(\unit_memory/DRAM/n1787 ) );
  OAI22_X1 U3813 ( .A1(n294), .A2(n481), .B1(\unit_memory/DRAM/n2761 ), .B2(
        n484), .ZN(\unit_memory/DRAM/n1786 ) );
  OAI22_X1 U3814 ( .A1(n297), .A2(n481), .B1(\unit_memory/DRAM/n2762 ), .B2(
        n484), .ZN(\unit_memory/DRAM/n1785 ) );
  OAI22_X1 U3815 ( .A1(n300), .A2(n481), .B1(\unit_memory/DRAM/n2763 ), .B2(
        n485), .ZN(\unit_memory/DRAM/n1784 ) );
  OAI22_X1 U3816 ( .A1(n303), .A2(n481), .B1(\unit_memory/DRAM/n2764 ), .B2(
        n485), .ZN(\unit_memory/DRAM/n1783 ) );
  OAI22_X1 U3817 ( .A1(n306), .A2(n481), .B1(\unit_memory/DRAM/n2765 ), .B2(
        n485), .ZN(\unit_memory/DRAM/n1782 ) );
  OAI22_X1 U3818 ( .A1(n309), .A2(n481), .B1(\unit_memory/DRAM/n2766 ), .B2(
        n485), .ZN(\unit_memory/DRAM/n1781 ) );
  OAI22_X1 U3819 ( .A1(n312), .A2(n481), .B1(\unit_memory/DRAM/n2767 ), .B2(
        n486), .ZN(\unit_memory/DRAM/n1780 ) );
  OAI22_X1 U3820 ( .A1(n336), .A2(n480), .B1(\unit_memory/DRAM/n2775 ), .B2(
        n488), .ZN(\unit_memory/DRAM/n1772 ) );
  OAI22_X1 U3821 ( .A1(n250), .A2(n503), .B1(\unit_memory/DRAM/n2815 ), .B2(
        n504), .ZN(\unit_memory/DRAM/n1732 ) );
  OAI22_X1 U3822 ( .A1(n267), .A2(n502), .B1(\unit_memory/DRAM/n2816 ), .B2(
        n504), .ZN(\unit_memory/DRAM/n1731 ) );
  OAI22_X1 U3823 ( .A1(n270), .A2(n503), .B1(\unit_memory/DRAM/n2817 ), .B2(
        n504), .ZN(\unit_memory/DRAM/n1730 ) );
  OAI22_X1 U3824 ( .A1(n273), .A2(n502), .B1(\unit_memory/DRAM/n2818 ), .B2(
        n504), .ZN(\unit_memory/DRAM/n1729 ) );
  OAI22_X1 U3825 ( .A1(n276), .A2(n503), .B1(\unit_memory/DRAM/n2819 ), .B2(
        n505), .ZN(\unit_memory/DRAM/n1728 ) );
  OAI22_X1 U3826 ( .A1(n279), .A2(n502), .B1(\unit_memory/DRAM/n2820 ), .B2(
        n505), .ZN(\unit_memory/DRAM/n1727 ) );
  OAI22_X1 U3827 ( .A1(n282), .A2(n503), .B1(\unit_memory/DRAM/n2821 ), .B2(
        n505), .ZN(\unit_memory/DRAM/n1726 ) );
  OAI22_X1 U3828 ( .A1(n285), .A2(n502), .B1(\unit_memory/DRAM/n2822 ), .B2(
        n505), .ZN(\unit_memory/DRAM/n1725 ) );
  OAI22_X1 U3829 ( .A1(n288), .A2(n503), .B1(\unit_memory/DRAM/n2823 ), .B2(
        n506), .ZN(\unit_memory/DRAM/n1724 ) );
  OAI22_X1 U3830 ( .A1(n291), .A2(n503), .B1(\unit_memory/DRAM/n2824 ), .B2(
        n506), .ZN(\unit_memory/DRAM/n1723 ) );
  OAI22_X1 U3831 ( .A1(n294), .A2(n503), .B1(\unit_memory/DRAM/n2825 ), .B2(
        n506), .ZN(\unit_memory/DRAM/n1722 ) );
  OAI22_X1 U3832 ( .A1(n297), .A2(n503), .B1(\unit_memory/DRAM/n2826 ), .B2(
        n506), .ZN(\unit_memory/DRAM/n1721 ) );
  OAI22_X1 U3833 ( .A1(n300), .A2(n503), .B1(\unit_memory/DRAM/n2827 ), .B2(
        n507), .ZN(\unit_memory/DRAM/n1720 ) );
  OAI22_X1 U3834 ( .A1(n303), .A2(n503), .B1(\unit_memory/DRAM/n2828 ), .B2(
        n507), .ZN(\unit_memory/DRAM/n1719 ) );
  OAI22_X1 U3835 ( .A1(n306), .A2(n503), .B1(\unit_memory/DRAM/n2829 ), .B2(
        n507), .ZN(\unit_memory/DRAM/n1718 ) );
  OAI22_X1 U3836 ( .A1(n309), .A2(n503), .B1(\unit_memory/DRAM/n2830 ), .B2(
        n507), .ZN(\unit_memory/DRAM/n1717 ) );
  OAI22_X1 U3837 ( .A1(n312), .A2(n503), .B1(\unit_memory/DRAM/n2831 ), .B2(
        n508), .ZN(\unit_memory/DRAM/n1716 ) );
  OAI22_X1 U3838 ( .A1(n336), .A2(n502), .B1(\unit_memory/DRAM/n2839 ), .B2(
        n510), .ZN(\unit_memory/DRAM/n1708 ) );
  OAI22_X1 U3839 ( .A1(n312), .A2(n514), .B1(\unit_memory/DRAM/n2863 ), .B2(
        n519), .ZN(\unit_memory/DRAM/n1684 ) );
  OAI22_X1 U3840 ( .A1(n336), .A2(n513), .B1(\unit_memory/DRAM/n2871 ), .B2(
        n521), .ZN(\unit_memory/DRAM/n1676 ) );
  OAI22_X1 U3841 ( .A1(n1285), .A2(\unit_decode/n2117 ), .B1(
        \unit_decode/n3626 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_31/n5 )
         );
  OAI22_X1 U3842 ( .A1(n1285), .A2(n116), .B1(n1396), .B2(n1296), .ZN(
        \unit_decode/RD1reg/ffi_1/n5 ) );
  OAI22_X1 U3843 ( .A1(n1285), .A2(\unit_decode/n2192 ), .B1(n1375), .B2(n1296), .ZN(\unit_decode/RD1reg/ffi_2/n5 ) );
  OAI22_X1 U3844 ( .A1(n1285), .A2(\unit_decode/n2191 ), .B1(n1386), .B2(n1296), .ZN(\unit_decode/RD1reg/ffi_3/n5 ) );
  OAI22_X1 U3845 ( .A1(n1289), .A2(\unit_decode/n2190 ), .B1(n1397), .B2(n1296), .ZN(\unit_decode/RD1reg/ffi_4/n5 ) );
  OAI22_X1 U3846 ( .A1(n1290), .A2(\unit_decode/n1109 ), .B1(n1302), .B2(
        \unit_decode/n239 ), .ZN(\unit_decode/Breg/ffi_0/n5 ) );
  INV_X1 U3847 ( .A(\unit_decode/registerB[0] ), .ZN(\unit_decode/n1109 ) );
  OAI22_X1 U3848 ( .A1(n1290), .A2(\unit_decode/n1110 ), .B1(n1302), .B2(
        \unit_decode/n233 ), .ZN(\unit_decode/Breg/ffi_1/n5 ) );
  INV_X1 U3849 ( .A(\unit_decode/registerB[1] ), .ZN(\unit_decode/n1110 ) );
  OAI22_X1 U3850 ( .A1(n1289), .A2(\unit_decode/n1111 ), .B1(n1301), .B2(
        \unit_decode/n227 ), .ZN(\unit_decode/Breg/ffi_2/n5 ) );
  INV_X1 U3851 ( .A(\unit_decode/registerB[2] ), .ZN(\unit_decode/n1111 ) );
  OAI22_X1 U3852 ( .A1(n1288), .A2(\unit_decode/n1112 ), .B1(n1301), .B2(
        \unit_decode/n235 ), .ZN(\unit_decode/Breg/ffi_3/n5 ) );
  INV_X1 U3853 ( .A(\unit_decode/registerB[3] ), .ZN(\unit_decode/n1112 ) );
  OAI22_X1 U3854 ( .A1(n1288), .A2(\unit_decode/n1113 ), .B1(n1300), .B2(
        \unit_decode/n221 ), .ZN(\unit_decode/Breg/ffi_4/n5 ) );
  INV_X1 U3855 ( .A(\unit_decode/registerB[4] ), .ZN(\unit_decode/n1113 ) );
  OAI22_X1 U3856 ( .A1(n1288), .A2(\unit_decode/n1114 ), .B1(n1300), .B2(
        \unit_decode/n223 ), .ZN(\unit_decode/Breg/ffi_5/n5 ) );
  INV_X1 U3857 ( .A(\unit_decode/registerB[5] ), .ZN(\unit_decode/n1114 ) );
  OAI22_X1 U3858 ( .A1(n1288), .A2(\unit_decode/n1115 ), .B1(n1300), .B2(
        \unit_decode/n207 ), .ZN(\unit_decode/Breg/ffi_6/n5 ) );
  INV_X1 U3859 ( .A(\unit_decode/registerB[6] ), .ZN(\unit_decode/n1115 ) );
  OAI22_X1 U3860 ( .A1(n1288), .A2(\unit_decode/n1116 ), .B1(n1300), .B2(
        \unit_decode/n219 ), .ZN(\unit_decode/Breg/ffi_7/n5 ) );
  INV_X1 U3861 ( .A(\unit_decode/registerB[7] ), .ZN(\unit_decode/n1116 ) );
  OAI22_X1 U3862 ( .A1(n1288), .A2(\unit_decode/n1117 ), .B1(n1300), .B2(
        \unit_decode/n3624 ), .ZN(\unit_decode/Breg/ffi_8/n5 ) );
  INV_X1 U3863 ( .A(\unit_decode/registerB[8] ), .ZN(\unit_decode/n1117 ) );
  OAI22_X1 U3864 ( .A1(n1288), .A2(\unit_decode/n1118 ), .B1(n1300), .B2(
        \unit_decode/n3623 ), .ZN(\unit_decode/Breg/ffi_9/n5 ) );
  INV_X1 U3865 ( .A(\unit_decode/registerB[9] ), .ZN(\unit_decode/n1118 ) );
  OAI22_X1 U3866 ( .A1(n1290), .A2(\unit_decode/n1119 ), .B1(n1302), .B2(
        \unit_decode/n3622 ), .ZN(\unit_decode/Breg/ffi_10/n5 ) );
  INV_X1 U3867 ( .A(\unit_decode/registerB[10] ), .ZN(\unit_decode/n1119 ) );
  OAI22_X1 U3868 ( .A1(n1290), .A2(\unit_decode/n1120 ), .B1(n1302), .B2(
        \unit_decode/n3558 ), .ZN(\unit_decode/Breg/ffi_11/n5 ) );
  INV_X1 U3869 ( .A(\unit_decode/registerB[11] ), .ZN(\unit_decode/n1120 ) );
  OAI22_X1 U3870 ( .A1(n1290), .A2(\unit_decode/n1121 ), .B1(n1302), .B2(
        \unit_decode/n3557 ), .ZN(\unit_decode/Breg/ffi_12/n5 ) );
  INV_X1 U3871 ( .A(\unit_decode/registerB[12] ), .ZN(\unit_decode/n1121 ) );
  OAI22_X1 U3872 ( .A1(n1290), .A2(\unit_decode/n1122 ), .B1(n1302), .B2(
        \unit_decode/n3556 ), .ZN(\unit_decode/Breg/ffi_13/n5 ) );
  INV_X1 U3873 ( .A(\unit_decode/registerB[13] ), .ZN(\unit_decode/n1122 ) );
  OAI22_X1 U3874 ( .A1(n1290), .A2(\unit_decode/n1123 ), .B1(n1302), .B2(
        \unit_decode/n3555 ), .ZN(\unit_decode/Breg/ffi_14/n5 ) );
  INV_X1 U3875 ( .A(\unit_decode/registerB[14] ), .ZN(\unit_decode/n1123 ) );
  OAI22_X1 U3876 ( .A1(n1290), .A2(\unit_decode/n1124 ), .B1(n1302), .B2(
        \unit_decode/n3554 ), .ZN(\unit_decode/Breg/ffi_15/n5 ) );
  INV_X1 U3877 ( .A(\unit_decode/registerB[15] ), .ZN(\unit_decode/n1124 ) );
  OAI22_X1 U3878 ( .A1(n1290), .A2(\unit_decode/n1125 ), .B1(n1302), .B2(
        \unit_decode/n3553 ), .ZN(\unit_decode/Breg/ffi_16/n5 ) );
  INV_X1 U3879 ( .A(\unit_decode/registerB[16] ), .ZN(\unit_decode/n1125 ) );
  OAI22_X1 U3880 ( .A1(n1290), .A2(\unit_decode/n1126 ), .B1(n1302), .B2(
        \unit_decode/n3552 ), .ZN(\unit_decode/Breg/ffi_17/n5 ) );
  INV_X1 U3881 ( .A(\unit_decode/registerB[17] ), .ZN(\unit_decode/n1126 ) );
  OAI22_X1 U3882 ( .A1(n1289), .A2(\unit_decode/n1127 ), .B1(n1302), .B2(
        \unit_decode/n3551 ), .ZN(\unit_decode/Breg/ffi_18/n5 ) );
  INV_X1 U3883 ( .A(\unit_decode/registerB[18] ), .ZN(\unit_decode/n1127 ) );
  OAI22_X1 U3884 ( .A1(n1289), .A2(\unit_decode/n1128 ), .B1(n1302), .B2(
        \unit_decode/n3550 ), .ZN(\unit_decode/Breg/ffi_19/n5 ) );
  INV_X1 U3885 ( .A(\unit_decode/registerB[19] ), .ZN(\unit_decode/n1128 ) );
  OAI22_X1 U3886 ( .A1(n1289), .A2(\unit_decode/n1129 ), .B1(n1301), .B2(
        \unit_decode/n3549 ), .ZN(\unit_decode/Breg/ffi_20/n5 ) );
  INV_X1 U3887 ( .A(\unit_decode/registerB[20] ), .ZN(\unit_decode/n1129 ) );
  OAI22_X1 U3888 ( .A1(n1289), .A2(\unit_decode/n1130 ), .B1(n1301), .B2(
        \unit_decode/n3548 ), .ZN(\unit_decode/Breg/ffi_21/n5 ) );
  INV_X1 U3889 ( .A(\unit_decode/registerB[21] ), .ZN(\unit_decode/n1130 ) );
  OAI22_X1 U3890 ( .A1(n1289), .A2(\unit_decode/n1131 ), .B1(n1301), .B2(
        \unit_decode/n3547 ), .ZN(\unit_decode/Breg/ffi_22/n5 ) );
  INV_X1 U3891 ( .A(\unit_decode/registerB[22] ), .ZN(\unit_decode/n1131 ) );
  OAI22_X1 U3892 ( .A1(n1289), .A2(\unit_decode/n1132 ), .B1(n1301), .B2(
        \unit_decode/n3546 ), .ZN(\unit_decode/Breg/ffi_23/n5 ) );
  INV_X1 U3893 ( .A(\unit_decode/registerB[23] ), .ZN(\unit_decode/n1132 ) );
  OAI22_X1 U3894 ( .A1(n1289), .A2(\unit_decode/n1133 ), .B1(n1301), .B2(
        \unit_decode/n3545 ), .ZN(\unit_decode/Breg/ffi_24/n5 ) );
  INV_X1 U3895 ( .A(\unit_decode/registerB[24] ), .ZN(\unit_decode/n1133 ) );
  OAI22_X1 U3896 ( .A1(n1289), .A2(\unit_decode/n1134 ), .B1(n1301), .B2(
        \unit_decode/n3544 ), .ZN(\unit_decode/Breg/ffi_25/n5 ) );
  INV_X1 U3897 ( .A(\unit_decode/registerB[25] ), .ZN(\unit_decode/n1134 ) );
  OAI22_X1 U3898 ( .A1(n1289), .A2(\unit_decode/n1135 ), .B1(n1301), .B2(
        \unit_decode/n3543 ), .ZN(\unit_decode/Breg/ffi_26/n5 ) );
  INV_X1 U3899 ( .A(\unit_decode/registerB[26] ), .ZN(\unit_decode/n1135 ) );
  OAI22_X1 U3900 ( .A1(n1289), .A2(\unit_decode/n1136 ), .B1(n1301), .B2(
        \unit_decode/n3542 ), .ZN(\unit_decode/Breg/ffi_27/n5 ) );
  INV_X1 U3901 ( .A(\unit_decode/registerB[27] ), .ZN(\unit_decode/n1136 ) );
  OAI22_X1 U3902 ( .A1(n1288), .A2(\unit_decode/n1137 ), .B1(n1301), .B2(
        \unit_decode/n3541 ), .ZN(\unit_decode/Breg/ffi_28/n5 ) );
  INV_X1 U3903 ( .A(\unit_decode/registerB[28] ), .ZN(\unit_decode/n1137 ) );
  OAI22_X1 U3904 ( .A1(n1288), .A2(\unit_decode/n1138 ), .B1(n1301), .B2(
        \unit_decode/n3540 ), .ZN(\unit_decode/Breg/ffi_29/n5 ) );
  INV_X1 U3905 ( .A(\unit_decode/registerB[29] ), .ZN(\unit_decode/n1138 ) );
  OAI22_X1 U3906 ( .A1(n1288), .A2(\unit_decode/n1139 ), .B1(n1301), .B2(
        \unit_decode/n3539 ), .ZN(\unit_decode/Breg/ffi_30/n5 ) );
  INV_X1 U3907 ( .A(\unit_decode/registerB[30] ), .ZN(\unit_decode/n1139 ) );
  OAI22_X1 U3908 ( .A1(n1288), .A2(\unit_decode/n1140 ), .B1(n1300), .B2(
        \unit_decode/n3538 ), .ZN(\unit_decode/Breg/ffi_31/n5 ) );
  INV_X1 U3909 ( .A(\unit_decode/registerB[31] ), .ZN(\unit_decode/n1140 ) );
  OAI22_X1 U3910 ( .A1(n1292), .A2(\unit_decode/n1143 ), .B1(n1304), .B2(
        \unit_decode/n193 ), .ZN(\unit_decode/Areg/ffi_2/n5 ) );
  INV_X1 U3911 ( .A(\unit_decode/registerA[2] ), .ZN(\unit_decode/n1143 ) );
  OAI22_X1 U3912 ( .A1(n1291), .A2(\unit_decode/n1144 ), .B1(n1303), .B2(
        \unit_decode/n215 ), .ZN(\unit_decode/Areg/ffi_3/n5 ) );
  INV_X1 U3913 ( .A(\unit_decode/registerA[3] ), .ZN(\unit_decode/n1144 ) );
  OAI22_X1 U3914 ( .A1(n1291), .A2(\unit_decode/n1145 ), .B1(n1303), .B2(
        \unit_decode/n3537 ), .ZN(\unit_decode/Areg/ffi_4/n5 ) );
  INV_X1 U3915 ( .A(\unit_decode/registerA[4] ), .ZN(\unit_decode/n1145 ) );
  OAI22_X1 U3916 ( .A1(n1291), .A2(\unit_decode/n1146 ), .B1(n1303), .B2(
        \unit_decode/n3536 ), .ZN(\unit_decode/Areg/ffi_5/n5 ) );
  INV_X1 U3917 ( .A(\unit_decode/registerA[5] ), .ZN(\unit_decode/n1146 ) );
  OAI22_X1 U3918 ( .A1(n1291), .A2(\unit_decode/n1147 ), .B1(n1303), .B2(
        \unit_decode/n3535 ), .ZN(\unit_decode/Areg/ffi_6/n5 ) );
  INV_X1 U3919 ( .A(\unit_decode/registerA[6] ), .ZN(\unit_decode/n1147 ) );
  OAI22_X1 U3920 ( .A1(n1291), .A2(\unit_decode/n1148 ), .B1(n1303), .B2(
        \unit_decode/n3534 ), .ZN(\unit_decode/Areg/ffi_7/n5 ) );
  INV_X1 U3921 ( .A(\unit_decode/registerA[7] ), .ZN(\unit_decode/n1148 ) );
  OAI22_X1 U3922 ( .A1(n1290), .A2(\unit_decode/n1149 ), .B1(n1303), .B2(
        \unit_decode/n3533 ), .ZN(\unit_decode/Areg/ffi_8/n5 ) );
  INV_X1 U3923 ( .A(\unit_decode/registerA[8] ), .ZN(\unit_decode/n1149 ) );
  OAI22_X1 U3924 ( .A1(n1290), .A2(\unit_decode/n1150 ), .B1(n1302), .B2(
        \unit_decode/n3532 ), .ZN(\unit_decode/Areg/ffi_9/n5 ) );
  INV_X1 U3925 ( .A(\unit_decode/registerA[9] ), .ZN(\unit_decode/n1150 ) );
  OAI22_X1 U3926 ( .A1(n1287), .A2(\unit_decode/n1154 ), .B1(n1304), .B2(
        \unit_decode/n3528 ), .ZN(\unit_decode/Areg/ffi_13/n5 ) );
  INV_X1 U3927 ( .A(\unit_decode/registerA[13] ), .ZN(\unit_decode/n1154 ) );
  OAI22_X1 U3928 ( .A1(n1292), .A2(\unit_decode/n1155 ), .B1(n1304), .B2(
        \unit_decode/n3527 ), .ZN(\unit_decode/Areg/ffi_14/n5 ) );
  INV_X1 U3929 ( .A(\unit_decode/registerA[14] ), .ZN(\unit_decode/n1155 ) );
  OAI22_X1 U3930 ( .A1(n1292), .A2(\unit_decode/n1156 ), .B1(n1304), .B2(
        \unit_decode/n3526 ), .ZN(\unit_decode/Areg/ffi_15/n5 ) );
  INV_X1 U3931 ( .A(\unit_decode/registerA[15] ), .ZN(\unit_decode/n1156 ) );
  OAI22_X1 U3932 ( .A1(n1292), .A2(\unit_decode/n1157 ), .B1(n1304), .B2(
        \unit_decode/n3525 ), .ZN(\unit_decode/Areg/ffi_16/n5 ) );
  INV_X1 U3933 ( .A(\unit_decode/registerA[16] ), .ZN(\unit_decode/n1157 ) );
  OAI22_X1 U3934 ( .A1(n1292), .A2(\unit_decode/n1158 ), .B1(n1304), .B2(
        \unit_decode/n3524 ), .ZN(\unit_decode/Areg/ffi_17/n5 ) );
  INV_X1 U3935 ( .A(\unit_decode/registerA[17] ), .ZN(\unit_decode/n1158 ) );
  OAI22_X1 U3936 ( .A1(n1292), .A2(\unit_decode/n1159 ), .B1(n1304), .B2(
        \unit_decode/n3523 ), .ZN(\unit_decode/Areg/ffi_18/n5 ) );
  INV_X1 U3937 ( .A(\unit_decode/registerA[18] ), .ZN(\unit_decode/n1159 ) );
  OAI22_X1 U3938 ( .A1(n1292), .A2(\unit_decode/n1160 ), .B1(n1304), .B2(
        \unit_decode/n3599 ), .ZN(\unit_decode/Areg/ffi_19/n5 ) );
  INV_X1 U3939 ( .A(\unit_decode/registerA[19] ), .ZN(\unit_decode/n1160 ) );
  OAI22_X1 U3940 ( .A1(n1292), .A2(\unit_decode/n1161 ), .B1(n1304), .B2(
        \unit_decode/n3598 ), .ZN(\unit_decode/Areg/ffi_20/n5 ) );
  INV_X1 U3941 ( .A(\unit_decode/registerA[20] ), .ZN(\unit_decode/n1161 ) );
  OAI22_X1 U3942 ( .A1(n1292), .A2(\unit_decode/n1162 ), .B1(n1304), .B2(
        \unit_decode/n3597 ), .ZN(\unit_decode/Areg/ffi_21/n5 ) );
  INV_X1 U3943 ( .A(\unit_decode/registerA[21] ), .ZN(\unit_decode/n1162 ) );
  OAI22_X1 U3944 ( .A1(n1292), .A2(\unit_decode/n1163 ), .B1(n1304), .B2(
        \unit_decode/n3596 ), .ZN(\unit_decode/Areg/ffi_22/n5 ) );
  INV_X1 U3945 ( .A(\unit_decode/registerA[22] ), .ZN(\unit_decode/n1163 ) );
  OAI22_X1 U3946 ( .A1(n1292), .A2(\unit_decode/n1164 ), .B1(n1304), .B2(
        \unit_decode/n3595 ), .ZN(\unit_decode/Areg/ffi_23/n5 ) );
  INV_X1 U3947 ( .A(\unit_decode/registerA[23] ), .ZN(\unit_decode/n1164 ) );
  OAI22_X1 U3948 ( .A1(n1292), .A2(\unit_decode/n1165 ), .B1(n1304), .B2(
        \unit_decode/n3594 ), .ZN(\unit_decode/Areg/ffi_24/n5 ) );
  INV_X1 U3949 ( .A(\unit_decode/registerA[24] ), .ZN(\unit_decode/n1165 ) );
  OAI22_X1 U3950 ( .A1(n1291), .A2(\unit_decode/n1166 ), .B1(n1303), .B2(
        \unit_decode/n3593 ), .ZN(\unit_decode/Areg/ffi_25/n5 ) );
  INV_X1 U3951 ( .A(\unit_decode/registerA[25] ), .ZN(\unit_decode/n1166 ) );
  OAI22_X1 U3952 ( .A1(n1291), .A2(\unit_decode/n1167 ), .B1(n1303), .B2(
        \unit_decode/n3592 ), .ZN(\unit_decode/Areg/ffi_26/n5 ) );
  INV_X1 U3953 ( .A(\unit_decode/registerA[26] ), .ZN(\unit_decode/n1167 ) );
  OAI22_X1 U3954 ( .A1(n1291), .A2(\unit_decode/n1168 ), .B1(n1303), .B2(
        \unit_decode/n3591 ), .ZN(\unit_decode/Areg/ffi_27/n5 ) );
  INV_X1 U3955 ( .A(\unit_decode/registerA[27] ), .ZN(\unit_decode/n1168 ) );
  OAI22_X1 U3956 ( .A1(n1291), .A2(\unit_decode/n1169 ), .B1(n1303), .B2(
        \unit_decode/n3590 ), .ZN(\unit_decode/Areg/ffi_28/n5 ) );
  INV_X1 U3957 ( .A(\unit_decode/registerA[28] ), .ZN(\unit_decode/n1169 ) );
  OAI22_X1 U3958 ( .A1(n1291), .A2(\unit_decode/n1170 ), .B1(n1303), .B2(
        \unit_decode/n3589 ), .ZN(\unit_decode/Areg/ffi_29/n5 ) );
  INV_X1 U3959 ( .A(\unit_decode/registerA[29] ), .ZN(\unit_decode/n1170 ) );
  OAI22_X1 U3960 ( .A1(n1291), .A2(\unit_decode/n1171 ), .B1(n1303), .B2(
        \unit_decode/n3588 ), .ZN(\unit_decode/Areg/ffi_30/n5 ) );
  INV_X1 U3961 ( .A(\unit_decode/registerA[30] ), .ZN(\unit_decode/n1171 ) );
  OAI22_X1 U3962 ( .A1(n1291), .A2(\unit_decode/n1172 ), .B1(n1303), .B2(
        \unit_decode/n3587 ), .ZN(\unit_decode/Areg/ffi_31/n5 ) );
  INV_X1 U3963 ( .A(\unit_decode/registerA[31] ), .ZN(\unit_decode/n1172 ) );
  OAI22_X1 U3964 ( .A1(n1288), .A2(n70), .B1(\unit_decode/n201 ), .B2(n1299), 
        .ZN(\unit_decode/NPC1reg/ffi_0/n5 ) );
  OAI22_X1 U3965 ( .A1(n1287), .A2(\unit_decode/n2147 ), .B1(
        \unit_decode/n205 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_1/n5 )
         );
  OAI22_X1 U3966 ( .A1(n1287), .A2(\unit_decode/n2146 ), .B1(
        \unit_decode/n195 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_2/n5 )
         );
  OAI22_X1 U3967 ( .A1(n1286), .A2(\unit_decode/n2145 ), .B1(
        \unit_decode/n217 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_3/n5 )
         );
  OAI22_X1 U3968 ( .A1(n1285), .A2(\unit_decode/n2144 ), .B1(
        \unit_decode/n3586 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_4/n5 )
         );
  OAI22_X1 U3969 ( .A1(n1285), .A2(\unit_decode/n2143 ), .B1(
        \unit_decode/n3585 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_5/n5 )
         );
  OAI22_X1 U3970 ( .A1(n1285), .A2(\unit_decode/n2142 ), .B1(
        \unit_decode/n3584 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_6/n5 )
         );
  OAI22_X1 U3971 ( .A1(n1285), .A2(\unit_decode/n2141 ), .B1(
        \unit_decode/n3583 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_7/n5 )
         );
  OAI22_X1 U3972 ( .A1(n1285), .A2(\unit_decode/n2140 ), .B1(
        \unit_decode/n3582 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_8/n5 )
         );
  OAI22_X1 U3973 ( .A1(n1285), .A2(\unit_decode/n2139 ), .B1(
        \unit_decode/n3581 ), .B2(n1296), .ZN(\unit_decode/NPC1reg/ffi_9/n5 )
         );
  OAI22_X1 U3974 ( .A1(n1287), .A2(\unit_decode/n2138 ), .B1(
        \unit_decode/n3580 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_10/n5 )
         );
  OAI22_X1 U3975 ( .A1(n1287), .A2(\unit_decode/n2137 ), .B1(
        \unit_decode/n3579 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_11/n5 )
         );
  OAI22_X1 U3976 ( .A1(n1287), .A2(\unit_decode/n2136 ), .B1(
        \unit_decode/n3578 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_12/n5 )
         );
  OAI22_X1 U3977 ( .A1(n1287), .A2(\unit_decode/n2135 ), .B1(
        \unit_decode/n3577 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_13/n5 )
         );
  OAI22_X1 U3978 ( .A1(n1287), .A2(\unit_decode/n2134 ), .B1(
        \unit_decode/n3576 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_14/n5 )
         );
  OAI22_X1 U3979 ( .A1(n1287), .A2(\unit_decode/n2133 ), .B1(
        \unit_decode/n3575 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_15/n5 )
         );
  OAI22_X1 U3980 ( .A1(n1287), .A2(\unit_decode/n2132 ), .B1(
        \unit_decode/n3574 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_16/n5 )
         );
  OAI22_X1 U3981 ( .A1(n1287), .A2(\unit_decode/n2131 ), .B1(
        \unit_decode/n3573 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_17/n5 )
         );
  OAI22_X1 U3982 ( .A1(n1287), .A2(\unit_decode/n2130 ), .B1(
        \unit_decode/n3572 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_18/n5 )
         );
  OAI22_X1 U3983 ( .A1(n1287), .A2(\unit_decode/n2129 ), .B1(
        \unit_decode/n3571 ), .B2(n1298), .ZN(\unit_decode/NPC1reg/ffi_19/n5 )
         );
  OAI22_X1 U3984 ( .A1(n1286), .A2(\unit_decode/n2128 ), .B1(
        \unit_decode/n3570 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_20/n5 )
         );
  OAI22_X1 U3985 ( .A1(n1286), .A2(\unit_decode/n2127 ), .B1(
        \unit_decode/n3569 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_21/n5 )
         );
  OAI22_X1 U3986 ( .A1(n1286), .A2(\unit_decode/n2126 ), .B1(
        \unit_decode/n3568 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_22/n5 )
         );
  OAI22_X1 U3987 ( .A1(n1286), .A2(\unit_decode/n2125 ), .B1(
        \unit_decode/n3567 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_23/n5 )
         );
  OAI22_X1 U3988 ( .A1(n1286), .A2(\unit_decode/n2124 ), .B1(
        \unit_decode/n3566 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_24/n5 )
         );
  OAI22_X1 U3989 ( .A1(n1286), .A2(\unit_decode/n2123 ), .B1(
        \unit_decode/n3565 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_25/n5 )
         );
  OAI22_X1 U3990 ( .A1(n1286), .A2(\unit_decode/n2122 ), .B1(
        \unit_decode/n3564 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_26/n5 )
         );
  OAI22_X1 U3991 ( .A1(n1286), .A2(\unit_decode/n2121 ), .B1(
        \unit_decode/n3563 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_27/n5 )
         );
  OAI22_X1 U3992 ( .A1(n1286), .A2(\unit_decode/n2120 ), .B1(
        \unit_decode/n3562 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_28/n5 )
         );
  OAI22_X1 U3993 ( .A1(n1286), .A2(\unit_decode/n2119 ), .B1(
        \unit_decode/n3561 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_29/n5 )
         );
  OAI22_X1 U3994 ( .A1(n1286), .A2(\unit_decode/n2118 ), .B1(
        \unit_decode/n3560 ), .B2(n1297), .ZN(\unit_decode/NPC1reg/ffi_30/n5 )
         );
  OAI22_X1 U3995 ( .A1(\unit_memory/DRAM/n3359 ), .A2(n692), .B1(n249), .B2(
        n698), .ZN(\unit_memory/DRAM/n1188 ) );
  OAI22_X1 U3996 ( .A1(\unit_memory/DRAM/n3360 ), .A2(n692), .B1(n266), .B2(
        n694), .ZN(\unit_memory/DRAM/n1187 ) );
  OAI22_X1 U3997 ( .A1(\unit_memory/DRAM/n3361 ), .A2(n692), .B1(n269), .B2(
        n694), .ZN(\unit_memory/DRAM/n1186 ) );
  OAI22_X1 U3998 ( .A1(\unit_memory/DRAM/n3362 ), .A2(n692), .B1(n272), .B2(
        n694), .ZN(\unit_memory/DRAM/n1185 ) );
  OAI22_X1 U3999 ( .A1(\unit_memory/DRAM/n3363 ), .A2(n692), .B1(n275), .B2(
        n695), .ZN(\unit_memory/DRAM/n1184 ) );
  OAI22_X1 U4000 ( .A1(\unit_memory/DRAM/n3364 ), .A2(n692), .B1(n278), .B2(
        n695), .ZN(\unit_memory/DRAM/n1183 ) );
  OAI22_X1 U4001 ( .A1(\unit_memory/DRAM/n3365 ), .A2(n692), .B1(n281), .B2(
        n695), .ZN(\unit_memory/DRAM/n1182 ) );
  OAI22_X1 U4002 ( .A1(\unit_memory/DRAM/n3366 ), .A2(n692), .B1(n284), .B2(
        n695), .ZN(\unit_memory/DRAM/n1181 ) );
  OAI22_X1 U4003 ( .A1(\unit_memory/DRAM/n3367 ), .A2(n692), .B1(n287), .B2(
        n696), .ZN(\unit_memory/DRAM/n1180 ) );
  OAI22_X1 U4004 ( .A1(\unit_memory/DRAM/n3368 ), .A2(n692), .B1(n290), .B2(
        n696), .ZN(\unit_memory/DRAM/n1179 ) );
  OAI22_X1 U4005 ( .A1(\unit_memory/DRAM/n3369 ), .A2(n692), .B1(n293), .B2(
        n696), .ZN(\unit_memory/DRAM/n1178 ) );
  OAI22_X1 U4006 ( .A1(\unit_memory/DRAM/n3370 ), .A2(n692), .B1(n296), .B2(
        n696), .ZN(\unit_memory/DRAM/n1177 ) );
  OAI22_X1 U4007 ( .A1(\unit_memory/DRAM/n3371 ), .A2(n693), .B1(n299), .B2(
        n697), .ZN(\unit_memory/DRAM/n1176 ) );
  OAI22_X1 U4008 ( .A1(\unit_memory/DRAM/n3372 ), .A2(n693), .B1(n302), .B2(
        n697), .ZN(\unit_memory/DRAM/n1175 ) );
  OAI22_X1 U4009 ( .A1(\unit_memory/DRAM/n3373 ), .A2(n693), .B1(n305), .B2(
        n697), .ZN(\unit_memory/DRAM/n1174 ) );
  OAI22_X1 U4010 ( .A1(\unit_memory/DRAM/n3374 ), .A2(n693), .B1(n308), .B2(
        n697), .ZN(\unit_memory/DRAM/n1173 ) );
  OAI22_X1 U4011 ( .A1(\unit_memory/DRAM/n3375 ), .A2(n693), .B1(n311), .B2(
        n698), .ZN(\unit_memory/DRAM/n1172 ) );
  OAI22_X1 U4012 ( .A1(\unit_memory/DRAM/n3376 ), .A2(n693), .B1(n314), .B2(
        n698), .ZN(\unit_memory/DRAM/n1171 ) );
  OAI22_X1 U4013 ( .A1(\unit_memory/DRAM/n3377 ), .A2(n693), .B1(n317), .B2(
        n698), .ZN(\unit_memory/DRAM/n1170 ) );
  OAI22_X1 U4014 ( .A1(\unit_memory/DRAM/n3378 ), .A2(n693), .B1(n320), .B2(
        n699), .ZN(\unit_memory/DRAM/n1169 ) );
  OAI22_X1 U4015 ( .A1(\unit_memory/DRAM/n3379 ), .A2(n693), .B1(n323), .B2(
        n699), .ZN(\unit_memory/DRAM/n1168 ) );
  OAI22_X1 U4016 ( .A1(\unit_memory/DRAM/n3380 ), .A2(n693), .B1(n326), .B2(
        n699), .ZN(\unit_memory/DRAM/n1167 ) );
  OAI22_X1 U4017 ( .A1(\unit_memory/DRAM/n3381 ), .A2(n693), .B1(n329), .B2(
        n699), .ZN(\unit_memory/DRAM/n1166 ) );
  OAI22_X1 U4018 ( .A1(\unit_memory/DRAM/n3382 ), .A2(n693), .B1(n332), .B2(
        n700), .ZN(\unit_memory/DRAM/n1165 ) );
  OAI22_X1 U4019 ( .A1(\unit_memory/DRAM/n3383 ), .A2(n693), .B1(n335), .B2(
        n700), .ZN(\unit_memory/DRAM/n1164 ) );
  OAI22_X1 U4020 ( .A1(\unit_memory/DRAM/n3384 ), .A2(n693), .B1(n338), .B2(
        n700), .ZN(\unit_memory/DRAM/n1163 ) );
  OAI22_X1 U4021 ( .A1(\unit_memory/DRAM/n3385 ), .A2(n692), .B1(n341), .B2(
        n700), .ZN(\unit_memory/DRAM/n1162 ) );
  OAI22_X1 U4022 ( .A1(\unit_memory/DRAM/n3386 ), .A2(n693), .B1(n344), .B2(
        n701), .ZN(\unit_memory/DRAM/n1161 ) );
  OAI22_X1 U4023 ( .A1(\unit_memory/DRAM/n3387 ), .A2(n692), .B1(n347), .B2(
        n701), .ZN(\unit_memory/DRAM/n1160 ) );
  OAI22_X1 U4024 ( .A1(\unit_memory/DRAM/n3388 ), .A2(n693), .B1(n350), .B2(
        n701), .ZN(\unit_memory/DRAM/n1159 ) );
  OAI22_X1 U4025 ( .A1(\unit_memory/DRAM/n3389 ), .A2(n692), .B1(n353), .B2(
        n701), .ZN(\unit_memory/DRAM/n1158 ) );
  NAND2_X1 U4026 ( .A1(wr_data[19]), .A2(n1346), .ZN(\unit_decode/n2208 ) );
  NAND2_X1 U4027 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_19/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_19/Y1 ), .ZN(wr_data[19]) );
  NAND2_X1 U4028 ( .A1(n1309), .A2(npc2_out[19]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_19/Y1 ) );
  NAND2_X1 U4029 ( .A1(n1306), .A2(\unit_memory/wb_prime[19] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_19/Y2 ) );
  NAND2_X1 U4030 ( .A1(wr_data[17]), .A2(n1346), .ZN(\unit_decode/n2210 ) );
  NAND2_X1 U4031 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_17/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_17/Y1 ), .ZN(wr_data[17]) );
  NAND2_X1 U4032 ( .A1(n1309), .A2(npc2_out[17]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_17/Y1 ) );
  NAND2_X1 U4033 ( .A1(n1306), .A2(\unit_memory/wb_prime[17] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_17/Y2 ) );
  NAND2_X1 U4034 ( .A1(wr_data[16]), .A2(n1346), .ZN(\unit_decode/n2211 ) );
  NAND2_X1 U4035 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_16/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_16/Y1 ), .ZN(wr_data[16]) );
  NAND2_X1 U4036 ( .A1(n1310), .A2(npc2_out[16]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_16/Y1 ) );
  NAND2_X1 U4037 ( .A1(n1306), .A2(\unit_memory/wb_prime[16] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_16/Y2 ) );
  NAND2_X1 U4038 ( .A1(wr_data[15]), .A2(n1345), .ZN(\unit_decode/n2212 ) );
  NAND2_X1 U4039 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_15/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_15/Y1 ), .ZN(wr_data[15]) );
  NAND2_X1 U4040 ( .A1(n1310), .A2(npc2_out[15]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_15/Y1 ) );
  NAND2_X1 U4041 ( .A1(n1306), .A2(\unit_memory/wb_prime[15] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_15/Y2 ) );
  NAND2_X1 U4042 ( .A1(wr_data[14]), .A2(n1346), .ZN(\unit_decode/n2213 ) );
  NAND2_X1 U4043 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_14/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_14/Y1 ), .ZN(wr_data[14]) );
  NAND2_X1 U4044 ( .A1(n1310), .A2(npc2_out[14]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_14/Y1 ) );
  NAND2_X1 U4045 ( .A1(n1306), .A2(\unit_memory/wb_prime[14] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_14/Y2 ) );
  NAND2_X1 U4046 ( .A1(wr_data[13]), .A2(n1345), .ZN(\unit_decode/n2214 ) );
  NAND2_X1 U4047 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_13/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_13/Y1 ), .ZN(wr_data[13]) );
  NAND2_X1 U4048 ( .A1(n1310), .A2(npc2_out[13]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_13/Y1 ) );
  NAND2_X1 U4049 ( .A1(n1306), .A2(\unit_memory/wb_prime[13] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_13/Y2 ) );
  NAND2_X1 U4050 ( .A1(wr_data[12]), .A2(n1346), .ZN(\unit_decode/n2215 ) );
  NAND2_X1 U4051 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_12/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_12/Y1 ), .ZN(wr_data[12]) );
  NAND2_X1 U4052 ( .A1(n1310), .A2(npc2_out[12]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_12/Y1 ) );
  NAND2_X1 U4053 ( .A1(n1306), .A2(\unit_memory/wb_prime[12] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_12/Y2 ) );
  NAND2_X1 U4054 ( .A1(wr_data[11]), .A2(n1345), .ZN(\unit_decode/n2216 ) );
  NAND2_X1 U4055 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_11/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_11/Y1 ), .ZN(wr_data[11]) );
  NAND2_X1 U4056 ( .A1(n1311), .A2(npc2_out[11]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_11/Y1 ) );
  NAND2_X1 U4057 ( .A1(n33), .A2(\unit_memory/wb_prime[11] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_11/Y2 ) );
  NAND2_X1 U4058 ( .A1(wr_data[10]), .A2(n1346), .ZN(\unit_decode/n2217 ) );
  NAND2_X1 U4059 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_10/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_10/Y1 ), .ZN(wr_data[10]) );
  NAND2_X1 U4060 ( .A1(n1311), .A2(npc2_out[10]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_10/Y1 ) );
  NAND2_X1 U4061 ( .A1(n33), .A2(\unit_memory/wb_prime[10] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_10/Y2 ) );
  NAND2_X1 U4062 ( .A1(wr_data[9]), .A2(n1346), .ZN(\unit_decode/n2218 ) );
  NAND2_X1 U4063 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_9/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_9/Y1 ), .ZN(wr_data[9]) );
  NAND2_X1 U4064 ( .A1(n1311), .A2(npc2_out[9]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_9/Y1 ) );
  NAND2_X1 U4065 ( .A1(n33), .A2(\unit_memory/wb_prime[9] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_9/Y2 ) );
  NAND2_X1 U4066 ( .A1(wr_data[8]), .A2(n1346), .ZN(\unit_decode/n2219 ) );
  NAND2_X1 U4067 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_8/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_8/Y1 ), .ZN(wr_data[8]) );
  NAND2_X1 U4068 ( .A1(n1311), .A2(npc2_out[8]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_8/Y1 ) );
  NAND2_X1 U4069 ( .A1(n33), .A2(\unit_memory/wb_prime[8] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_8/Y2 ) );
  NAND2_X1 U4070 ( .A1(wr_data[7]), .A2(n1345), .ZN(\unit_decode/n2220 ) );
  NAND2_X1 U4071 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_7/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_7/Y1 ), .ZN(wr_data[7]) );
  NAND2_X1 U4072 ( .A1(n1311), .A2(npc2_out[7]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_7/Y1 ) );
  NAND2_X1 U4073 ( .A1(n33), .A2(\unit_memory/wb_prime[7] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_7/Y2 ) );
  NAND2_X1 U4074 ( .A1(wr_data[6]), .A2(n1346), .ZN(\unit_decode/n2221 ) );
  NAND2_X1 U4075 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_6/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_6/Y1 ), .ZN(wr_data[6]) );
  NAND2_X1 U4076 ( .A1(n1312), .A2(npc2_out[6]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_6/Y1 ) );
  NAND2_X1 U4077 ( .A1(n33), .A2(\unit_memory/wb_prime[6] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_6/Y2 ) );
  NAND2_X1 U4078 ( .A1(wr_data[5]), .A2(n1345), .ZN(\unit_decode/n2222 ) );
  NAND2_X1 U4079 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_5/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_5/Y1 ), .ZN(wr_data[5]) );
  NAND2_X1 U4080 ( .A1(n1312), .A2(npc2_out[5]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_5/Y1 ) );
  NAND2_X1 U4081 ( .A1(n33), .A2(\unit_memory/wb_prime[5] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_5/Y2 ) );
  NAND2_X1 U4082 ( .A1(wr_data[4]), .A2(n1345), .ZN(\unit_decode/n2223 ) );
  NAND2_X1 U4083 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_4/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_4/Y1 ), .ZN(wr_data[4]) );
  NAND2_X1 U4084 ( .A1(n1312), .A2(npc2_out[4]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_4/Y1 ) );
  NAND2_X1 U4085 ( .A1(n33), .A2(\unit_memory/wb_prime[4] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_4/Y2 ) );
  NAND2_X1 U4086 ( .A1(wr_data[3]), .A2(n1345), .ZN(\unit_decode/n2224 ) );
  NAND2_X1 U4087 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_3/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_3/Y1 ), .ZN(wr_data[3]) );
  NAND2_X1 U4088 ( .A1(n1312), .A2(npc2_out[3]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_3/Y1 ) );
  NAND2_X1 U4089 ( .A1(n33), .A2(\unit_memory/wb_prime[3] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_3/Y2 ) );
  NAND2_X1 U4090 ( .A1(wr_data[2]), .A2(n1345), .ZN(\unit_decode/n2225 ) );
  NAND2_X1 U4091 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_2/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_2/Y1 ), .ZN(wr_data[2]) );
  NAND2_X1 U4092 ( .A1(n1312), .A2(npc2_out[2]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_2/Y1 ) );
  NAND2_X1 U4093 ( .A1(n33), .A2(\unit_memory/wb_prime[2] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_2/Y2 ) );
  NAND2_X1 U4094 ( .A1(wr_data[23]), .A2(n1346), .ZN(\unit_decode/n2204 ) );
  NAND2_X1 U4095 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_23/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_23/Y1 ), .ZN(wr_data[23]) );
  NAND2_X1 U4096 ( .A1(n1308), .A2(npc2_out[23]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_23/Y1 ) );
  NAND2_X1 U4097 ( .A1(n1306), .A2(\unit_memory/wb_prime[23] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_23/Y2 ) );
  NAND2_X1 U4098 ( .A1(wr_data[22]), .A2(n1347), .ZN(\unit_decode/n2205 ) );
  NAND2_X1 U4099 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_22/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_22/Y1 ), .ZN(wr_data[22]) );
  NAND2_X1 U4100 ( .A1(n1308), .A2(npc2_out[22]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_22/Y1 ) );
  NAND2_X1 U4101 ( .A1(n1306), .A2(\unit_memory/wb_prime[22] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_22/Y2 ) );
  NAND2_X1 U4102 ( .A1(wr_data[21]), .A2(n1347), .ZN(\unit_decode/n2206 ) );
  NAND2_X1 U4103 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_21/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_21/Y1 ), .ZN(wr_data[21]) );
  NAND2_X1 U4104 ( .A1(n1309), .A2(npc2_out[21]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_21/Y1 ) );
  NAND2_X1 U4105 ( .A1(n1306), .A2(\unit_memory/wb_prime[21] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_21/Y2 ) );
  NAND2_X1 U4106 ( .A1(wr_data[20]), .A2(n1347), .ZN(\unit_decode/n2207 ) );
  NAND2_X1 U4107 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_20/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_20/Y1 ), .ZN(wr_data[20]) );
  NAND2_X1 U4108 ( .A1(n1309), .A2(npc2_out[20]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_20/Y1 ) );
  NAND2_X1 U4109 ( .A1(n1306), .A2(\unit_memory/wb_prime[20] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_20/Y2 ) );
  NAND2_X1 U4110 ( .A1(wr_data[18]), .A2(n1347), .ZN(\unit_decode/n2209 ) );
  NAND2_X1 U4111 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_18/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_18/Y1 ), .ZN(wr_data[18]) );
  NAND2_X1 U4112 ( .A1(n1309), .A2(npc2_out[18]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_18/Y1 ) );
  NAND2_X1 U4113 ( .A1(n1306), .A2(\unit_memory/wb_prime[18] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_18/Y2 ) );
  NAND2_X1 U4114 ( .A1(wr_data[31]), .A2(n1346), .ZN(\unit_decode/n2195 ) );
  NAND2_X1 U4115 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_31/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_31/Y1 ), .ZN(wr_data[31]) );
  NAND2_X1 U4116 ( .A1(n1307), .A2(npc2_out[31]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_31/Y1 ) );
  NAND2_X1 U4117 ( .A1(n33), .A2(\unit_memory/wb_prime[31] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_31/Y2 ) );
  NAND2_X1 U4118 ( .A1(wr_data[30]), .A2(n1347), .ZN(\unit_decode/n2197 ) );
  NAND2_X1 U4119 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_30/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_30/Y1 ), .ZN(wr_data[30]) );
  NAND2_X1 U4120 ( .A1(n1307), .A2(npc2_out[30]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_30/Y1 ) );
  NAND2_X1 U4121 ( .A1(n33), .A2(\unit_memory/wb_prime[30] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_30/Y2 ) );
  NAND2_X1 U4122 ( .A1(wr_data[29]), .A2(n1347), .ZN(\unit_decode/n2198 ) );
  NAND2_X1 U4123 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_29/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_29/Y1 ), .ZN(wr_data[29]) );
  NAND2_X1 U4124 ( .A1(n1307), .A2(npc2_out[29]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_29/Y1 ) );
  NAND2_X1 U4125 ( .A1(n33), .A2(\unit_memory/wb_prime[29] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_29/Y2 ) );
  NAND2_X1 U4126 ( .A1(wr_data[28]), .A2(n1347), .ZN(\unit_decode/n2199 ) );
  NAND2_X1 U4127 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_28/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_28/Y1 ), .ZN(wr_data[28]) );
  NAND2_X1 U4128 ( .A1(n1307), .A2(npc2_out[28]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_28/Y1 ) );
  NAND2_X1 U4129 ( .A1(n33), .A2(\unit_memory/wb_prime[28] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_28/Y2 ) );
  NAND2_X1 U4130 ( .A1(wr_data[27]), .A2(n1346), .ZN(\unit_decode/n2200 ) );
  NAND2_X1 U4131 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_27/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_27/Y1 ), .ZN(wr_data[27]) );
  NAND2_X1 U4132 ( .A1(n1307), .A2(npc2_out[27]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_27/Y1 ) );
  NAND2_X1 U4133 ( .A1(n33), .A2(\unit_memory/wb_prime[27] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_27/Y2 ) );
  NAND2_X1 U4134 ( .A1(wr_data[26]), .A2(n1347), .ZN(\unit_decode/n2201 ) );
  NAND2_X1 U4135 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_26/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_26/Y1 ), .ZN(wr_data[26]) );
  NAND2_X1 U4136 ( .A1(n1308), .A2(npc2_out[26]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_26/Y1 ) );
  NAND2_X1 U4137 ( .A1(n33), .A2(\unit_memory/wb_prime[26] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_26/Y2 ) );
  NAND2_X1 U4138 ( .A1(wr_data[25]), .A2(n1347), .ZN(\unit_decode/n2202 ) );
  NAND2_X1 U4139 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_25/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_25/Y1 ), .ZN(wr_data[25]) );
  NAND2_X1 U4140 ( .A1(n1308), .A2(npc2_out[25]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_25/Y1 ) );
  NAND2_X1 U4141 ( .A1(n33), .A2(\unit_memory/wb_prime[25] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_25/Y2 ) );
  NAND2_X1 U4142 ( .A1(wr_data[24]), .A2(n1347), .ZN(\unit_decode/n2203 ) );
  NAND2_X1 U4143 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_24/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_24/Y1 ), .ZN(wr_data[24]) );
  NAND2_X1 U4144 ( .A1(n1308), .A2(npc2_out[24]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_24/Y1 ) );
  NAND2_X1 U4145 ( .A1(n33), .A2(\unit_memory/wb_prime[24] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_24/Y2 ) );
  BUF_X1 U4146 ( .A(cw_mem[6]), .Z(n1317) );
  BUF_X1 U4147 ( .A(cw_mem[6]), .Z(n1318) );
  BUF_X1 U4148 ( .A(cw_mem[6]), .Z(n1319) );
  BUF_X1 U4149 ( .A(cw_mem[6]), .Z(n1320) );
  BUF_X1 U4150 ( .A(cw_mem[6]), .Z(n1315) );
  BUF_X1 U4151 ( .A(cw_mem[6]), .Z(n1316) );
  BUF_X1 U4152 ( .A(cw_mem[3]), .Z(n1307) );
  BUF_X1 U4153 ( .A(cw_mem[3]), .Z(n1309) );
  BUF_X1 U4154 ( .A(cw_mem[3]), .Z(n1310) );
  BUF_X1 U4155 ( .A(cw_mem[3]), .Z(n1311) );
  BUF_X1 U4156 ( .A(cw_mem[3]), .Z(n1312) );
  BUF_X1 U4157 ( .A(cw_mem[3]), .Z(n1308) );
  BUF_X1 U4158 ( .A(cw_mem[6]), .Z(n1321) );
  BUF_X1 U4159 ( .A(cw_mem[3]), .Z(n1313) );
  NAND2_X1 U4160 ( .A1(\unit_fetch/pc_regout[4] ), .A2(n1697), .ZN(
        \unit_fetch/n682 ) );
  NAND2_X1 U4161 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_2/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_2/Y1 ), .ZN(
        \unit_memory/wb_prime[2] ) );
  NAND2_X1 U4162 ( .A1(n1321), .A2(\unit_memory/DataMemOut[2] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_2/Y1 ) );
  NAND2_X1 U4163 ( .A1(n1314), .A2(aluout_regn[2]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_2/Y2 ) );
  NAND2_X1 U4164 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_24/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_24/Y1 ), .ZN(
        \unit_memory/wb_prime[24] ) );
  NAND2_X1 U4165 ( .A1(n1316), .A2(\unit_memory/DataMemOut[24] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_24/Y1 ) );
  NAND2_X1 U4166 ( .A1(n34), .A2(aluout_regn[24]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_24/Y2 ) );
  NAND2_X1 U4167 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_22/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_22/Y1 ), .ZN(
        \unit_memory/wb_prime[22] ) );
  NAND2_X1 U4168 ( .A1(n1317), .A2(\unit_memory/DataMemOut[22] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_22/Y1 ) );
  NAND2_X1 U4169 ( .A1(n34), .A2(aluout_regn[22]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_22/Y2 ) );
  NAND2_X1 U4170 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_21/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_21/Y1 ), .ZN(
        \unit_memory/wb_prime[21] ) );
  NAND2_X1 U4171 ( .A1(n1317), .A2(\unit_memory/DataMemOut[21] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_21/Y1 ) );
  NAND2_X1 U4172 ( .A1(n34), .A2(aluout_regn[21]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_21/Y2 ) );
  NAND2_X1 U4173 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_20/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_20/Y1 ), .ZN(
        \unit_memory/wb_prime[20] ) );
  NAND2_X1 U4174 ( .A1(n1317), .A2(\unit_memory/DataMemOut[20] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_20/Y1 ) );
  NAND2_X1 U4175 ( .A1(n34), .A2(aluout_regn[20]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_20/Y2 ) );
  NAND2_X1 U4176 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_19/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_19/Y1 ), .ZN(
        \unit_memory/wb_prime[19] ) );
  NAND2_X1 U4177 ( .A1(n1317), .A2(\unit_memory/DataMemOut[19] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_19/Y1 ) );
  NAND2_X1 U4178 ( .A1(n34), .A2(aluout_regn[19]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_19/Y2 ) );
  NAND2_X1 U4179 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_18/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_18/Y1 ), .ZN(
        \unit_memory/wb_prime[18] ) );
  NAND2_X1 U4180 ( .A1(n1317), .A2(\unit_memory/DataMemOut[18] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_18/Y1 ) );
  NAND2_X1 U4181 ( .A1(n34), .A2(aluout_regn[18]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_18/Y2 ) );
  NAND2_X1 U4182 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_17/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_17/Y1 ), .ZN(
        \unit_memory/wb_prime[17] ) );
  NAND2_X1 U4183 ( .A1(n1318), .A2(\unit_memory/DataMemOut[17] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_17/Y1 ) );
  NAND2_X1 U4184 ( .A1(n34), .A2(aluout_regn[17]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_17/Y2 ) );
  NAND2_X1 U4185 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_16/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_16/Y1 ), .ZN(
        \unit_memory/wb_prime[16] ) );
  NAND2_X1 U4186 ( .A1(n1318), .A2(\unit_memory/DataMemOut[16] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_16/Y1 ) );
  NAND2_X1 U4187 ( .A1(n34), .A2(aluout_regn[16]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_16/Y2 ) );
  NAND2_X1 U4188 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_15/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_15/Y1 ), .ZN(
        \unit_memory/wb_prime[15] ) );
  NAND2_X1 U4189 ( .A1(n1318), .A2(\unit_memory/DataMemOut[15] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_15/Y1 ) );
  NAND2_X1 U4190 ( .A1(n34), .A2(aluout_regn[15]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_15/Y2 ) );
  NAND2_X1 U4191 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_14/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_14/Y1 ), .ZN(
        \unit_memory/wb_prime[14] ) );
  NAND2_X1 U4192 ( .A1(n1318), .A2(\unit_memory/DataMemOut[14] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_14/Y1 ) );
  NAND2_X1 U4193 ( .A1(n34), .A2(aluout_regn[14]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_14/Y2 ) );
  NAND2_X1 U4194 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_13/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_13/Y1 ), .ZN(
        \unit_memory/wb_prime[13] ) );
  NAND2_X1 U4195 ( .A1(n1318), .A2(\unit_memory/DataMemOut[13] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_13/Y1 ) );
  NAND2_X1 U4196 ( .A1(n34), .A2(aluout_regn[13]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_13/Y2 ) );
  NAND2_X1 U4197 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_12/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_12/Y1 ), .ZN(
        \unit_memory/wb_prime[12] ) );
  NAND2_X1 U4198 ( .A1(n1319), .A2(\unit_memory/DataMemOut[12] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_12/Y1 ) );
  NAND2_X1 U4199 ( .A1(n1314), .A2(aluout_regn[12]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_12/Y2 ) );
  NAND2_X1 U4200 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_11/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_11/Y1 ), .ZN(
        \unit_memory/wb_prime[11] ) );
  NAND2_X1 U4201 ( .A1(n1319), .A2(\unit_memory/DataMemOut[11] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_11/Y1 ) );
  NAND2_X1 U4202 ( .A1(n1314), .A2(aluout_regn[11]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_11/Y2 ) );
  NAND2_X1 U4203 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_10/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_10/Y1 ), .ZN(
        \unit_memory/wb_prime[10] ) );
  NAND2_X1 U4204 ( .A1(n1319), .A2(\unit_memory/DataMemOut[10] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_10/Y1 ) );
  NAND2_X1 U4205 ( .A1(n1314), .A2(aluout_regn[10]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_10/Y2 ) );
  NAND2_X1 U4206 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_9/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_9/Y1 ), .ZN(
        \unit_memory/wb_prime[9] ) );
  NAND2_X1 U4207 ( .A1(n1319), .A2(\unit_memory/DataMemOut[9] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_9/Y1 ) );
  NAND2_X1 U4208 ( .A1(n1314), .A2(aluout_regn[9]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_9/Y2 ) );
  NAND2_X1 U4209 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_8/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_8/Y1 ), .ZN(
        \unit_memory/wb_prime[8] ) );
  NAND2_X1 U4210 ( .A1(n1319), .A2(\unit_memory/DataMemOut[8] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_8/Y1 ) );
  NAND2_X1 U4211 ( .A1(n1314), .A2(aluout_regn[8]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_8/Y2 ) );
  NAND2_X1 U4212 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_7/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_7/Y1 ), .ZN(
        \unit_memory/wb_prime[7] ) );
  NAND2_X1 U4213 ( .A1(n1320), .A2(\unit_memory/DataMemOut[7] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_7/Y1 ) );
  NAND2_X1 U4214 ( .A1(n1314), .A2(aluout_regn[7]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_7/Y2 ) );
  NAND2_X1 U4215 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_6/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_6/Y1 ), .ZN(
        \unit_memory/wb_prime[6] ) );
  NAND2_X1 U4216 ( .A1(n1320), .A2(\unit_memory/DataMemOut[6] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_6/Y1 ) );
  NAND2_X1 U4217 ( .A1(n1314), .A2(aluout_regn[6]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_6/Y2 ) );
  NAND2_X1 U4218 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_5/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_5/Y1 ), .ZN(
        \unit_memory/wb_prime[5] ) );
  NAND2_X1 U4219 ( .A1(n1320), .A2(\unit_memory/DataMemOut[5] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_5/Y1 ) );
  NAND2_X1 U4220 ( .A1(n1314), .A2(aluout_regn[5]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_5/Y2 ) );
  NAND2_X1 U4221 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_4/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_4/Y1 ), .ZN(
        \unit_memory/wb_prime[4] ) );
  NAND2_X1 U4222 ( .A1(n1320), .A2(\unit_memory/DataMemOut[4] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_4/Y1 ) );
  NAND2_X1 U4223 ( .A1(n1314), .A2(aluout_regn[4]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_4/Y2 ) );
  NAND2_X1 U4224 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_3/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_3/Y1 ), .ZN(
        \unit_memory/wb_prime[3] ) );
  NAND2_X1 U4225 ( .A1(n1320), .A2(\unit_memory/DataMemOut[3] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_3/Y1 ) );
  NAND2_X1 U4226 ( .A1(n1314), .A2(aluout_regn[3]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_3/Y2 ) );
  NAND2_X1 U4227 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_1/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_1/Y1 ), .ZN(
        \unit_memory/wb_prime[1] ) );
  NAND2_X1 U4228 ( .A1(n1321), .A2(\unit_memory/DataMemOut[1] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_1/Y1 ) );
  NAND2_X1 U4229 ( .A1(n1314), .A2(aluout_regn[1]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_1/Y2 ) );
  NAND2_X1 U4230 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_23/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_23/Y1 ), .ZN(
        \unit_memory/wb_prime[23] ) );
  NAND2_X1 U4231 ( .A1(n1316), .A2(\unit_memory/DataMemOut[23] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_23/Y1 ) );
  NAND2_X1 U4232 ( .A1(n34), .A2(aluout_regn[23]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_23/Y2 ) );
  INV_X1 U4233 ( .A(wr_address[2]), .ZN(\unit_decode/n2183 ) );
  INV_X1 U4234 ( .A(wr_address[0]), .ZN(\unit_decode/n2185 ) );
  INV_X1 U4235 ( .A(wr_address[1]), .ZN(\unit_decode/n2184 ) );
  INV_X1 U4236 ( .A(aluout_regn[0]), .ZN(\unit_memory/DRAM/n552 ) );
  OAI21_X1 U4237 ( .B1(\unit_decode/n3603 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_26/n5 ) );
  OAI21_X1 U4238 ( .B1(\unit_decode/n3602 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_27/n5 ) );
  OAI21_X1 U4239 ( .B1(\unit_decode/n3559 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_28/n5 ) );
  OAI21_X1 U4240 ( .B1(\unit_decode/n3601 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_29/n5 ) );
  OAI21_X1 U4241 ( .B1(\unit_decode/n3600 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_30/n5 ) );
  OAI21_X1 U4242 ( .B1(\unit_decode/n3625 ), .B2(n1299), .A(
        \unit_decode/n3519 ), .ZN(\unit_decode/IMMreg/ffi_31/n5 ) );
  NOR2_X1 U4243 ( .A1(n108), .A2(n109), .ZN(\unit_memory/DRAM/n771 ) );
  AND2_X1 U4244 ( .A1(cw_mem[4]), .A2(n135), .ZN(\unit_decode/n2244 ) );
  AND2_X1 U4245 ( .A1(aluout_regn[4]), .A2(\unit_memory/DRAM/n546 ), .ZN(
        \unit_memory/DRAM/n792 ) );
  AND2_X1 U4246 ( .A1(aluout_regn[4]), .A2(aluout_regn[3]), .ZN(
        \unit_memory/DRAM/n809 ) );
  AND2_X1 U4247 ( .A1(\unit_fetch/pc_regout[2] ), .A2(n36), .ZN(n111) );
  NOR2_X1 U4248 ( .A1(n1333), .A2(\unit_control/n385 ), .ZN(
        \unit_control/uut_third_stage/ffi_15/n5 ) );
  NOR2_X1 U4249 ( .A1(n1333), .A2(\unit_control/n391 ), .ZN(
        \unit_control/uut_third_stage/ffi_5/n5 ) );
  NOR2_X1 U4250 ( .A1(n1333), .A2(\unit_control/n393 ), .ZN(
        \unit_control/uut_third_stage/ffi_3/n5 ) );
  NOR2_X1 U4251 ( .A1(n1337), .A2(\unit_control/n387 ), .ZN(
        \unit_control/uut_third_stage/ffi_13/n5 ) );
  NOR2_X1 U4252 ( .A1(n1333), .A2(\unit_control/n378 ), .ZN(
        \unit_control/uut_third_stage/ffi_11/n5 ) );
  NOR2_X1 U4253 ( .A1(\unit_control/uut_third_stage/ffi_19/n2 ), .A2(n1328), 
        .ZN(\unit_control/uut_third_stage/ffi_19/n6 ) );
  NOR2_X1 U4254 ( .A1(\unit_control/uut_third_stage/ffi_17/n2 ), .A2(n1328), 
        .ZN(\unit_control/uut_third_stage/ffi_17/n6 ) );
  NOR2_X1 U4255 ( .A1(\unit_control/uut_third_stage/ffi_12/n2 ), .A2(n1327), 
        .ZN(\unit_control/uut_third_stage/ffi_12/n5 ) );
  NOR2_X1 U4256 ( .A1(n1329), .A2(\unit_control/n398 ), .ZN(
        \unit_control/uut_fourth_stage/ffi_7/n5 ) );
  NOR2_X1 U4257 ( .A1(n1329), .A2(\unit_control/n399 ), .ZN(
        \unit_control/uut_fourth_stage/ffi_5/n5 ) );
  NOR2_X1 U4258 ( .A1(n1329), .A2(\unit_control/n383 ), .ZN(
        \unit_control/uut_fourth_stage/ffi_3/n6 ) );
  NOR2_X1 U4259 ( .A1(n1334), .A2(\unit_control/n381 ), .ZN(
        \unit_control/uut_third_stage/ffi_9/n6 ) );
  NOR2_X1 U4260 ( .A1(n1330), .A2(\unit_control/n386 ), .ZN(
        \unit_control/uut_third_stage/ffi_14/n5 ) );
  NOR2_X1 U4261 ( .A1(n1334), .A2(\unit_control/n389 ), .ZN(
        \unit_control/uut_third_stage/ffi_7/n5 ) );
  NOR2_X1 U4262 ( .A1(n1331), .A2(\unit_control/n390 ), .ZN(
        \unit_control/uut_third_stage/ffi_6/n5 ) );
  NOR2_X1 U4263 ( .A1(n1331), .A2(\unit_control/n392 ), .ZN(
        \unit_control/uut_third_stage/ffi_4/n5 ) );
  NOR2_X1 U4264 ( .A1(n1332), .A2(\unit_control/n382 ), .ZN(
        \unit_control/uut_fourth_stage/ffi_6/n6 ) );
  NOR2_X1 U4265 ( .A1(n1332), .A2(\unit_control/n400 ), .ZN(
        \unit_control/uut_fourth_stage/ffi_4/n5 ) );
  NOR2_X1 U4266 ( .A1(n1330), .A2(\unit_control/n379 ), .ZN(
        \unit_control/uut_third_stage/ffi_10/n5 ) );
  INV_X1 U4267 ( .A(aluout_regn[3]), .ZN(\unit_memory/DRAM/n546 ) );
  NAND2_X1 U4268 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_31/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_31/Y1 ), .ZN(
        \unit_memory/wb_prime[31] ) );
  NAND2_X1 U4269 ( .A1(n1315), .A2(\unit_memory/DataMemOut[31] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_31/Y1 ) );
  NAND2_X1 U4270 ( .A1(n34), .A2(aluout_regn[31]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_31/Y2 ) );
  NAND2_X1 U4271 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_30/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_30/Y1 ), .ZN(
        \unit_memory/wb_prime[30] ) );
  NAND2_X1 U4272 ( .A1(n1315), .A2(\unit_memory/DataMemOut[30] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_30/Y1 ) );
  NAND2_X1 U4273 ( .A1(n34), .A2(aluout_regn[30]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_30/Y2 ) );
  NAND2_X1 U4274 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_29/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_29/Y1 ), .ZN(
        \unit_memory/wb_prime[29] ) );
  NAND2_X1 U4275 ( .A1(n1315), .A2(\unit_memory/DataMemOut[29] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_29/Y1 ) );
  NAND2_X1 U4276 ( .A1(n34), .A2(aluout_regn[29]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_29/Y2 ) );
  NAND2_X1 U4277 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_28/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_28/Y1 ), .ZN(
        \unit_memory/wb_prime[28] ) );
  NAND2_X1 U4278 ( .A1(n1315), .A2(\unit_memory/DataMemOut[28] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_28/Y1 ) );
  NAND2_X1 U4279 ( .A1(n34), .A2(aluout_regn[28]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_28/Y2 ) );
  NAND2_X1 U4280 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_27/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_27/Y1 ), .ZN(
        \unit_memory/wb_prime[27] ) );
  NAND2_X1 U4281 ( .A1(n1316), .A2(\unit_memory/DataMemOut[27] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_27/Y1 ) );
  NAND2_X1 U4282 ( .A1(n34), .A2(aluout_regn[27]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_27/Y2 ) );
  NAND2_X1 U4283 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_26/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_26/Y1 ), .ZN(
        \unit_memory/wb_prime[26] ) );
  NAND2_X1 U4284 ( .A1(n1316), .A2(\unit_memory/DataMemOut[26] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_26/Y1 ) );
  NAND2_X1 U4285 ( .A1(n34), .A2(aluout_regn[26]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_26/Y2 ) );
  NAND2_X1 U4286 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_25/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_25/Y1 ), .ZN(
        \unit_memory/wb_prime[25] ) );
  NAND2_X1 U4287 ( .A1(n1316), .A2(\unit_memory/DataMemOut[25] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_25/Y1 ) );
  NAND2_X1 U4288 ( .A1(n34), .A2(aluout_regn[25]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_25/Y2 ) );
  NAND2_X1 U4289 ( .A1(\unit_memory/MUX21_ALMEM/MUX21GENI_0/Y2 ), .A2(
        \unit_memory/MUX21_ALMEM/MUX21GENI_0/Y1 ), .ZN(
        \unit_memory/wb_prime[0] ) );
  NAND2_X1 U4290 ( .A1(n1315), .A2(\unit_memory/DataMemOut[0] ), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_0/Y1 ) );
  NAND2_X1 U4291 ( .A1(n34), .A2(aluout_regn[0]), .ZN(
        \unit_memory/MUX21_ALMEM/MUX21GENI_0/Y2 ) );
  INV_X1 U4292 ( .A(wr_address[4]), .ZN(\unit_decode/n2165 ) );
  INV_X1 U4293 ( .A(wr_address[3]), .ZN(\unit_decode/n2182 ) );
  OR2_X1 U4294 ( .A1(n1647), .A2(n1697), .ZN(n1498) );
  NAND2_X1 U4295 ( .A1(wr_data[1]), .A2(n1345), .ZN(\unit_decode/n2226 ) );
  NAND2_X1 U4296 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_1/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_1/Y1 ), .ZN(wr_data[1]) );
  NAND2_X1 U4297 ( .A1(n1313), .A2(npc2_out[1]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_1/Y1 ) );
  NAND2_X1 U4298 ( .A1(n33), .A2(\unit_memory/wb_prime[1] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_1/Y2 ) );
  NAND2_X1 U4299 ( .A1(wr_data[0]), .A2(n1345), .ZN(\unit_decode/n2227 ) );
  NAND2_X1 U4300 ( .A1(\unit_memory/MUX21_NPCWB/MUX21GENI_0/Y2 ), .A2(
        \unit_memory/MUX21_NPCWB/MUX21GENI_0/Y1 ), .ZN(wr_data[0]) );
  NAND2_X1 U4301 ( .A1(n1313), .A2(npc2_out[0]), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_0/Y1 ) );
  NAND2_X1 U4302 ( .A1(n33), .A2(\unit_memory/wb_prime[0] ), .ZN(
        \unit_memory/MUX21_NPCWB/MUX21GENI_0/Y2 ) );
  NOR3_X1 U4303 ( .A1(IR_OUT[24]), .A2(IR_OUT[25]), .A3(\unit_decode/n2093 ), 
        .ZN(\unit_decode/n3489 ) );
  NOR3_X1 U4304 ( .A1(\unit_decode/n2093 ), .A2(IR_OUT[25]), .A3(
        \unit_decode/n2092 ), .ZN(\unit_decode/n3495 ) );
  NOR3_X1 U4305 ( .A1(IR_OUT[24]), .A2(IR_OUT[25]), .A3(IR_OUT[23]), .ZN(
        \unit_decode/n3505 ) );
  NOR3_X1 U4306 ( .A1(IR_OUT[23]), .A2(IR_OUT[25]), .A3(\unit_decode/n2092 ), 
        .ZN(\unit_decode/n3507 ) );
  NOR3_X1 U4307 ( .A1(IR_OUT[19]), .A2(IR_OUT[20]), .A3(\unit_decode/n2098 ), 
        .ZN(\unit_decode/n2869 ) );
  NOR3_X1 U4308 ( .A1(\unit_decode/n2098 ), .A2(IR_OUT[20]), .A3(
        \unit_decode/n2097 ), .ZN(\unit_decode/n2875 ) );
  NOR3_X1 U4309 ( .A1(\unit_decode/n2098 ), .A2(IR_OUT[19]), .A3(
        \unit_decode/n2096 ), .ZN(\unit_decode/n2877 ) );
  NOR3_X1 U4310 ( .A1(IR_OUT[19]), .A2(IR_OUT[20]), .A3(IR_OUT[18]), .ZN(
        \unit_decode/n2885 ) );
  NOR3_X1 U4311 ( .A1(IR_OUT[18]), .A2(IR_OUT[20]), .A3(\unit_decode/n2097 ), 
        .ZN(\unit_decode/n2887 ) );
  NOR3_X1 U4312 ( .A1(IR_OUT[18]), .A2(IR_OUT[19]), .A3(\unit_decode/n2096 ), 
        .ZN(\unit_decode/n2889 ) );
  NOR3_X1 U4313 ( .A1(\unit_decode/n2097 ), .A2(IR_OUT[18]), .A3(
        \unit_decode/n2096 ), .ZN(\unit_decode/n2891 ) );
  NOR3_X1 U4314 ( .A1(\unit_decode/n2093 ), .A2(IR_OUT[24]), .A3(
        \unit_decode/n2091 ), .ZN(\unit_decode/n3497 ) );
  NOR3_X1 U4315 ( .A1(IR_OUT[23]), .A2(IR_OUT[24]), .A3(\unit_decode/n2091 ), 
        .ZN(\unit_decode/n3509 ) );
  NOR3_X1 U4316 ( .A1(\unit_decode/n2092 ), .A2(IR_OUT[23]), .A3(
        \unit_decode/n2091 ), .ZN(\unit_decode/n3511 ) );
  NOR2_X1 U4317 ( .A1(IR_OUT[21]), .A2(IR_OUT[22]), .ZN(\unit_decode/n3491 )
         );
  NOR2_X1 U4318 ( .A1(IR_OUT[16]), .A2(IR_OUT[17]), .ZN(\unit_decode/n2871 )
         );
  NOR2_X1 U4319 ( .A1(\unit_decode/n2100 ), .A2(IR_OUT[17]), .ZN(
        \unit_decode/n2870 ) );
  AOI221_X1 U4320 ( .B1(n147), .B2(\unit_memory/DRAM/n50 ), .C1(n160), .C2(
        \unit_memory/DRAM/n306 ), .A(\unit_memory/DRAM/n588 ), .ZN(
        \unit_memory/DRAM/n587 ) );
  OAI22_X1 U4321 ( .A1(\unit_memory/DRAM/n2672 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2416 ), .B2(n186), .ZN(\unit_memory/DRAM/n588 ) );
  AOI221_X1 U4322 ( .B1(n147), .B2(\unit_memory/DRAM/n18 ), .C1(n160), .C2(
        \unit_memory/DRAM/n274 ), .A(\unit_memory/DRAM/n592 ), .ZN(
        \unit_memory/DRAM/n591 ) );
  OAI22_X1 U4323 ( .A1(\unit_memory/DRAM/n2640 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2384 ), .B2(n186), .ZN(\unit_memory/DRAM/n592 ) );
  AOI221_X1 U4324 ( .B1(n147), .B2(\unit_memory/DRAM/n51 ), .C1(n160), .C2(
        \unit_memory/DRAM/n307 ), .A(\unit_memory/DRAM/n609 ), .ZN(
        \unit_memory/DRAM/n608 ) );
  OAI22_X1 U4325 ( .A1(\unit_memory/DRAM/n2673 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2417 ), .B2(n186), .ZN(\unit_memory/DRAM/n609 ) );
  AOI221_X1 U4326 ( .B1(n147), .B2(\unit_memory/DRAM/n19 ), .C1(n160), .C2(
        \unit_memory/DRAM/n275 ), .A(\unit_memory/DRAM/n613 ), .ZN(
        \unit_memory/DRAM/n612 ) );
  OAI22_X1 U4327 ( .A1(\unit_memory/DRAM/n2641 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2385 ), .B2(n186), .ZN(\unit_memory/DRAM/n613 ) );
  AOI221_X1 U4328 ( .B1(n147), .B2(\unit_memory/DRAM/n52 ), .C1(n160), .C2(
        \unit_memory/DRAM/n308 ), .A(\unit_memory/DRAM/n630 ), .ZN(
        \unit_memory/DRAM/n629 ) );
  OAI22_X1 U4329 ( .A1(\unit_memory/DRAM/n2674 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2418 ), .B2(n186), .ZN(\unit_memory/DRAM/n630 ) );
  AOI221_X1 U4330 ( .B1(n147), .B2(\unit_memory/DRAM/n20 ), .C1(n160), .C2(
        \unit_memory/DRAM/n276 ), .A(\unit_memory/DRAM/n634 ), .ZN(
        \unit_memory/DRAM/n633 ) );
  OAI22_X1 U4331 ( .A1(\unit_memory/DRAM/n2642 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2386 ), .B2(n186), .ZN(\unit_memory/DRAM/n634 ) );
  AOI221_X1 U4332 ( .B1(n148), .B2(\unit_memory/DRAM/n53 ), .C1(n161), .C2(
        \unit_memory/DRAM/n309 ), .A(\unit_memory/DRAM/n651 ), .ZN(
        \unit_memory/DRAM/n650 ) );
  OAI22_X1 U4333 ( .A1(\unit_memory/DRAM/n2675 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2419 ), .B2(n187), .ZN(\unit_memory/DRAM/n651 ) );
  AOI221_X1 U4334 ( .B1(n148), .B2(\unit_memory/DRAM/n21 ), .C1(n161), .C2(
        \unit_memory/DRAM/n277 ), .A(\unit_memory/DRAM/n655 ), .ZN(
        \unit_memory/DRAM/n654 ) );
  OAI22_X1 U4335 ( .A1(\unit_memory/DRAM/n2643 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2387 ), .B2(n187), .ZN(\unit_memory/DRAM/n655 ) );
  AOI221_X1 U4336 ( .B1(n148), .B2(\unit_memory/DRAM/n54 ), .C1(n161), .C2(
        \unit_memory/DRAM/n310 ), .A(\unit_memory/DRAM/n672 ), .ZN(
        \unit_memory/DRAM/n671 ) );
  OAI22_X1 U4337 ( .A1(\unit_memory/DRAM/n2676 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2420 ), .B2(n187), .ZN(\unit_memory/DRAM/n672 ) );
  AOI221_X1 U4338 ( .B1(n148), .B2(\unit_memory/DRAM/n22 ), .C1(n161), .C2(
        \unit_memory/DRAM/n278 ), .A(\unit_memory/DRAM/n676 ), .ZN(
        \unit_memory/DRAM/n675 ) );
  OAI22_X1 U4339 ( .A1(\unit_memory/DRAM/n2644 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2388 ), .B2(n187), .ZN(\unit_memory/DRAM/n676 ) );
  AOI221_X1 U4340 ( .B1(n148), .B2(\unit_memory/DRAM/n55 ), .C1(n161), .C2(
        \unit_memory/DRAM/n311 ), .A(\unit_memory/DRAM/n693 ), .ZN(
        \unit_memory/DRAM/n692 ) );
  OAI22_X1 U4341 ( .A1(\unit_memory/DRAM/n2677 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2421 ), .B2(n187), .ZN(\unit_memory/DRAM/n693 ) );
  AOI221_X1 U4342 ( .B1(n148), .B2(\unit_memory/DRAM/n23 ), .C1(n161), .C2(
        \unit_memory/DRAM/n279 ), .A(\unit_memory/DRAM/n697 ), .ZN(
        \unit_memory/DRAM/n696 ) );
  OAI22_X1 U4343 ( .A1(\unit_memory/DRAM/n2645 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2389 ), .B2(n187), .ZN(\unit_memory/DRAM/n697 ) );
  AOI221_X1 U4344 ( .B1(n149), .B2(\unit_memory/DRAM/n56 ), .C1(n162), .C2(
        \unit_memory/DRAM/n312 ), .A(\unit_memory/DRAM/n714 ), .ZN(
        \unit_memory/DRAM/n713 ) );
  OAI22_X1 U4345 ( .A1(\unit_memory/DRAM/n2678 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2422 ), .B2(n188), .ZN(\unit_memory/DRAM/n714 ) );
  AOI221_X1 U4346 ( .B1(n149), .B2(\unit_memory/DRAM/n24 ), .C1(n162), .C2(
        \unit_memory/DRAM/n280 ), .A(\unit_memory/DRAM/n718 ), .ZN(
        \unit_memory/DRAM/n717 ) );
  OAI22_X1 U4347 ( .A1(\unit_memory/DRAM/n2646 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2390 ), .B2(n188), .ZN(\unit_memory/DRAM/n718 ) );
  AOI221_X1 U4348 ( .B1(n150), .B2(\unit_memory/DRAM/n58 ), .C1(n163), .C2(
        \unit_memory/DRAM/n314 ), .A(\unit_memory/DRAM/n2235 ), .ZN(
        \unit_memory/DRAM/n2234 ) );
  OAI22_X1 U4349 ( .A1(\unit_memory/DRAM/n2680 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2424 ), .B2(n189), .ZN(\unit_memory/DRAM/n2235 ) );
  AOI221_X1 U4350 ( .B1(n151), .B2(\unit_memory/DRAM/n26 ), .C1(n164), .C2(
        \unit_memory/DRAM/n282 ), .A(\unit_memory/DRAM/n2239 ), .ZN(
        \unit_memory/DRAM/n2238 ) );
  OAI22_X1 U4351 ( .A1(\unit_memory/DRAM/n2648 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2392 ), .B2(n190), .ZN(\unit_memory/DRAM/n2239 ) );
  AOI221_X1 U4352 ( .B1(n152), .B2(\unit_memory/DRAM/n59 ), .C1(n165), .C2(
        \unit_memory/DRAM/n315 ), .A(\unit_memory/DRAM/n2256 ), .ZN(
        \unit_memory/DRAM/n2255 ) );
  OAI22_X1 U4353 ( .A1(\unit_memory/DRAM/n2681 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2425 ), .B2(n191), .ZN(\unit_memory/DRAM/n2256 ) );
  AOI221_X1 U4354 ( .B1(n152), .B2(\unit_memory/DRAM/n27 ), .C1(n165), .C2(
        \unit_memory/DRAM/n283 ), .A(\unit_memory/DRAM/n2260 ), .ZN(
        \unit_memory/DRAM/n2259 ) );
  OAI22_X1 U4355 ( .A1(\unit_memory/DRAM/n2649 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2393 ), .B2(n191), .ZN(\unit_memory/DRAM/n2260 ) );
  AOI221_X1 U4356 ( .B1(n152), .B2(\unit_memory/DRAM/n60 ), .C1(n165), .C2(
        \unit_memory/DRAM/n316 ), .A(\unit_memory/DRAM/n2277 ), .ZN(
        \unit_memory/DRAM/n2276 ) );
  OAI22_X1 U4357 ( .A1(\unit_memory/DRAM/n2682 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2426 ), .B2(n191), .ZN(\unit_memory/DRAM/n2277 ) );
  AOI221_X1 U4358 ( .B1(n151), .B2(\unit_memory/DRAM/n28 ), .C1(n164), .C2(
        \unit_memory/DRAM/n284 ), .A(\unit_memory/DRAM/n2281 ), .ZN(
        \unit_memory/DRAM/n2280 ) );
  OAI22_X1 U4359 ( .A1(\unit_memory/DRAM/n2650 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2394 ), .B2(n190), .ZN(\unit_memory/DRAM/n2281 ) );
  AOI221_X1 U4360 ( .B1(n151), .B2(\unit_memory/DRAM/n61 ), .C1(n164), .C2(
        \unit_memory/DRAM/n317 ), .A(\unit_memory/DRAM/n2298 ), .ZN(
        \unit_memory/DRAM/n2297 ) );
  OAI22_X1 U4361 ( .A1(\unit_memory/DRAM/n2683 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2427 ), .B2(n190), .ZN(\unit_memory/DRAM/n2298 ) );
  AOI221_X1 U4362 ( .B1(n152), .B2(\unit_memory/DRAM/n29 ), .C1(n165), .C2(
        \unit_memory/DRAM/n285 ), .A(\unit_memory/DRAM/n2302 ), .ZN(
        \unit_memory/DRAM/n2301 ) );
  OAI22_X1 U4363 ( .A1(\unit_memory/DRAM/n2651 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2395 ), .B2(n191), .ZN(\unit_memory/DRAM/n2302 ) );
  AOI221_X1 U4364 ( .B1(n152), .B2(\unit_memory/DRAM/n62 ), .C1(n165), .C2(
        \unit_memory/DRAM/n318 ), .A(\unit_memory/DRAM/n2319 ), .ZN(
        \unit_memory/DRAM/n2318 ) );
  OAI22_X1 U4365 ( .A1(\unit_memory/DRAM/n2684 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2428 ), .B2(n191), .ZN(\unit_memory/DRAM/n2319 ) );
  AOI221_X1 U4366 ( .B1(n150), .B2(\unit_memory/DRAM/n30 ), .C1(n163), .C2(
        \unit_memory/DRAM/n286 ), .A(\unit_memory/DRAM/n2323 ), .ZN(
        \unit_memory/DRAM/n2322 ) );
  OAI22_X1 U4367 ( .A1(\unit_memory/DRAM/n2652 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2396 ), .B2(n189), .ZN(\unit_memory/DRAM/n2323 ) );
  AOI221_X1 U4368 ( .B1(n152), .B2(\unit_memory/DRAM/n63 ), .C1(n165), .C2(
        \unit_memory/DRAM/n319 ), .A(\unit_memory/DRAM/n2340 ), .ZN(
        \unit_memory/DRAM/n2339 ) );
  OAI22_X1 U4369 ( .A1(\unit_memory/DRAM/n2685 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2429 ), .B2(n191), .ZN(\unit_memory/DRAM/n2340 ) );
  AOI221_X1 U4370 ( .B1(n151), .B2(\unit_memory/DRAM/n31 ), .C1(n164), .C2(
        \unit_memory/DRAM/n287 ), .A(\unit_memory/DRAM/n2344 ), .ZN(
        \unit_memory/DRAM/n2343 ) );
  OAI22_X1 U4371 ( .A1(\unit_memory/DRAM/n2653 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2397 ), .B2(n190), .ZN(\unit_memory/DRAM/n2344 ) );
  AOI221_X1 U4372 ( .B1(n150), .B2(\unit_memory/DRAM/n64 ), .C1(n163), .C2(
        \unit_memory/DRAM/n320 ), .A(\unit_memory/DRAM/n2361 ), .ZN(
        \unit_memory/DRAM/n2360 ) );
  OAI22_X1 U4373 ( .A1(\unit_memory/DRAM/n2686 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2430 ), .B2(n189), .ZN(\unit_memory/DRAM/n2361 ) );
  AOI221_X1 U4374 ( .B1(n147), .B2(\unit_memory/DRAM/n32 ), .C1(n160), .C2(
        \unit_memory/DRAM/n288 ), .A(\unit_memory/DRAM/n2365 ), .ZN(
        \unit_memory/DRAM/n2364 ) );
  OAI22_X1 U4375 ( .A1(\unit_memory/DRAM/n2654 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2398 ), .B2(n186), .ZN(\unit_memory/DRAM/n2365 ) );
  AOI221_X1 U4376 ( .B1(n199), .B2(\unit_memory/DRAM/n178 ), .C1(n212), .C2(
        \unit_memory/DRAM/n434 ), .A(\unit_memory/DRAM/n589 ), .ZN(
        \unit_memory/DRAM/n586 ) );
  OAI22_X1 U4377 ( .A1(\unit_memory/DRAM/n2800 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2544 ), .B2(n238), .ZN(\unit_memory/DRAM/n589 ) );
  AOI221_X1 U4378 ( .B1(n199), .B2(\unit_memory/DRAM/n146 ), .C1(n212), .C2(
        \unit_memory/DRAM/n402 ), .A(\unit_memory/DRAM/n593 ), .ZN(
        \unit_memory/DRAM/n590 ) );
  OAI22_X1 U4379 ( .A1(\unit_memory/DRAM/n2768 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2512 ), .B2(n238), .ZN(\unit_memory/DRAM/n593 ) );
  AOI221_X1 U4380 ( .B1(n199), .B2(\unit_memory/DRAM/n179 ), .C1(n212), .C2(
        \unit_memory/DRAM/n435 ), .A(\unit_memory/DRAM/n610 ), .ZN(
        \unit_memory/DRAM/n607 ) );
  OAI22_X1 U4381 ( .A1(\unit_memory/DRAM/n2801 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2545 ), .B2(n238), .ZN(\unit_memory/DRAM/n610 ) );
  AOI221_X1 U4382 ( .B1(n199), .B2(\unit_memory/DRAM/n147 ), .C1(n212), .C2(
        \unit_memory/DRAM/n403 ), .A(\unit_memory/DRAM/n614 ), .ZN(
        \unit_memory/DRAM/n611 ) );
  OAI22_X1 U4383 ( .A1(\unit_memory/DRAM/n2769 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2513 ), .B2(n238), .ZN(\unit_memory/DRAM/n614 ) );
  AOI221_X1 U4384 ( .B1(n199), .B2(\unit_memory/DRAM/n180 ), .C1(n212), .C2(
        \unit_memory/DRAM/n436 ), .A(\unit_memory/DRAM/n631 ), .ZN(
        \unit_memory/DRAM/n628 ) );
  OAI22_X1 U4385 ( .A1(\unit_memory/DRAM/n2802 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2546 ), .B2(n238), .ZN(\unit_memory/DRAM/n631 ) );
  AOI221_X1 U4386 ( .B1(n199), .B2(\unit_memory/DRAM/n148 ), .C1(n212), .C2(
        \unit_memory/DRAM/n404 ), .A(\unit_memory/DRAM/n635 ), .ZN(
        \unit_memory/DRAM/n632 ) );
  OAI22_X1 U4387 ( .A1(\unit_memory/DRAM/n2770 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2514 ), .B2(n238), .ZN(\unit_memory/DRAM/n635 ) );
  AOI221_X1 U4388 ( .B1(n200), .B2(\unit_memory/DRAM/n181 ), .C1(n213), .C2(
        \unit_memory/DRAM/n437 ), .A(\unit_memory/DRAM/n652 ), .ZN(
        \unit_memory/DRAM/n649 ) );
  OAI22_X1 U4389 ( .A1(\unit_memory/DRAM/n2803 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2547 ), .B2(n239), .ZN(\unit_memory/DRAM/n652 ) );
  AOI221_X1 U4390 ( .B1(n200), .B2(\unit_memory/DRAM/n149 ), .C1(n213), .C2(
        \unit_memory/DRAM/n405 ), .A(\unit_memory/DRAM/n656 ), .ZN(
        \unit_memory/DRAM/n653 ) );
  OAI22_X1 U4391 ( .A1(\unit_memory/DRAM/n2771 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2515 ), .B2(n239), .ZN(\unit_memory/DRAM/n656 ) );
  AOI221_X1 U4392 ( .B1(n200), .B2(\unit_memory/DRAM/n182 ), .C1(n213), .C2(
        \unit_memory/DRAM/n438 ), .A(\unit_memory/DRAM/n673 ), .ZN(
        \unit_memory/DRAM/n670 ) );
  OAI22_X1 U4393 ( .A1(\unit_memory/DRAM/n2804 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2548 ), .B2(n239), .ZN(\unit_memory/DRAM/n673 ) );
  AOI221_X1 U4394 ( .B1(n200), .B2(\unit_memory/DRAM/n150 ), .C1(n213), .C2(
        \unit_memory/DRAM/n406 ), .A(\unit_memory/DRAM/n677 ), .ZN(
        \unit_memory/DRAM/n674 ) );
  OAI22_X1 U4395 ( .A1(\unit_memory/DRAM/n2772 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2516 ), .B2(n239), .ZN(\unit_memory/DRAM/n677 ) );
  AOI221_X1 U4396 ( .B1(n200), .B2(\unit_memory/DRAM/n183 ), .C1(n213), .C2(
        \unit_memory/DRAM/n439 ), .A(\unit_memory/DRAM/n694 ), .ZN(
        \unit_memory/DRAM/n691 ) );
  OAI22_X1 U4397 ( .A1(\unit_memory/DRAM/n2805 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2549 ), .B2(n239), .ZN(\unit_memory/DRAM/n694 ) );
  AOI221_X1 U4398 ( .B1(n200), .B2(\unit_memory/DRAM/n151 ), .C1(n213), .C2(
        \unit_memory/DRAM/n407 ), .A(\unit_memory/DRAM/n698 ), .ZN(
        \unit_memory/DRAM/n695 ) );
  OAI22_X1 U4399 ( .A1(\unit_memory/DRAM/n2773 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2517 ), .B2(n239), .ZN(\unit_memory/DRAM/n698 ) );
  AOI221_X1 U4400 ( .B1(n201), .B2(\unit_memory/DRAM/n184 ), .C1(n214), .C2(
        \unit_memory/DRAM/n440 ), .A(\unit_memory/DRAM/n715 ), .ZN(
        \unit_memory/DRAM/n712 ) );
  OAI22_X1 U4401 ( .A1(\unit_memory/DRAM/n2806 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2550 ), .B2(n240), .ZN(\unit_memory/DRAM/n715 ) );
  AOI221_X1 U4402 ( .B1(n201), .B2(\unit_memory/DRAM/n152 ), .C1(n214), .C2(
        \unit_memory/DRAM/n408 ), .A(\unit_memory/DRAM/n719 ), .ZN(
        \unit_memory/DRAM/n716 ) );
  OAI22_X1 U4403 ( .A1(\unit_memory/DRAM/n2774 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2518 ), .B2(n240), .ZN(\unit_memory/DRAM/n719 ) );
  AOI221_X1 U4404 ( .B1(n202), .B2(\unit_memory/DRAM/n186 ), .C1(n215), .C2(
        \unit_memory/DRAM/n442 ), .A(\unit_memory/DRAM/n2236 ), .ZN(
        \unit_memory/DRAM/n2233 ) );
  OAI22_X1 U4405 ( .A1(\unit_memory/DRAM/n2808 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2552 ), .B2(n241), .ZN(\unit_memory/DRAM/n2236 ) );
  AOI221_X1 U4406 ( .B1(n203), .B2(\unit_memory/DRAM/n154 ), .C1(n216), .C2(
        \unit_memory/DRAM/n410 ), .A(\unit_memory/DRAM/n2240 ), .ZN(
        \unit_memory/DRAM/n2237 ) );
  OAI22_X1 U4407 ( .A1(\unit_memory/DRAM/n2776 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2520 ), .B2(n242), .ZN(\unit_memory/DRAM/n2240 ) );
  AOI221_X1 U4408 ( .B1(n204), .B2(\unit_memory/DRAM/n187 ), .C1(n217), .C2(
        \unit_memory/DRAM/n443 ), .A(\unit_memory/DRAM/n2257 ), .ZN(
        \unit_memory/DRAM/n2254 ) );
  OAI22_X1 U4409 ( .A1(\unit_memory/DRAM/n2809 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2553 ), .B2(n243), .ZN(\unit_memory/DRAM/n2257 ) );
  AOI221_X1 U4410 ( .B1(n204), .B2(\unit_memory/DRAM/n155 ), .C1(n217), .C2(
        \unit_memory/DRAM/n411 ), .A(\unit_memory/DRAM/n2261 ), .ZN(
        \unit_memory/DRAM/n2258 ) );
  OAI22_X1 U4411 ( .A1(\unit_memory/DRAM/n2777 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2521 ), .B2(n243), .ZN(\unit_memory/DRAM/n2261 ) );
  AOI221_X1 U4412 ( .B1(n204), .B2(\unit_memory/DRAM/n188 ), .C1(n217), .C2(
        \unit_memory/DRAM/n444 ), .A(\unit_memory/DRAM/n2278 ), .ZN(
        \unit_memory/DRAM/n2275 ) );
  OAI22_X1 U4413 ( .A1(\unit_memory/DRAM/n2810 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2554 ), .B2(n243), .ZN(\unit_memory/DRAM/n2278 ) );
  AOI221_X1 U4414 ( .B1(n203), .B2(\unit_memory/DRAM/n156 ), .C1(n216), .C2(
        \unit_memory/DRAM/n412 ), .A(\unit_memory/DRAM/n2282 ), .ZN(
        \unit_memory/DRAM/n2279 ) );
  OAI22_X1 U4415 ( .A1(\unit_memory/DRAM/n2778 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2522 ), .B2(n242), .ZN(\unit_memory/DRAM/n2282 ) );
  AOI221_X1 U4416 ( .B1(n203), .B2(\unit_memory/DRAM/n189 ), .C1(n216), .C2(
        \unit_memory/DRAM/n445 ), .A(\unit_memory/DRAM/n2299 ), .ZN(
        \unit_memory/DRAM/n2296 ) );
  OAI22_X1 U4417 ( .A1(\unit_memory/DRAM/n2811 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2555 ), .B2(n242), .ZN(\unit_memory/DRAM/n2299 ) );
  AOI221_X1 U4418 ( .B1(n204), .B2(\unit_memory/DRAM/n157 ), .C1(n217), .C2(
        \unit_memory/DRAM/n413 ), .A(\unit_memory/DRAM/n2303 ), .ZN(
        \unit_memory/DRAM/n2300 ) );
  OAI22_X1 U4419 ( .A1(\unit_memory/DRAM/n2779 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2523 ), .B2(n243), .ZN(\unit_memory/DRAM/n2303 ) );
  AOI221_X1 U4420 ( .B1(n204), .B2(\unit_memory/DRAM/n190 ), .C1(n217), .C2(
        \unit_memory/DRAM/n446 ), .A(\unit_memory/DRAM/n2320 ), .ZN(
        \unit_memory/DRAM/n2317 ) );
  OAI22_X1 U4421 ( .A1(\unit_memory/DRAM/n2812 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2556 ), .B2(n243), .ZN(\unit_memory/DRAM/n2320 ) );
  AOI221_X1 U4422 ( .B1(n202), .B2(\unit_memory/DRAM/n158 ), .C1(n215), .C2(
        \unit_memory/DRAM/n414 ), .A(\unit_memory/DRAM/n2324 ), .ZN(
        \unit_memory/DRAM/n2321 ) );
  OAI22_X1 U4423 ( .A1(\unit_memory/DRAM/n2780 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2524 ), .B2(n241), .ZN(\unit_memory/DRAM/n2324 ) );
  AOI221_X1 U4424 ( .B1(n204), .B2(\unit_memory/DRAM/n191 ), .C1(n217), .C2(
        \unit_memory/DRAM/n447 ), .A(\unit_memory/DRAM/n2341 ), .ZN(
        \unit_memory/DRAM/n2338 ) );
  OAI22_X1 U4425 ( .A1(\unit_memory/DRAM/n2813 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2557 ), .B2(n243), .ZN(\unit_memory/DRAM/n2341 ) );
  AOI221_X1 U4426 ( .B1(n203), .B2(\unit_memory/DRAM/n159 ), .C1(n216), .C2(
        \unit_memory/DRAM/n415 ), .A(\unit_memory/DRAM/n2345 ), .ZN(
        \unit_memory/DRAM/n2342 ) );
  OAI22_X1 U4427 ( .A1(\unit_memory/DRAM/n2781 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2525 ), .B2(n242), .ZN(\unit_memory/DRAM/n2345 ) );
  AOI221_X1 U4428 ( .B1(n202), .B2(\unit_memory/DRAM/n192 ), .C1(n215), .C2(
        \unit_memory/DRAM/n448 ), .A(\unit_memory/DRAM/n2362 ), .ZN(
        \unit_memory/DRAM/n2359 ) );
  OAI22_X1 U4429 ( .A1(\unit_memory/DRAM/n2814 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2558 ), .B2(n241), .ZN(\unit_memory/DRAM/n2362 ) );
  AOI221_X1 U4430 ( .B1(n199), .B2(\unit_memory/DRAM/n160 ), .C1(n212), .C2(
        \unit_memory/DRAM/n416 ), .A(\unit_memory/DRAM/n2366 ), .ZN(
        \unit_memory/DRAM/n2363 ) );
  OAI22_X1 U4431 ( .A1(\unit_memory/DRAM/n2782 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2526 ), .B2(n238), .ZN(\unit_memory/DRAM/n2366 ) );
  OAI221_X1 U4432 ( .B1(\unit_decode/n1907 ), .B2(n1095), .C1(
        \unit_decode/n1899 ), .C2(n1098), .A(\unit_decode/n2436 ), .ZN(
        \unit_decode/n2435 ) );
  AOI22_X1 U4433 ( .A1(n1101), .A2(\unit_decode/n4114 ), .B1(n1102), .B2(
        \unit_decode/n3682 ), .ZN(\unit_decode/n2436 ) );
  OAI221_X1 U4434 ( .B1(\unit_decode/n1939 ), .B2(n1143), .C1(
        \unit_decode/n1931 ), .C2(n1146), .A(\unit_decode/n2444 ), .ZN(
        \unit_decode/n2443 ) );
  AOI22_X1 U4435 ( .A1(n1149), .A2(\unit_decode/n4112 ), .B1(n1150), .B2(
        \unit_decode/n3862 ), .ZN(\unit_decode/n2444 ) );
  OAI221_X1 U4436 ( .B1(\unit_decode/n1906 ), .B2(n1095), .C1(
        \unit_decode/n1898 ), .C2(n1098), .A(\unit_decode/n2418 ), .ZN(
        \unit_decode/n2417 ) );
  AOI22_X1 U4437 ( .A1(n1101), .A2(\unit_decode/n4110 ), .B1(n1102), .B2(
        \unit_decode/n3676 ), .ZN(\unit_decode/n2418 ) );
  OAI221_X1 U4438 ( .B1(\unit_decode/n1938 ), .B2(n1143), .C1(
        \unit_decode/n1930 ), .C2(n1146), .A(\unit_decode/n2426 ), .ZN(
        \unit_decode/n2425 ) );
  AOI22_X1 U4439 ( .A1(n1149), .A2(\unit_decode/n4108 ), .B1(n1150), .B2(
        \unit_decode/n3856 ), .ZN(\unit_decode/n2426 ) );
  OAI221_X1 U4440 ( .B1(\unit_decode/n1905 ), .B2(n1095), .C1(
        \unit_decode/n1897 ), .C2(n1098), .A(\unit_decode/n2400 ), .ZN(
        \unit_decode/n2399 ) );
  AOI22_X1 U4441 ( .A1(n1101), .A2(\unit_decode/n4106 ), .B1(n1102), .B2(
        \unit_decode/n3670 ), .ZN(\unit_decode/n2400 ) );
  OAI221_X1 U4442 ( .B1(\unit_decode/n1937 ), .B2(n1143), .C1(
        \unit_decode/n1929 ), .C2(n1146), .A(\unit_decode/n2408 ), .ZN(
        \unit_decode/n2407 ) );
  AOI22_X1 U4443 ( .A1(n1149), .A2(\unit_decode/n4104 ), .B1(n1150), .B2(
        \unit_decode/n3850 ), .ZN(\unit_decode/n2408 ) );
  OAI221_X1 U4444 ( .B1(\unit_decode/n1904 ), .B2(n1095), .C1(
        \unit_decode/n1896 ), .C2(n1098), .A(\unit_decode/n2382 ), .ZN(
        \unit_decode/n2381 ) );
  AOI22_X1 U4445 ( .A1(n1101), .A2(\unit_decode/n4102 ), .B1(n1102), .B2(
        \unit_decode/n3664 ), .ZN(\unit_decode/n2382 ) );
  OAI221_X1 U4446 ( .B1(\unit_decode/n1936 ), .B2(n1143), .C1(
        \unit_decode/n1928 ), .C2(n1146), .A(\unit_decode/n2390 ), .ZN(
        \unit_decode/n2389 ) );
  AOI22_X1 U4447 ( .A1(n1149), .A2(\unit_decode/n4100 ), .B1(n1150), .B2(
        \unit_decode/n3844 ), .ZN(\unit_decode/n2390 ) );
  OAI221_X1 U4448 ( .B1(\unit_decode/n1903 ), .B2(n1095), .C1(
        \unit_decode/n1895 ), .C2(n1098), .A(\unit_decode/n2364 ), .ZN(
        \unit_decode/n2363 ) );
  AOI22_X1 U4449 ( .A1(n1101), .A2(\unit_decode/n4098 ), .B1(n1102), .B2(
        \unit_decode/n3658 ), .ZN(\unit_decode/n2364 ) );
  OAI221_X1 U4450 ( .B1(\unit_decode/n1935 ), .B2(n1143), .C1(
        \unit_decode/n1927 ), .C2(n1146), .A(\unit_decode/n2372 ), .ZN(
        \unit_decode/n2371 ) );
  AOI22_X1 U4451 ( .A1(n1149), .A2(\unit_decode/n4096 ), .B1(n1150), .B2(
        \unit_decode/n3838 ), .ZN(\unit_decode/n2372 ) );
  OAI221_X1 U4452 ( .B1(\unit_decode/n1902 ), .B2(n1095), .C1(
        \unit_decode/n1894 ), .C2(n1098), .A(\unit_decode/n2346 ), .ZN(
        \unit_decode/n2345 ) );
  AOI22_X1 U4453 ( .A1(n1101), .A2(\unit_decode/n4094 ), .B1(n1102), .B2(
        \unit_decode/n3652 ), .ZN(\unit_decode/n2346 ) );
  OAI221_X1 U4454 ( .B1(\unit_decode/n1934 ), .B2(n1143), .C1(
        \unit_decode/n1926 ), .C2(n1146), .A(\unit_decode/n2354 ), .ZN(
        \unit_decode/n2353 ) );
  AOI22_X1 U4455 ( .A1(n1149), .A2(\unit_decode/n4092 ), .B1(n1150), .B2(
        \unit_decode/n3832 ), .ZN(\unit_decode/n2354 ) );
  OAI221_X1 U4456 ( .B1(\unit_decode/n1901 ), .B2(n1095), .C1(
        \unit_decode/n1893 ), .C2(n1098), .A(\unit_decode/n2328 ), .ZN(
        \unit_decode/n2327 ) );
  AOI22_X1 U4457 ( .A1(n1101), .A2(\unit_decode/n4018 ), .B1(n1102), .B2(
        \unit_decode/n3634 ), .ZN(\unit_decode/n2328 ) );
  OAI221_X1 U4458 ( .B1(\unit_decode/n1933 ), .B2(n1143), .C1(
        \unit_decode/n1925 ), .C2(n1146), .A(\unit_decode/n2336 ), .ZN(
        \unit_decode/n2335 ) );
  AOI22_X1 U4459 ( .A1(n1149), .A2(\unit_decode/n4016 ), .B1(n1150), .B2(
        \unit_decode/n3646 ), .ZN(\unit_decode/n2336 ) );
  OAI221_X1 U4460 ( .B1(\unit_decode/n1900 ), .B2(n1095), .C1(
        \unit_decode/n1892 ), .C2(n1098), .A(\unit_decode/n2280 ), .ZN(
        \unit_decode/n2277 ) );
  AOI22_X1 U4461 ( .A1(n1101), .A2(\unit_decode/n4014 ), .B1(n1102), .B2(
        \unit_decode/n3628 ), .ZN(\unit_decode/n2280 ) );
  OAI221_X1 U4462 ( .B1(\unit_decode/n1932 ), .B2(n1143), .C1(
        \unit_decode/n1924 ), .C2(n1146), .A(\unit_decode/n2304 ), .ZN(
        \unit_decode/n2301 ) );
  AOI22_X1 U4463 ( .A1(n1149), .A2(\unit_decode/n4012 ), .B1(n1150), .B2(
        \unit_decode/n3640 ), .ZN(\unit_decode/n2304 ) );
  OAI221_X1 U4464 ( .B1(\unit_decode/n1907 ), .B2(n1191), .C1(
        \unit_decode/n1899 ), .C2(n1194), .A(\unit_decode/n3056 ), .ZN(
        \unit_decode/n3055 ) );
  AOI22_X1 U4465 ( .A1(n1197), .A2(\unit_decode/n4114 ), .B1(n1198), .B2(
        \unit_decode/n3682 ), .ZN(\unit_decode/n3056 ) );
  OAI221_X1 U4466 ( .B1(\unit_decode/n1939 ), .B2(n1239), .C1(
        \unit_decode/n1931 ), .C2(n1242), .A(\unit_decode/n3064 ), .ZN(
        \unit_decode/n3063 ) );
  AOI22_X1 U4467 ( .A1(n1245), .A2(\unit_decode/n4112 ), .B1(n1246), .B2(
        \unit_decode/n3862 ), .ZN(\unit_decode/n3064 ) );
  OAI221_X1 U4468 ( .B1(\unit_decode/n1906 ), .B2(n1191), .C1(
        \unit_decode/n1898 ), .C2(n1194), .A(\unit_decode/n3038 ), .ZN(
        \unit_decode/n3037 ) );
  AOI22_X1 U4469 ( .A1(n1197), .A2(\unit_decode/n4110 ), .B1(n1198), .B2(
        \unit_decode/n3676 ), .ZN(\unit_decode/n3038 ) );
  OAI221_X1 U4470 ( .B1(\unit_decode/n1938 ), .B2(n1239), .C1(
        \unit_decode/n1930 ), .C2(n1242), .A(\unit_decode/n3046 ), .ZN(
        \unit_decode/n3045 ) );
  AOI22_X1 U4471 ( .A1(n1245), .A2(\unit_decode/n4108 ), .B1(n1246), .B2(
        \unit_decode/n3856 ), .ZN(\unit_decode/n3046 ) );
  OAI221_X1 U4472 ( .B1(\unit_decode/n1905 ), .B2(n1191), .C1(
        \unit_decode/n1897 ), .C2(n1194), .A(\unit_decode/n3020 ), .ZN(
        \unit_decode/n3019 ) );
  AOI22_X1 U4473 ( .A1(n1197), .A2(\unit_decode/n4106 ), .B1(n1198), .B2(
        \unit_decode/n3670 ), .ZN(\unit_decode/n3020 ) );
  OAI221_X1 U4474 ( .B1(\unit_decode/n1937 ), .B2(n1239), .C1(
        \unit_decode/n1929 ), .C2(n1242), .A(\unit_decode/n3028 ), .ZN(
        \unit_decode/n3027 ) );
  AOI22_X1 U4475 ( .A1(n1245), .A2(\unit_decode/n4104 ), .B1(n1246), .B2(
        \unit_decode/n3850 ), .ZN(\unit_decode/n3028 ) );
  OAI221_X1 U4476 ( .B1(\unit_decode/n1904 ), .B2(n1191), .C1(
        \unit_decode/n1896 ), .C2(n1194), .A(\unit_decode/n3002 ), .ZN(
        \unit_decode/n3001 ) );
  AOI22_X1 U4477 ( .A1(n1197), .A2(\unit_decode/n4102 ), .B1(n1198), .B2(
        \unit_decode/n3664 ), .ZN(\unit_decode/n3002 ) );
  OAI221_X1 U4478 ( .B1(\unit_decode/n1936 ), .B2(n1239), .C1(
        \unit_decode/n1928 ), .C2(n1242), .A(\unit_decode/n3010 ), .ZN(
        \unit_decode/n3009 ) );
  AOI22_X1 U4479 ( .A1(n1245), .A2(\unit_decode/n4100 ), .B1(n1246), .B2(
        \unit_decode/n3844 ), .ZN(\unit_decode/n3010 ) );
  OAI221_X1 U4480 ( .B1(\unit_decode/n1903 ), .B2(n1191), .C1(
        \unit_decode/n1895 ), .C2(n1194), .A(\unit_decode/n2984 ), .ZN(
        \unit_decode/n2983 ) );
  AOI22_X1 U4481 ( .A1(n1197), .A2(\unit_decode/n4098 ), .B1(n1198), .B2(
        \unit_decode/n3658 ), .ZN(\unit_decode/n2984 ) );
  OAI221_X1 U4482 ( .B1(\unit_decode/n1935 ), .B2(n1239), .C1(
        \unit_decode/n1927 ), .C2(n1242), .A(\unit_decode/n2992 ), .ZN(
        \unit_decode/n2991 ) );
  AOI22_X1 U4483 ( .A1(n1245), .A2(\unit_decode/n4096 ), .B1(n1246), .B2(
        \unit_decode/n3838 ), .ZN(\unit_decode/n2992 ) );
  OAI221_X1 U4484 ( .B1(\unit_decode/n1902 ), .B2(n1191), .C1(
        \unit_decode/n1894 ), .C2(n1194), .A(\unit_decode/n2966 ), .ZN(
        \unit_decode/n2965 ) );
  AOI22_X1 U4485 ( .A1(n1197), .A2(\unit_decode/n4094 ), .B1(n1198), .B2(
        \unit_decode/n3652 ), .ZN(\unit_decode/n2966 ) );
  OAI221_X1 U4486 ( .B1(\unit_decode/n1934 ), .B2(n1239), .C1(
        \unit_decode/n1926 ), .C2(n1242), .A(\unit_decode/n2974 ), .ZN(
        \unit_decode/n2973 ) );
  AOI22_X1 U4487 ( .A1(n1245), .A2(\unit_decode/n4092 ), .B1(n1246), .B2(
        \unit_decode/n3832 ), .ZN(\unit_decode/n2974 ) );
  OAI221_X1 U4488 ( .B1(\unit_decode/n1901 ), .B2(n1191), .C1(
        \unit_decode/n1893 ), .C2(n1194), .A(\unit_decode/n2948 ), .ZN(
        \unit_decode/n2947 ) );
  AOI22_X1 U4489 ( .A1(n1197), .A2(\unit_decode/n4018 ), .B1(n1198), .B2(
        \unit_decode/n3634 ), .ZN(\unit_decode/n2948 ) );
  OAI221_X1 U4490 ( .B1(\unit_decode/n1933 ), .B2(n1239), .C1(
        \unit_decode/n1925 ), .C2(n1242), .A(\unit_decode/n2956 ), .ZN(
        \unit_decode/n2955 ) );
  AOI22_X1 U4491 ( .A1(n1245), .A2(\unit_decode/n4016 ), .B1(n1246), .B2(
        \unit_decode/n3646 ), .ZN(\unit_decode/n2956 ) );
  OAI221_X1 U4492 ( .B1(\unit_decode/n1900 ), .B2(n1191), .C1(
        \unit_decode/n1892 ), .C2(n1194), .A(\unit_decode/n2900 ), .ZN(
        \unit_decode/n2897 ) );
  AOI22_X1 U4493 ( .A1(n1197), .A2(\unit_decode/n4014 ), .B1(n1198), .B2(
        \unit_decode/n3628 ), .ZN(\unit_decode/n2900 ) );
  OAI221_X1 U4494 ( .B1(\unit_decode/n1932 ), .B2(n1239), .C1(
        \unit_decode/n1924 ), .C2(n1242), .A(\unit_decode/n2924 ), .ZN(
        \unit_decode/n2921 ) );
  AOI22_X1 U4495 ( .A1(n1245), .A2(\unit_decode/n4012 ), .B1(n1246), .B2(
        \unit_decode/n3640 ), .ZN(\unit_decode/n2924 ) );
  OAI221_X1 U4496 ( .B1(\unit_decode/n1580 ), .B2(n1093), .C1(
        \unit_decode/n1556 ), .C2(n1096), .A(\unit_decode/n2868 ), .ZN(
        \unit_decode/n2867 ) );
  AOI22_X1 U4497 ( .A1(n1099), .A2(\unit_decode/n4090 ), .B1(n1104), .B2(
        \unit_decode/n3826 ), .ZN(\unit_decode/n2868 ) );
  OAI221_X1 U4498 ( .B1(\unit_decode/n1676 ), .B2(n1141), .C1(
        \unit_decode/n1652 ), .C2(n1144), .A(\unit_decode/n2884 ), .ZN(
        \unit_decode/n2883 ) );
  AOI22_X1 U4499 ( .A1(n1147), .A2(\unit_decode/n4088 ), .B1(n1152), .B2(
        \unit_decode/n4006 ), .ZN(\unit_decode/n2884 ) );
  OAI221_X1 U4500 ( .B1(\unit_decode/n1581 ), .B2(n1093), .C1(
        \unit_decode/n1557 ), .C2(n1096), .A(\unit_decode/n2850 ), .ZN(
        \unit_decode/n2849 ) );
  AOI22_X1 U4501 ( .A1(n1099), .A2(\unit_decode/n4086 ), .B1(n1104), .B2(
        \unit_decode/n3820 ), .ZN(\unit_decode/n2850 ) );
  OAI221_X1 U4502 ( .B1(\unit_decode/n1677 ), .B2(n1141), .C1(
        \unit_decode/n1653 ), .C2(n1144), .A(\unit_decode/n2858 ), .ZN(
        \unit_decode/n2857 ) );
  AOI22_X1 U4503 ( .A1(n1147), .A2(\unit_decode/n4084 ), .B1(n1152), .B2(
        \unit_decode/n4000 ), .ZN(\unit_decode/n2858 ) );
  OAI221_X1 U4504 ( .B1(\unit_decode/n1582 ), .B2(n1093), .C1(
        \unit_decode/n1558 ), .C2(n1096), .A(\unit_decode/n2832 ), .ZN(
        \unit_decode/n2831 ) );
  AOI22_X1 U4505 ( .A1(n1099), .A2(\unit_decode/n4082 ), .B1(n1104), .B2(
        \unit_decode/n3814 ), .ZN(\unit_decode/n2832 ) );
  OAI221_X1 U4506 ( .B1(\unit_decode/n1678 ), .B2(n1141), .C1(
        \unit_decode/n1654 ), .C2(n1144), .A(\unit_decode/n2840 ), .ZN(
        \unit_decode/n2839 ) );
  AOI22_X1 U4507 ( .A1(n1147), .A2(\unit_decode/n4080 ), .B1(n1152), .B2(
        \unit_decode/n3994 ), .ZN(\unit_decode/n2840 ) );
  OAI221_X1 U4508 ( .B1(\unit_decode/n1583 ), .B2(n1093), .C1(
        \unit_decode/n1559 ), .C2(n1096), .A(\unit_decode/n2814 ), .ZN(
        \unit_decode/n2813 ) );
  AOI22_X1 U4509 ( .A1(n1099), .A2(\unit_decode/n4078 ), .B1(n1104), .B2(
        \unit_decode/n3808 ), .ZN(\unit_decode/n2814 ) );
  OAI221_X1 U4510 ( .B1(\unit_decode/n1679 ), .B2(n1141), .C1(
        \unit_decode/n1655 ), .C2(n1144), .A(\unit_decode/n2822 ), .ZN(
        \unit_decode/n2821 ) );
  AOI22_X1 U4511 ( .A1(n1147), .A2(\unit_decode/n4076 ), .B1(n1152), .B2(
        \unit_decode/n3988 ), .ZN(\unit_decode/n2822 ) );
  OAI221_X1 U4512 ( .B1(\unit_decode/n1584 ), .B2(n1093), .C1(
        \unit_decode/n1560 ), .C2(n1096), .A(\unit_decode/n2796 ), .ZN(
        \unit_decode/n2795 ) );
  AOI22_X1 U4513 ( .A1(n1099), .A2(\unit_decode/n4074 ), .B1(n1104), .B2(
        \unit_decode/n3802 ), .ZN(\unit_decode/n2796 ) );
  OAI221_X1 U4514 ( .B1(\unit_decode/n1680 ), .B2(n1141), .C1(
        \unit_decode/n1656 ), .C2(n1144), .A(\unit_decode/n2804 ), .ZN(
        \unit_decode/n2803 ) );
  AOI22_X1 U4515 ( .A1(n1147), .A2(\unit_decode/n4072 ), .B1(n1152), .B2(
        \unit_decode/n3982 ), .ZN(\unit_decode/n2804 ) );
  OAI221_X1 U4516 ( .B1(\unit_decode/n1585 ), .B2(n1093), .C1(
        \unit_decode/n1561 ), .C2(n1096), .A(\unit_decode/n2778 ), .ZN(
        \unit_decode/n2777 ) );
  AOI22_X1 U4517 ( .A1(n1099), .A2(\unit_decode/n4070 ), .B1(n1104), .B2(
        \unit_decode/n3796 ), .ZN(\unit_decode/n2778 ) );
  OAI221_X1 U4518 ( .B1(\unit_decode/n1681 ), .B2(n1141), .C1(
        \unit_decode/n1657 ), .C2(n1144), .A(\unit_decode/n2786 ), .ZN(
        \unit_decode/n2785 ) );
  AOI22_X1 U4519 ( .A1(n1147), .A2(\unit_decode/n4068 ), .B1(n1152), .B2(
        \unit_decode/n3976 ), .ZN(\unit_decode/n2786 ) );
  OAI221_X1 U4520 ( .B1(\unit_decode/n1586 ), .B2(n1093), .C1(
        \unit_decode/n1562 ), .C2(n1096), .A(\unit_decode/n2760 ), .ZN(
        \unit_decode/n2759 ) );
  AOI22_X1 U4521 ( .A1(n1099), .A2(\unit_decode/n4066 ), .B1(n1104), .B2(
        \unit_decode/n3790 ), .ZN(\unit_decode/n2760 ) );
  OAI221_X1 U4522 ( .B1(\unit_decode/n1682 ), .B2(n1141), .C1(
        \unit_decode/n1658 ), .C2(n1144), .A(\unit_decode/n2768 ), .ZN(
        \unit_decode/n2767 ) );
  AOI22_X1 U4523 ( .A1(n1147), .A2(\unit_decode/n4064 ), .B1(n1152), .B2(
        \unit_decode/n3970 ), .ZN(\unit_decode/n2768 ) );
  OAI221_X1 U4524 ( .B1(\unit_decode/n1587 ), .B2(n1093), .C1(
        \unit_decode/n1563 ), .C2(n1096), .A(\unit_decode/n2742 ), .ZN(
        \unit_decode/n2741 ) );
  AOI22_X1 U4525 ( .A1(n1099), .A2(\unit_decode/n4062 ), .B1(n1104), .B2(
        \unit_decode/n3784 ), .ZN(\unit_decode/n2742 ) );
  OAI221_X1 U4526 ( .B1(\unit_decode/n1683 ), .B2(n1141), .C1(
        \unit_decode/n1659 ), .C2(n1144), .A(\unit_decode/n2750 ), .ZN(
        \unit_decode/n2749 ) );
  AOI22_X1 U4527 ( .A1(n1147), .A2(\unit_decode/n4060 ), .B1(n1152), .B2(
        \unit_decode/n3964 ), .ZN(\unit_decode/n2750 ) );
  OAI221_X1 U4528 ( .B1(\unit_decode/n1588 ), .B2(n1093), .C1(
        \unit_decode/n1564 ), .C2(n1096), .A(\unit_decode/n2724 ), .ZN(
        \unit_decode/n2723 ) );
  AOI22_X1 U4529 ( .A1(n1099), .A2(\unit_decode/n4058 ), .B1(n1103), .B2(
        \unit_decode/n3778 ), .ZN(\unit_decode/n2724 ) );
  OAI221_X1 U4530 ( .B1(\unit_decode/n1684 ), .B2(n1141), .C1(
        \unit_decode/n1660 ), .C2(n1144), .A(\unit_decode/n2732 ), .ZN(
        \unit_decode/n2731 ) );
  AOI22_X1 U4531 ( .A1(n1147), .A2(\unit_decode/n4056 ), .B1(n1151), .B2(
        \unit_decode/n3958 ), .ZN(\unit_decode/n2732 ) );
  OAI221_X1 U4532 ( .B1(\unit_decode/n1589 ), .B2(n1093), .C1(
        \unit_decode/n1565 ), .C2(n1096), .A(\unit_decode/n2706 ), .ZN(
        \unit_decode/n2705 ) );
  AOI22_X1 U4533 ( .A1(n1099), .A2(\unit_decode/n4054 ), .B1(n1103), .B2(
        \unit_decode/n3772 ), .ZN(\unit_decode/n2706 ) );
  OAI221_X1 U4534 ( .B1(\unit_decode/n1685 ), .B2(n1141), .C1(
        \unit_decode/n1661 ), .C2(n1144), .A(\unit_decode/n2714 ), .ZN(
        \unit_decode/n2713 ) );
  AOI22_X1 U4535 ( .A1(n1147), .A2(\unit_decode/n4052 ), .B1(n1151), .B2(
        \unit_decode/n3952 ), .ZN(\unit_decode/n2714 ) );
  OAI221_X1 U4536 ( .B1(\unit_decode/n1590 ), .B2(n1093), .C1(
        \unit_decode/n1566 ), .C2(n1096), .A(\unit_decode/n2688 ), .ZN(
        \unit_decode/n2687 ) );
  AOI22_X1 U4537 ( .A1(n1099), .A2(\unit_decode/n4050 ), .B1(n1103), .B2(
        \unit_decode/n3766 ), .ZN(\unit_decode/n2688 ) );
  OAI221_X1 U4538 ( .B1(\unit_decode/n1686 ), .B2(n1141), .C1(
        \unit_decode/n1662 ), .C2(n1144), .A(\unit_decode/n2696 ), .ZN(
        \unit_decode/n2695 ) );
  AOI22_X1 U4539 ( .A1(n1147), .A2(\unit_decode/n4048 ), .B1(n1151), .B2(
        \unit_decode/n3946 ), .ZN(\unit_decode/n2696 ) );
  OAI221_X1 U4540 ( .B1(\unit_decode/n1591 ), .B2(n1093), .C1(
        \unit_decode/n1567 ), .C2(n1096), .A(\unit_decode/n2670 ), .ZN(
        \unit_decode/n2669 ) );
  AOI22_X1 U4541 ( .A1(n1099), .A2(\unit_decode/n4046 ), .B1(n1103), .B2(
        \unit_decode/n3760 ), .ZN(\unit_decode/n2670 ) );
  OAI221_X1 U4542 ( .B1(\unit_decode/n1687 ), .B2(n1141), .C1(
        \unit_decode/n1663 ), .C2(n1144), .A(\unit_decode/n2678 ), .ZN(
        \unit_decode/n2677 ) );
  AOI22_X1 U4543 ( .A1(n1147), .A2(\unit_decode/n4044 ), .B1(n1151), .B2(
        \unit_decode/n3940 ), .ZN(\unit_decode/n2678 ) );
  OAI221_X1 U4544 ( .B1(\unit_decode/n1592 ), .B2(n1094), .C1(
        \unit_decode/n1568 ), .C2(n1097), .A(\unit_decode/n2652 ), .ZN(
        \unit_decode/n2651 ) );
  AOI22_X1 U4545 ( .A1(n1100), .A2(\unit_decode/n4042 ), .B1(n1103), .B2(
        \unit_decode/n3754 ), .ZN(\unit_decode/n2652 ) );
  OAI221_X1 U4546 ( .B1(\unit_decode/n1688 ), .B2(n1142), .C1(
        \unit_decode/n1664 ), .C2(n1145), .A(\unit_decode/n2660 ), .ZN(
        \unit_decode/n2659 ) );
  AOI22_X1 U4547 ( .A1(n1148), .A2(\unit_decode/n4040 ), .B1(n1151), .B2(
        \unit_decode/n3934 ), .ZN(\unit_decode/n2660 ) );
  OAI221_X1 U4548 ( .B1(\unit_decode/n1593 ), .B2(n1094), .C1(
        \unit_decode/n1569 ), .C2(n1097), .A(\unit_decode/n2634 ), .ZN(
        \unit_decode/n2633 ) );
  AOI22_X1 U4549 ( .A1(n1100), .A2(\unit_decode/n4038 ), .B1(n1103), .B2(
        \unit_decode/n3748 ), .ZN(\unit_decode/n2634 ) );
  OAI221_X1 U4550 ( .B1(\unit_decode/n1689 ), .B2(n1142), .C1(
        \unit_decode/n1665 ), .C2(n1145), .A(\unit_decode/n2642 ), .ZN(
        \unit_decode/n2641 ) );
  AOI22_X1 U4551 ( .A1(n1148), .A2(\unit_decode/n4036 ), .B1(n1151), .B2(
        \unit_decode/n3928 ), .ZN(\unit_decode/n2642 ) );
  OAI221_X1 U4552 ( .B1(\unit_decode/n1594 ), .B2(n1094), .C1(
        \unit_decode/n1570 ), .C2(n1097), .A(\unit_decode/n2616 ), .ZN(
        \unit_decode/n2615 ) );
  AOI22_X1 U4553 ( .A1(n1100), .A2(\unit_decode/n4034 ), .B1(n1103), .B2(
        \unit_decode/n3742 ), .ZN(\unit_decode/n2616 ) );
  OAI221_X1 U4554 ( .B1(\unit_decode/n1690 ), .B2(n1142), .C1(
        \unit_decode/n1666 ), .C2(n1145), .A(\unit_decode/n2624 ), .ZN(
        \unit_decode/n2623 ) );
  AOI22_X1 U4555 ( .A1(n1148), .A2(\unit_decode/n4032 ), .B1(n1151), .B2(
        \unit_decode/n3922 ), .ZN(\unit_decode/n2624 ) );
  OAI221_X1 U4556 ( .B1(\unit_decode/n1595 ), .B2(n1094), .C1(
        \unit_decode/n1571 ), .C2(n1097), .A(\unit_decode/n2598 ), .ZN(
        \unit_decode/n2597 ) );
  AOI22_X1 U4557 ( .A1(n1100), .A2(\unit_decode/n4030 ), .B1(n1103), .B2(
        \unit_decode/n3736 ), .ZN(\unit_decode/n2598 ) );
  OAI221_X1 U4558 ( .B1(\unit_decode/n1691 ), .B2(n1142), .C1(
        \unit_decode/n1667 ), .C2(n1145), .A(\unit_decode/n2606 ), .ZN(
        \unit_decode/n2605 ) );
  AOI22_X1 U4559 ( .A1(n1148), .A2(\unit_decode/n4028 ), .B1(n1151), .B2(
        \unit_decode/n3916 ), .ZN(\unit_decode/n2606 ) );
  OAI221_X1 U4560 ( .B1(\unit_decode/n1596 ), .B2(n1094), .C1(
        \unit_decode/n1572 ), .C2(n1097), .A(\unit_decode/n2580 ), .ZN(
        \unit_decode/n2579 ) );
  AOI22_X1 U4561 ( .A1(n1100), .A2(\unit_decode/n4026 ), .B1(n1103), .B2(
        \unit_decode/n3730 ), .ZN(\unit_decode/n2580 ) );
  OAI221_X1 U4562 ( .B1(\unit_decode/n1692 ), .B2(n1142), .C1(
        \unit_decode/n1668 ), .C2(n1145), .A(\unit_decode/n2588 ), .ZN(
        \unit_decode/n2587 ) );
  AOI22_X1 U4563 ( .A1(n1148), .A2(\unit_decode/n4024 ), .B1(n1151), .B2(
        \unit_decode/n3910 ), .ZN(\unit_decode/n2588 ) );
  OAI221_X1 U4564 ( .B1(\unit_decode/n1597 ), .B2(n1094), .C1(
        \unit_decode/n1573 ), .C2(n1097), .A(\unit_decode/n2562 ), .ZN(
        \unit_decode/n2561 ) );
  AOI22_X1 U4565 ( .A1(n1100), .A2(\unit_decode/n4022 ), .B1(n1103), .B2(
        \unit_decode/n3724 ), .ZN(\unit_decode/n2562 ) );
  OAI221_X1 U4566 ( .B1(\unit_decode/n1693 ), .B2(n1142), .C1(
        \unit_decode/n1669 ), .C2(n1145), .A(\unit_decode/n2570 ), .ZN(
        \unit_decode/n2569 ) );
  AOI22_X1 U4567 ( .A1(n1148), .A2(\unit_decode/n4020 ), .B1(n1151), .B2(
        \unit_decode/n3904 ), .ZN(\unit_decode/n2570 ) );
  OAI221_X1 U4568 ( .B1(\unit_decode/n1598 ), .B2(n1094), .C1(
        \unit_decode/n1574 ), .C2(n1097), .A(\unit_decode/n2544 ), .ZN(
        \unit_decode/n2543 ) );
  AOI22_X1 U4569 ( .A1(n1100), .A2(\unit_decode/n4138 ), .B1(n1103), .B2(
        \unit_decode/n3718 ), .ZN(\unit_decode/n2544 ) );
  OAI221_X1 U4570 ( .B1(\unit_decode/n1694 ), .B2(n1142), .C1(
        \unit_decode/n1670 ), .C2(n1145), .A(\unit_decode/n2552 ), .ZN(
        \unit_decode/n2551 ) );
  AOI22_X1 U4571 ( .A1(n1148), .A2(\unit_decode/n4136 ), .B1(n1151), .B2(
        \unit_decode/n3898 ), .ZN(\unit_decode/n2552 ) );
  OAI221_X1 U4572 ( .B1(\unit_decode/n1599 ), .B2(n1094), .C1(
        \unit_decode/n1575 ), .C2(n1097), .A(\unit_decode/n2526 ), .ZN(
        \unit_decode/n2525 ) );
  AOI22_X1 U4573 ( .A1(n1100), .A2(\unit_decode/n4134 ), .B1(n1103), .B2(
        \unit_decode/n3712 ), .ZN(\unit_decode/n2526 ) );
  OAI221_X1 U4574 ( .B1(\unit_decode/n1695 ), .B2(n1142), .C1(
        \unit_decode/n1671 ), .C2(n1145), .A(\unit_decode/n2534 ), .ZN(
        \unit_decode/n2533 ) );
  AOI22_X1 U4575 ( .A1(n1148), .A2(\unit_decode/n4132 ), .B1(n1151), .B2(
        \unit_decode/n3892 ), .ZN(\unit_decode/n2534 ) );
  OAI221_X1 U4576 ( .B1(\unit_decode/n1600 ), .B2(n1094), .C1(
        \unit_decode/n1576 ), .C2(n1097), .A(\unit_decode/n2508 ), .ZN(
        \unit_decode/n2507 ) );
  AOI22_X1 U4577 ( .A1(n1100), .A2(\unit_decode/n4130 ), .B1(n1102), .B2(
        \unit_decode/n3706 ), .ZN(\unit_decode/n2508 ) );
  OAI221_X1 U4578 ( .B1(\unit_decode/n1696 ), .B2(n1142), .C1(
        \unit_decode/n1672 ), .C2(n1145), .A(\unit_decode/n2516 ), .ZN(
        \unit_decode/n2515 ) );
  AOI22_X1 U4579 ( .A1(n1148), .A2(\unit_decode/n4128 ), .B1(n1150), .B2(
        \unit_decode/n3886 ), .ZN(\unit_decode/n2516 ) );
  OAI221_X1 U4580 ( .B1(\unit_decode/n1601 ), .B2(n1094), .C1(
        \unit_decode/n1577 ), .C2(n1097), .A(\unit_decode/n2490 ), .ZN(
        \unit_decode/n2489 ) );
  AOI22_X1 U4581 ( .A1(n1100), .A2(\unit_decode/n4126 ), .B1(n1102), .B2(
        \unit_decode/n3700 ), .ZN(\unit_decode/n2490 ) );
  OAI221_X1 U4582 ( .B1(\unit_decode/n1697 ), .B2(n1142), .C1(
        \unit_decode/n1673 ), .C2(n1145), .A(\unit_decode/n2498 ), .ZN(
        \unit_decode/n2497 ) );
  AOI22_X1 U4583 ( .A1(n1148), .A2(\unit_decode/n4124 ), .B1(n1150), .B2(
        \unit_decode/n3880 ), .ZN(\unit_decode/n2498 ) );
  OAI221_X1 U4584 ( .B1(\unit_decode/n1602 ), .B2(n1094), .C1(
        \unit_decode/n1578 ), .C2(n1097), .A(\unit_decode/n2472 ), .ZN(
        \unit_decode/n2471 ) );
  AOI22_X1 U4585 ( .A1(n1100), .A2(\unit_decode/n4122 ), .B1(n1102), .B2(
        \unit_decode/n3694 ), .ZN(\unit_decode/n2472 ) );
  OAI221_X1 U4586 ( .B1(\unit_decode/n1698 ), .B2(n1142), .C1(
        \unit_decode/n1674 ), .C2(n1145), .A(\unit_decode/n2480 ), .ZN(
        \unit_decode/n2479 ) );
  AOI22_X1 U4587 ( .A1(n1148), .A2(\unit_decode/n4120 ), .B1(n1150), .B2(
        \unit_decode/n3874 ), .ZN(\unit_decode/n2480 ) );
  OAI221_X1 U4588 ( .B1(\unit_decode/n1603 ), .B2(n1094), .C1(
        \unit_decode/n1579 ), .C2(n1097), .A(\unit_decode/n2454 ), .ZN(
        \unit_decode/n2453 ) );
  AOI22_X1 U4589 ( .A1(n1100), .A2(\unit_decode/n4118 ), .B1(n1102), .B2(
        \unit_decode/n3688 ), .ZN(\unit_decode/n2454 ) );
  OAI221_X1 U4590 ( .B1(\unit_decode/n1699 ), .B2(n1142), .C1(
        \unit_decode/n1675 ), .C2(n1145), .A(\unit_decode/n2462 ), .ZN(
        \unit_decode/n2461 ) );
  AOI22_X1 U4591 ( .A1(n1148), .A2(\unit_decode/n4116 ), .B1(n1150), .B2(
        \unit_decode/n3868 ), .ZN(\unit_decode/n2462 ) );
  OAI221_X1 U4592 ( .B1(\unit_decode/n1580 ), .B2(n1189), .C1(
        \unit_decode/n1556 ), .C2(n1192), .A(\unit_decode/n3488 ), .ZN(
        \unit_decode/n3487 ) );
  AOI22_X1 U4593 ( .A1(n1195), .A2(\unit_decode/n4090 ), .B1(n1200), .B2(
        \unit_decode/n3826 ), .ZN(\unit_decode/n3488 ) );
  OAI221_X1 U4594 ( .B1(\unit_decode/n1676 ), .B2(n1237), .C1(
        \unit_decode/n1652 ), .C2(n1240), .A(\unit_decode/n3504 ), .ZN(
        \unit_decode/n3503 ) );
  AOI22_X1 U4595 ( .A1(n1243), .A2(\unit_decode/n4088 ), .B1(n1248), .B2(
        \unit_decode/n4006 ), .ZN(\unit_decode/n3504 ) );
  OAI221_X1 U4596 ( .B1(\unit_decode/n1581 ), .B2(n1189), .C1(
        \unit_decode/n1557 ), .C2(n1192), .A(\unit_decode/n3470 ), .ZN(
        \unit_decode/n3469 ) );
  AOI22_X1 U4597 ( .A1(n1195), .A2(\unit_decode/n4086 ), .B1(n1200), .B2(
        \unit_decode/n3820 ), .ZN(\unit_decode/n3470 ) );
  OAI221_X1 U4598 ( .B1(\unit_decode/n1677 ), .B2(n1237), .C1(
        \unit_decode/n1653 ), .C2(n1240), .A(\unit_decode/n3478 ), .ZN(
        \unit_decode/n3477 ) );
  AOI22_X1 U4599 ( .A1(n1243), .A2(\unit_decode/n4084 ), .B1(n1248), .B2(
        \unit_decode/n4000 ), .ZN(\unit_decode/n3478 ) );
  OAI221_X1 U4600 ( .B1(\unit_decode/n1582 ), .B2(n1189), .C1(
        \unit_decode/n1558 ), .C2(n1192), .A(\unit_decode/n3452 ), .ZN(
        \unit_decode/n3451 ) );
  AOI22_X1 U4601 ( .A1(n1195), .A2(\unit_decode/n4082 ), .B1(n1200), .B2(
        \unit_decode/n3814 ), .ZN(\unit_decode/n3452 ) );
  OAI221_X1 U4602 ( .B1(\unit_decode/n1678 ), .B2(n1237), .C1(
        \unit_decode/n1654 ), .C2(n1240), .A(\unit_decode/n3460 ), .ZN(
        \unit_decode/n3459 ) );
  AOI22_X1 U4603 ( .A1(n1243), .A2(\unit_decode/n4080 ), .B1(n1248), .B2(
        \unit_decode/n3994 ), .ZN(\unit_decode/n3460 ) );
  OAI221_X1 U4604 ( .B1(\unit_decode/n1583 ), .B2(n1189), .C1(
        \unit_decode/n1559 ), .C2(n1192), .A(\unit_decode/n3434 ), .ZN(
        \unit_decode/n3433 ) );
  AOI22_X1 U4605 ( .A1(n1195), .A2(\unit_decode/n4078 ), .B1(n1200), .B2(
        \unit_decode/n3808 ), .ZN(\unit_decode/n3434 ) );
  OAI221_X1 U4606 ( .B1(\unit_decode/n1679 ), .B2(n1237), .C1(
        \unit_decode/n1655 ), .C2(n1240), .A(\unit_decode/n3442 ), .ZN(
        \unit_decode/n3441 ) );
  AOI22_X1 U4607 ( .A1(n1243), .A2(\unit_decode/n4076 ), .B1(n1248), .B2(
        \unit_decode/n3988 ), .ZN(\unit_decode/n3442 ) );
  OAI221_X1 U4608 ( .B1(\unit_decode/n1584 ), .B2(n1189), .C1(
        \unit_decode/n1560 ), .C2(n1192), .A(\unit_decode/n3416 ), .ZN(
        \unit_decode/n3415 ) );
  AOI22_X1 U4609 ( .A1(n1195), .A2(\unit_decode/n4074 ), .B1(n1200), .B2(
        \unit_decode/n3802 ), .ZN(\unit_decode/n3416 ) );
  OAI221_X1 U4610 ( .B1(\unit_decode/n1680 ), .B2(n1237), .C1(
        \unit_decode/n1656 ), .C2(n1240), .A(\unit_decode/n3424 ), .ZN(
        \unit_decode/n3423 ) );
  AOI22_X1 U4611 ( .A1(n1243), .A2(\unit_decode/n4072 ), .B1(n1248), .B2(
        \unit_decode/n3982 ), .ZN(\unit_decode/n3424 ) );
  OAI221_X1 U4612 ( .B1(\unit_decode/n1585 ), .B2(n1189), .C1(
        \unit_decode/n1561 ), .C2(n1192), .A(\unit_decode/n3398 ), .ZN(
        \unit_decode/n3397 ) );
  AOI22_X1 U4613 ( .A1(n1195), .A2(\unit_decode/n4070 ), .B1(n1200), .B2(
        \unit_decode/n3796 ), .ZN(\unit_decode/n3398 ) );
  OAI221_X1 U4614 ( .B1(\unit_decode/n1681 ), .B2(n1237), .C1(
        \unit_decode/n1657 ), .C2(n1240), .A(\unit_decode/n3406 ), .ZN(
        \unit_decode/n3405 ) );
  AOI22_X1 U4615 ( .A1(n1243), .A2(\unit_decode/n4068 ), .B1(n1248), .B2(
        \unit_decode/n3976 ), .ZN(\unit_decode/n3406 ) );
  OAI221_X1 U4616 ( .B1(\unit_decode/n1586 ), .B2(n1189), .C1(
        \unit_decode/n1562 ), .C2(n1192), .A(\unit_decode/n3380 ), .ZN(
        \unit_decode/n3379 ) );
  AOI22_X1 U4617 ( .A1(n1195), .A2(\unit_decode/n4066 ), .B1(n1200), .B2(
        \unit_decode/n3790 ), .ZN(\unit_decode/n3380 ) );
  OAI221_X1 U4618 ( .B1(\unit_decode/n1682 ), .B2(n1237), .C1(
        \unit_decode/n1658 ), .C2(n1240), .A(\unit_decode/n3388 ), .ZN(
        \unit_decode/n3387 ) );
  AOI22_X1 U4619 ( .A1(n1243), .A2(\unit_decode/n4064 ), .B1(n1248), .B2(
        \unit_decode/n3970 ), .ZN(\unit_decode/n3388 ) );
  OAI221_X1 U4620 ( .B1(\unit_decode/n1587 ), .B2(n1189), .C1(
        \unit_decode/n1563 ), .C2(n1192), .A(\unit_decode/n3362 ), .ZN(
        \unit_decode/n3361 ) );
  AOI22_X1 U4621 ( .A1(n1195), .A2(\unit_decode/n4062 ), .B1(n1200), .B2(
        \unit_decode/n3784 ), .ZN(\unit_decode/n3362 ) );
  OAI221_X1 U4622 ( .B1(\unit_decode/n1683 ), .B2(n1237), .C1(
        \unit_decode/n1659 ), .C2(n1240), .A(\unit_decode/n3370 ), .ZN(
        \unit_decode/n3369 ) );
  AOI22_X1 U4623 ( .A1(n1243), .A2(\unit_decode/n4060 ), .B1(n1248), .B2(
        \unit_decode/n3964 ), .ZN(\unit_decode/n3370 ) );
  OAI221_X1 U4624 ( .B1(\unit_decode/n1588 ), .B2(n1189), .C1(
        \unit_decode/n1564 ), .C2(n1192), .A(\unit_decode/n3344 ), .ZN(
        \unit_decode/n3343 ) );
  AOI22_X1 U4625 ( .A1(n1195), .A2(\unit_decode/n4058 ), .B1(n1199), .B2(
        \unit_decode/n3778 ), .ZN(\unit_decode/n3344 ) );
  OAI221_X1 U4626 ( .B1(\unit_decode/n1684 ), .B2(n1237), .C1(
        \unit_decode/n1660 ), .C2(n1240), .A(\unit_decode/n3352 ), .ZN(
        \unit_decode/n3351 ) );
  AOI22_X1 U4627 ( .A1(n1243), .A2(\unit_decode/n4056 ), .B1(n1247), .B2(
        \unit_decode/n3958 ), .ZN(\unit_decode/n3352 ) );
  OAI221_X1 U4628 ( .B1(\unit_decode/n1589 ), .B2(n1189), .C1(
        \unit_decode/n1565 ), .C2(n1192), .A(\unit_decode/n3326 ), .ZN(
        \unit_decode/n3325 ) );
  AOI22_X1 U4629 ( .A1(n1195), .A2(\unit_decode/n4054 ), .B1(n1199), .B2(
        \unit_decode/n3772 ), .ZN(\unit_decode/n3326 ) );
  OAI221_X1 U4630 ( .B1(\unit_decode/n1685 ), .B2(n1237), .C1(
        \unit_decode/n1661 ), .C2(n1240), .A(\unit_decode/n3334 ), .ZN(
        \unit_decode/n3333 ) );
  AOI22_X1 U4631 ( .A1(n1243), .A2(\unit_decode/n4052 ), .B1(n1247), .B2(
        \unit_decode/n3952 ), .ZN(\unit_decode/n3334 ) );
  OAI221_X1 U4632 ( .B1(\unit_decode/n1590 ), .B2(n1189), .C1(
        \unit_decode/n1566 ), .C2(n1192), .A(\unit_decode/n3308 ), .ZN(
        \unit_decode/n3307 ) );
  AOI22_X1 U4633 ( .A1(n1195), .A2(\unit_decode/n4050 ), .B1(n1199), .B2(
        \unit_decode/n3766 ), .ZN(\unit_decode/n3308 ) );
  OAI221_X1 U4634 ( .B1(\unit_decode/n1686 ), .B2(n1237), .C1(
        \unit_decode/n1662 ), .C2(n1240), .A(\unit_decode/n3316 ), .ZN(
        \unit_decode/n3315 ) );
  AOI22_X1 U4635 ( .A1(n1243), .A2(\unit_decode/n4048 ), .B1(n1247), .B2(
        \unit_decode/n3946 ), .ZN(\unit_decode/n3316 ) );
  OAI221_X1 U4636 ( .B1(\unit_decode/n1591 ), .B2(n1189), .C1(
        \unit_decode/n1567 ), .C2(n1192), .A(\unit_decode/n3290 ), .ZN(
        \unit_decode/n3289 ) );
  AOI22_X1 U4637 ( .A1(n1195), .A2(\unit_decode/n4046 ), .B1(n1199), .B2(
        \unit_decode/n3760 ), .ZN(\unit_decode/n3290 ) );
  OAI221_X1 U4638 ( .B1(\unit_decode/n1687 ), .B2(n1237), .C1(
        \unit_decode/n1663 ), .C2(n1240), .A(\unit_decode/n3298 ), .ZN(
        \unit_decode/n3297 ) );
  AOI22_X1 U4639 ( .A1(n1243), .A2(\unit_decode/n4044 ), .B1(n1247), .B2(
        \unit_decode/n3940 ), .ZN(\unit_decode/n3298 ) );
  OAI221_X1 U4640 ( .B1(\unit_decode/n1592 ), .B2(n1190), .C1(
        \unit_decode/n1568 ), .C2(n1193), .A(\unit_decode/n3272 ), .ZN(
        \unit_decode/n3271 ) );
  AOI22_X1 U4641 ( .A1(n1196), .A2(\unit_decode/n4042 ), .B1(n1199), .B2(
        \unit_decode/n3754 ), .ZN(\unit_decode/n3272 ) );
  OAI221_X1 U4642 ( .B1(\unit_decode/n1688 ), .B2(n1238), .C1(
        \unit_decode/n1664 ), .C2(n1241), .A(\unit_decode/n3280 ), .ZN(
        \unit_decode/n3279 ) );
  AOI22_X1 U4643 ( .A1(n1244), .A2(\unit_decode/n4040 ), .B1(n1247), .B2(
        \unit_decode/n3934 ), .ZN(\unit_decode/n3280 ) );
  OAI221_X1 U4644 ( .B1(\unit_decode/n1593 ), .B2(n1190), .C1(
        \unit_decode/n1569 ), .C2(n1193), .A(\unit_decode/n3254 ), .ZN(
        \unit_decode/n3253 ) );
  AOI22_X1 U4645 ( .A1(n1196), .A2(\unit_decode/n4038 ), .B1(n1199), .B2(
        \unit_decode/n3748 ), .ZN(\unit_decode/n3254 ) );
  OAI221_X1 U4646 ( .B1(\unit_decode/n1689 ), .B2(n1238), .C1(
        \unit_decode/n1665 ), .C2(n1241), .A(\unit_decode/n3262 ), .ZN(
        \unit_decode/n3261 ) );
  AOI22_X1 U4647 ( .A1(n1244), .A2(\unit_decode/n4036 ), .B1(n1247), .B2(
        \unit_decode/n3928 ), .ZN(\unit_decode/n3262 ) );
  OAI221_X1 U4648 ( .B1(\unit_decode/n1594 ), .B2(n1190), .C1(
        \unit_decode/n1570 ), .C2(n1193), .A(\unit_decode/n3236 ), .ZN(
        \unit_decode/n3235 ) );
  AOI22_X1 U4649 ( .A1(n1196), .A2(\unit_decode/n4034 ), .B1(n1199), .B2(
        \unit_decode/n3742 ), .ZN(\unit_decode/n3236 ) );
  OAI221_X1 U4650 ( .B1(\unit_decode/n1690 ), .B2(n1238), .C1(
        \unit_decode/n1666 ), .C2(n1241), .A(\unit_decode/n3244 ), .ZN(
        \unit_decode/n3243 ) );
  AOI22_X1 U4651 ( .A1(n1244), .A2(\unit_decode/n4032 ), .B1(n1247), .B2(
        \unit_decode/n3922 ), .ZN(\unit_decode/n3244 ) );
  OAI221_X1 U4652 ( .B1(\unit_decode/n1595 ), .B2(n1190), .C1(
        \unit_decode/n1571 ), .C2(n1193), .A(\unit_decode/n3218 ), .ZN(
        \unit_decode/n3217 ) );
  AOI22_X1 U4653 ( .A1(n1196), .A2(\unit_decode/n4030 ), .B1(n1199), .B2(
        \unit_decode/n3736 ), .ZN(\unit_decode/n3218 ) );
  OAI221_X1 U4654 ( .B1(\unit_decode/n1691 ), .B2(n1238), .C1(
        \unit_decode/n1667 ), .C2(n1241), .A(\unit_decode/n3226 ), .ZN(
        \unit_decode/n3225 ) );
  AOI22_X1 U4655 ( .A1(n1244), .A2(\unit_decode/n4028 ), .B1(n1247), .B2(
        \unit_decode/n3916 ), .ZN(\unit_decode/n3226 ) );
  OAI221_X1 U4656 ( .B1(\unit_decode/n1596 ), .B2(n1190), .C1(
        \unit_decode/n1572 ), .C2(n1193), .A(\unit_decode/n3200 ), .ZN(
        \unit_decode/n3199 ) );
  AOI22_X1 U4657 ( .A1(n1196), .A2(\unit_decode/n4026 ), .B1(n1199), .B2(
        \unit_decode/n3730 ), .ZN(\unit_decode/n3200 ) );
  OAI221_X1 U4658 ( .B1(\unit_decode/n1692 ), .B2(n1238), .C1(
        \unit_decode/n1668 ), .C2(n1241), .A(\unit_decode/n3208 ), .ZN(
        \unit_decode/n3207 ) );
  AOI22_X1 U4659 ( .A1(n1244), .A2(\unit_decode/n4024 ), .B1(n1247), .B2(
        \unit_decode/n3910 ), .ZN(\unit_decode/n3208 ) );
  OAI221_X1 U4660 ( .B1(\unit_decode/n1597 ), .B2(n1190), .C1(
        \unit_decode/n1573 ), .C2(n1193), .A(\unit_decode/n3182 ), .ZN(
        \unit_decode/n3181 ) );
  AOI22_X1 U4661 ( .A1(n1196), .A2(\unit_decode/n4022 ), .B1(n1199), .B2(
        \unit_decode/n3724 ), .ZN(\unit_decode/n3182 ) );
  OAI221_X1 U4662 ( .B1(\unit_decode/n1693 ), .B2(n1238), .C1(
        \unit_decode/n1669 ), .C2(n1241), .A(\unit_decode/n3190 ), .ZN(
        \unit_decode/n3189 ) );
  AOI22_X1 U4663 ( .A1(n1244), .A2(\unit_decode/n4020 ), .B1(n1247), .B2(
        \unit_decode/n3904 ), .ZN(\unit_decode/n3190 ) );
  OAI221_X1 U4664 ( .B1(\unit_decode/n1598 ), .B2(n1190), .C1(
        \unit_decode/n1574 ), .C2(n1193), .A(\unit_decode/n3164 ), .ZN(
        \unit_decode/n3163 ) );
  AOI22_X1 U4665 ( .A1(n1196), .A2(\unit_decode/n4138 ), .B1(n1199), .B2(
        \unit_decode/n3718 ), .ZN(\unit_decode/n3164 ) );
  OAI221_X1 U4666 ( .B1(\unit_decode/n1694 ), .B2(n1238), .C1(
        \unit_decode/n1670 ), .C2(n1241), .A(\unit_decode/n3172 ), .ZN(
        \unit_decode/n3171 ) );
  AOI22_X1 U4667 ( .A1(n1244), .A2(\unit_decode/n4136 ), .B1(n1247), .B2(
        \unit_decode/n3898 ), .ZN(\unit_decode/n3172 ) );
  OAI221_X1 U4668 ( .B1(\unit_decode/n1599 ), .B2(n1190), .C1(
        \unit_decode/n1575 ), .C2(n1193), .A(\unit_decode/n3146 ), .ZN(
        \unit_decode/n3145 ) );
  AOI22_X1 U4669 ( .A1(n1196), .A2(\unit_decode/n4134 ), .B1(n1199), .B2(
        \unit_decode/n3712 ), .ZN(\unit_decode/n3146 ) );
  OAI221_X1 U4670 ( .B1(\unit_decode/n1695 ), .B2(n1238), .C1(
        \unit_decode/n1671 ), .C2(n1241), .A(\unit_decode/n3154 ), .ZN(
        \unit_decode/n3153 ) );
  AOI22_X1 U4671 ( .A1(n1244), .A2(\unit_decode/n4132 ), .B1(n1247), .B2(
        \unit_decode/n3892 ), .ZN(\unit_decode/n3154 ) );
  OAI221_X1 U4672 ( .B1(\unit_decode/n1600 ), .B2(n1190), .C1(
        \unit_decode/n1576 ), .C2(n1193), .A(\unit_decode/n3128 ), .ZN(
        \unit_decode/n3127 ) );
  AOI22_X1 U4673 ( .A1(n1196), .A2(\unit_decode/n4130 ), .B1(n1198), .B2(
        \unit_decode/n3706 ), .ZN(\unit_decode/n3128 ) );
  OAI221_X1 U4674 ( .B1(\unit_decode/n1696 ), .B2(n1238), .C1(
        \unit_decode/n1672 ), .C2(n1241), .A(\unit_decode/n3136 ), .ZN(
        \unit_decode/n3135 ) );
  AOI22_X1 U4675 ( .A1(n1244), .A2(\unit_decode/n4128 ), .B1(n1246), .B2(
        \unit_decode/n3886 ), .ZN(\unit_decode/n3136 ) );
  OAI221_X1 U4676 ( .B1(\unit_decode/n1601 ), .B2(n1190), .C1(
        \unit_decode/n1577 ), .C2(n1193), .A(\unit_decode/n3110 ), .ZN(
        \unit_decode/n3109 ) );
  AOI22_X1 U4677 ( .A1(n1196), .A2(\unit_decode/n4126 ), .B1(n1198), .B2(
        \unit_decode/n3700 ), .ZN(\unit_decode/n3110 ) );
  OAI221_X1 U4678 ( .B1(\unit_decode/n1697 ), .B2(n1238), .C1(
        \unit_decode/n1673 ), .C2(n1241), .A(\unit_decode/n3118 ), .ZN(
        \unit_decode/n3117 ) );
  AOI22_X1 U4679 ( .A1(n1244), .A2(\unit_decode/n4124 ), .B1(n1246), .B2(
        \unit_decode/n3880 ), .ZN(\unit_decode/n3118 ) );
  OAI221_X1 U4680 ( .B1(\unit_decode/n1602 ), .B2(n1190), .C1(
        \unit_decode/n1578 ), .C2(n1193), .A(\unit_decode/n3092 ), .ZN(
        \unit_decode/n3091 ) );
  AOI22_X1 U4681 ( .A1(n1196), .A2(\unit_decode/n4122 ), .B1(n1198), .B2(
        \unit_decode/n3694 ), .ZN(\unit_decode/n3092 ) );
  OAI221_X1 U4682 ( .B1(\unit_decode/n1698 ), .B2(n1238), .C1(
        \unit_decode/n1674 ), .C2(n1241), .A(\unit_decode/n3100 ), .ZN(
        \unit_decode/n3099 ) );
  AOI22_X1 U4683 ( .A1(n1244), .A2(\unit_decode/n4120 ), .B1(n1246), .B2(
        \unit_decode/n3874 ), .ZN(\unit_decode/n3100 ) );
  OAI221_X1 U4684 ( .B1(\unit_decode/n1603 ), .B2(n1190), .C1(
        \unit_decode/n1579 ), .C2(n1193), .A(\unit_decode/n3074 ), .ZN(
        \unit_decode/n3073 ) );
  AOI22_X1 U4685 ( .A1(n1196), .A2(\unit_decode/n4118 ), .B1(n1198), .B2(
        \unit_decode/n3688 ), .ZN(\unit_decode/n3074 ) );
  OAI221_X1 U4686 ( .B1(\unit_decode/n1699 ), .B2(n1238), .C1(
        \unit_decode/n1675 ), .C2(n1241), .A(\unit_decode/n3082 ), .ZN(
        \unit_decode/n3081 ) );
  AOI22_X1 U4687 ( .A1(n1244), .A2(\unit_decode/n4116 ), .B1(n1246), .B2(
        \unit_decode/n3868 ), .ZN(\unit_decode/n3082 ) );
  OAI221_X1 U4688 ( .B1(\unit_decode/n1806 ), .B2(n1107), .C1(
        \unit_decode/n1798 ), .C2(n1110), .A(\unit_decode/n2437 ), .ZN(
        \unit_decode/n2434 ) );
  AOI22_X1 U4689 ( .A1(n1113), .A2(\unit_decode/n4113 ), .B1(n1114), .B2(
        \unit_decode/n3681 ), .ZN(\unit_decode/n2437 ) );
  OAI221_X1 U4690 ( .B1(\unit_decode/n1838 ), .B2(n1155), .C1(
        \unit_decode/n1830 ), .C2(n1158), .A(\unit_decode/n2445 ), .ZN(
        \unit_decode/n2442 ) );
  AOI22_X1 U4691 ( .A1(n1161), .A2(\unit_decode/n4111 ), .B1(n1162), .B2(
        \unit_decode/n3861 ), .ZN(\unit_decode/n2445 ) );
  OAI221_X1 U4692 ( .B1(\unit_decode/n1805 ), .B2(n1107), .C1(
        \unit_decode/n1797 ), .C2(n1110), .A(\unit_decode/n2419 ), .ZN(
        \unit_decode/n2416 ) );
  AOI22_X1 U4693 ( .A1(n1113), .A2(\unit_decode/n4109 ), .B1(n1114), .B2(
        \unit_decode/n3675 ), .ZN(\unit_decode/n2419 ) );
  OAI221_X1 U4694 ( .B1(\unit_decode/n1837 ), .B2(n1155), .C1(
        \unit_decode/n1829 ), .C2(n1158), .A(\unit_decode/n2427 ), .ZN(
        \unit_decode/n2424 ) );
  AOI22_X1 U4695 ( .A1(n1161), .A2(\unit_decode/n4107 ), .B1(n1162), .B2(
        \unit_decode/n3855 ), .ZN(\unit_decode/n2427 ) );
  OAI221_X1 U4696 ( .B1(\unit_decode/n1804 ), .B2(n1107), .C1(
        \unit_decode/n1796 ), .C2(n1110), .A(\unit_decode/n2401 ), .ZN(
        \unit_decode/n2398 ) );
  AOI22_X1 U4697 ( .A1(n1113), .A2(\unit_decode/n4105 ), .B1(n1114), .B2(
        \unit_decode/n3669 ), .ZN(\unit_decode/n2401 ) );
  OAI221_X1 U4698 ( .B1(\unit_decode/n1836 ), .B2(n1155), .C1(
        \unit_decode/n1828 ), .C2(n1158), .A(\unit_decode/n2409 ), .ZN(
        \unit_decode/n2406 ) );
  AOI22_X1 U4699 ( .A1(n1161), .A2(\unit_decode/n4103 ), .B1(n1162), .B2(
        \unit_decode/n3849 ), .ZN(\unit_decode/n2409 ) );
  OAI221_X1 U4700 ( .B1(\unit_decode/n1803 ), .B2(n1107), .C1(
        \unit_decode/n1795 ), .C2(n1110), .A(\unit_decode/n2383 ), .ZN(
        \unit_decode/n2380 ) );
  AOI22_X1 U4701 ( .A1(n1113), .A2(\unit_decode/n4101 ), .B1(n1114), .B2(
        \unit_decode/n3663 ), .ZN(\unit_decode/n2383 ) );
  OAI221_X1 U4702 ( .B1(\unit_decode/n1835 ), .B2(n1155), .C1(
        \unit_decode/n1827 ), .C2(n1158), .A(\unit_decode/n2391 ), .ZN(
        \unit_decode/n2388 ) );
  AOI22_X1 U4703 ( .A1(n1161), .A2(\unit_decode/n4099 ), .B1(n1162), .B2(
        \unit_decode/n3843 ), .ZN(\unit_decode/n2391 ) );
  OAI221_X1 U4704 ( .B1(\unit_decode/n1802 ), .B2(n1107), .C1(
        \unit_decode/n1794 ), .C2(n1110), .A(\unit_decode/n2365 ), .ZN(
        \unit_decode/n2362 ) );
  AOI22_X1 U4705 ( .A1(n1113), .A2(\unit_decode/n4097 ), .B1(n1114), .B2(
        \unit_decode/n3657 ), .ZN(\unit_decode/n2365 ) );
  OAI221_X1 U4706 ( .B1(\unit_decode/n1834 ), .B2(n1155), .C1(
        \unit_decode/n1826 ), .C2(n1158), .A(\unit_decode/n2373 ), .ZN(
        \unit_decode/n2370 ) );
  AOI22_X1 U4707 ( .A1(n1161), .A2(\unit_decode/n4095 ), .B1(n1162), .B2(
        \unit_decode/n3837 ), .ZN(\unit_decode/n2373 ) );
  OAI221_X1 U4708 ( .B1(\unit_decode/n1801 ), .B2(n1107), .C1(
        \unit_decode/n1793 ), .C2(n1110), .A(\unit_decode/n2347 ), .ZN(
        \unit_decode/n2344 ) );
  AOI22_X1 U4709 ( .A1(n1113), .A2(\unit_decode/n4093 ), .B1(n1114), .B2(
        \unit_decode/n3651 ), .ZN(\unit_decode/n2347 ) );
  OAI221_X1 U4710 ( .B1(\unit_decode/n1833 ), .B2(n1155), .C1(
        \unit_decode/n1825 ), .C2(n1158), .A(\unit_decode/n2355 ), .ZN(
        \unit_decode/n2352 ) );
  AOI22_X1 U4711 ( .A1(n1161), .A2(\unit_decode/n4091 ), .B1(n1162), .B2(
        \unit_decode/n3831 ), .ZN(\unit_decode/n2355 ) );
  OAI221_X1 U4712 ( .B1(\unit_decode/n1800 ), .B2(n1107), .C1(
        \unit_decode/n1792 ), .C2(n1110), .A(\unit_decode/n2329 ), .ZN(
        \unit_decode/n2326 ) );
  AOI22_X1 U4713 ( .A1(n1113), .A2(\unit_decode/n4017 ), .B1(n1114), .B2(
        \unit_decode/n3633 ), .ZN(\unit_decode/n2329 ) );
  OAI221_X1 U4714 ( .B1(\unit_decode/n1832 ), .B2(n1155), .C1(
        \unit_decode/n1824 ), .C2(n1158), .A(\unit_decode/n2337 ), .ZN(
        \unit_decode/n2334 ) );
  AOI22_X1 U4715 ( .A1(n1161), .A2(\unit_decode/n4015 ), .B1(n1162), .B2(
        \unit_decode/n3645 ), .ZN(\unit_decode/n2337 ) );
  OAI221_X1 U4716 ( .B1(\unit_decode/n1799 ), .B2(n1107), .C1(
        \unit_decode/n1791 ), .C2(n1110), .A(\unit_decode/n2285 ), .ZN(
        \unit_decode/n2276 ) );
  AOI22_X1 U4717 ( .A1(n1113), .A2(\unit_decode/n4013 ), .B1(n1114), .B2(
        \unit_decode/n3627 ), .ZN(\unit_decode/n2285 ) );
  OAI221_X1 U4718 ( .B1(\unit_decode/n1831 ), .B2(n1155), .C1(
        \unit_decode/n1823 ), .C2(n1158), .A(\unit_decode/n2309 ), .ZN(
        \unit_decode/n2300 ) );
  AOI22_X1 U4719 ( .A1(n1161), .A2(\unit_decode/n4011 ), .B1(n1162), .B2(
        \unit_decode/n3639 ), .ZN(\unit_decode/n2309 ) );
  OAI221_X1 U4720 ( .B1(\unit_decode/n1806 ), .B2(n1203), .C1(
        \unit_decode/n1798 ), .C2(n1206), .A(\unit_decode/n3057 ), .ZN(
        \unit_decode/n3054 ) );
  AOI22_X1 U4721 ( .A1(n1209), .A2(\unit_decode/n4113 ), .B1(n1210), .B2(
        \unit_decode/n3681 ), .ZN(\unit_decode/n3057 ) );
  OAI221_X1 U4722 ( .B1(\unit_decode/n1838 ), .B2(n1251), .C1(
        \unit_decode/n1830 ), .C2(n1254), .A(\unit_decode/n3065 ), .ZN(
        \unit_decode/n3062 ) );
  AOI22_X1 U4723 ( .A1(n1257), .A2(\unit_decode/n4111 ), .B1(n1258), .B2(
        \unit_decode/n3861 ), .ZN(\unit_decode/n3065 ) );
  OAI221_X1 U4724 ( .B1(\unit_decode/n1805 ), .B2(n1203), .C1(
        \unit_decode/n1797 ), .C2(n1206), .A(\unit_decode/n3039 ), .ZN(
        \unit_decode/n3036 ) );
  AOI22_X1 U4725 ( .A1(n1209), .A2(\unit_decode/n4109 ), .B1(n1210), .B2(
        \unit_decode/n3675 ), .ZN(\unit_decode/n3039 ) );
  OAI221_X1 U4726 ( .B1(\unit_decode/n1837 ), .B2(n1251), .C1(
        \unit_decode/n1829 ), .C2(n1254), .A(\unit_decode/n3047 ), .ZN(
        \unit_decode/n3044 ) );
  AOI22_X1 U4727 ( .A1(n1257), .A2(\unit_decode/n4107 ), .B1(n1258), .B2(
        \unit_decode/n3855 ), .ZN(\unit_decode/n3047 ) );
  OAI221_X1 U4728 ( .B1(\unit_decode/n1804 ), .B2(n1203), .C1(
        \unit_decode/n1796 ), .C2(n1206), .A(\unit_decode/n3021 ), .ZN(
        \unit_decode/n3018 ) );
  AOI22_X1 U4729 ( .A1(n1209), .A2(\unit_decode/n4105 ), .B1(n1210), .B2(
        \unit_decode/n3669 ), .ZN(\unit_decode/n3021 ) );
  OAI221_X1 U4730 ( .B1(\unit_decode/n1836 ), .B2(n1251), .C1(
        \unit_decode/n1828 ), .C2(n1254), .A(\unit_decode/n3029 ), .ZN(
        \unit_decode/n3026 ) );
  AOI22_X1 U4731 ( .A1(n1257), .A2(\unit_decode/n4103 ), .B1(n1258), .B2(
        \unit_decode/n3849 ), .ZN(\unit_decode/n3029 ) );
  OAI221_X1 U4732 ( .B1(\unit_decode/n1803 ), .B2(n1203), .C1(
        \unit_decode/n1795 ), .C2(n1206), .A(\unit_decode/n3003 ), .ZN(
        \unit_decode/n3000 ) );
  AOI22_X1 U4733 ( .A1(n1209), .A2(\unit_decode/n4101 ), .B1(n1210), .B2(
        \unit_decode/n3663 ), .ZN(\unit_decode/n3003 ) );
  OAI221_X1 U4734 ( .B1(\unit_decode/n1835 ), .B2(n1251), .C1(
        \unit_decode/n1827 ), .C2(n1254), .A(\unit_decode/n3011 ), .ZN(
        \unit_decode/n3008 ) );
  AOI22_X1 U4735 ( .A1(n1257), .A2(\unit_decode/n4099 ), .B1(n1258), .B2(
        \unit_decode/n3843 ), .ZN(\unit_decode/n3011 ) );
  OAI221_X1 U4736 ( .B1(\unit_decode/n1802 ), .B2(n1203), .C1(
        \unit_decode/n1794 ), .C2(n1206), .A(\unit_decode/n2985 ), .ZN(
        \unit_decode/n2982 ) );
  AOI22_X1 U4737 ( .A1(n1209), .A2(\unit_decode/n4097 ), .B1(n1210), .B2(
        \unit_decode/n3657 ), .ZN(\unit_decode/n2985 ) );
  OAI221_X1 U4738 ( .B1(\unit_decode/n1834 ), .B2(n1251), .C1(
        \unit_decode/n1826 ), .C2(n1254), .A(\unit_decode/n2993 ), .ZN(
        \unit_decode/n2990 ) );
  AOI22_X1 U4739 ( .A1(n1257), .A2(\unit_decode/n4095 ), .B1(n1258), .B2(
        \unit_decode/n3837 ), .ZN(\unit_decode/n2993 ) );
  OAI221_X1 U4740 ( .B1(\unit_decode/n1801 ), .B2(n1203), .C1(
        \unit_decode/n1793 ), .C2(n1206), .A(\unit_decode/n2967 ), .ZN(
        \unit_decode/n2964 ) );
  AOI22_X1 U4741 ( .A1(n1209), .A2(\unit_decode/n4093 ), .B1(n1210), .B2(
        \unit_decode/n3651 ), .ZN(\unit_decode/n2967 ) );
  OAI221_X1 U4742 ( .B1(\unit_decode/n1833 ), .B2(n1251), .C1(
        \unit_decode/n1825 ), .C2(n1254), .A(\unit_decode/n2975 ), .ZN(
        \unit_decode/n2972 ) );
  AOI22_X1 U4743 ( .A1(n1257), .A2(\unit_decode/n4091 ), .B1(n1258), .B2(
        \unit_decode/n3831 ), .ZN(\unit_decode/n2975 ) );
  OAI221_X1 U4744 ( .B1(\unit_decode/n1800 ), .B2(n1203), .C1(
        \unit_decode/n1792 ), .C2(n1206), .A(\unit_decode/n2949 ), .ZN(
        \unit_decode/n2946 ) );
  AOI22_X1 U4745 ( .A1(n1209), .A2(\unit_decode/n4017 ), .B1(n1210), .B2(
        \unit_decode/n3633 ), .ZN(\unit_decode/n2949 ) );
  OAI221_X1 U4746 ( .B1(\unit_decode/n1832 ), .B2(n1251), .C1(
        \unit_decode/n1824 ), .C2(n1254), .A(\unit_decode/n2957 ), .ZN(
        \unit_decode/n2954 ) );
  AOI22_X1 U4747 ( .A1(n1257), .A2(\unit_decode/n4015 ), .B1(n1258), .B2(
        \unit_decode/n3645 ), .ZN(\unit_decode/n2957 ) );
  OAI221_X1 U4748 ( .B1(\unit_decode/n1799 ), .B2(n1203), .C1(
        \unit_decode/n1791 ), .C2(n1206), .A(\unit_decode/n2905 ), .ZN(
        \unit_decode/n2896 ) );
  AOI22_X1 U4749 ( .A1(n1209), .A2(\unit_decode/n4013 ), .B1(n1210), .B2(
        \unit_decode/n3627 ), .ZN(\unit_decode/n2905 ) );
  OAI221_X1 U4750 ( .B1(\unit_decode/n1831 ), .B2(n1251), .C1(
        \unit_decode/n1823 ), .C2(n1254), .A(\unit_decode/n2929 ), .ZN(
        \unit_decode/n2920 ) );
  AOI22_X1 U4751 ( .A1(n1257), .A2(\unit_decode/n4011 ), .B1(n1258), .B2(
        \unit_decode/n3639 ), .ZN(\unit_decode/n2929 ) );
  OAI221_X1 U4752 ( .B1(\unit_decode/n1388 ), .B2(n1105), .C1(
        \unit_decode/n1365 ), .C2(n1108), .A(\unit_decode/n2874 ), .ZN(
        \unit_decode/n2866 ) );
  AOI22_X1 U4753 ( .A1(n1111), .A2(\unit_decode/n4089 ), .B1(n1116), .B2(
        \unit_decode/n3825 ), .ZN(\unit_decode/n2874 ) );
  OAI221_X1 U4754 ( .B1(\unit_decode/n1484 ), .B2(n1153), .C1(
        \unit_decode/n1460 ), .C2(n1156), .A(\unit_decode/n2886 ), .ZN(
        \unit_decode/n2882 ) );
  AOI22_X1 U4755 ( .A1(n1159), .A2(\unit_decode/n4087 ), .B1(n1164), .B2(
        \unit_decode/n4005 ), .ZN(\unit_decode/n2886 ) );
  OAI221_X1 U4756 ( .B1(\unit_decode/n1389 ), .B2(n1105), .C1(
        \unit_decode/n1366 ), .C2(n1108), .A(\unit_decode/n2851 ), .ZN(
        \unit_decode/n2848 ) );
  AOI22_X1 U4757 ( .A1(n1111), .A2(\unit_decode/n4085 ), .B1(n1116), .B2(
        \unit_decode/n3819 ), .ZN(\unit_decode/n2851 ) );
  OAI221_X1 U4758 ( .B1(\unit_decode/n1485 ), .B2(n1153), .C1(
        \unit_decode/n1461 ), .C2(n1156), .A(\unit_decode/n2859 ), .ZN(
        \unit_decode/n2856 ) );
  AOI22_X1 U4759 ( .A1(n1159), .A2(\unit_decode/n4083 ), .B1(n1164), .B2(
        \unit_decode/n3999 ), .ZN(\unit_decode/n2859 ) );
  OAI221_X1 U4760 ( .B1(\unit_decode/n1390 ), .B2(n1105), .C1(
        \unit_decode/n1367 ), .C2(n1108), .A(\unit_decode/n2833 ), .ZN(
        \unit_decode/n2830 ) );
  AOI22_X1 U4761 ( .A1(n1111), .A2(\unit_decode/n4081 ), .B1(n1116), .B2(
        \unit_decode/n3813 ), .ZN(\unit_decode/n2833 ) );
  OAI221_X1 U4762 ( .B1(\unit_decode/n1486 ), .B2(n1153), .C1(
        \unit_decode/n1462 ), .C2(n1156), .A(\unit_decode/n2841 ), .ZN(
        \unit_decode/n2838 ) );
  AOI22_X1 U4763 ( .A1(n1159), .A2(\unit_decode/n4079 ), .B1(n1164), .B2(
        \unit_decode/n3993 ), .ZN(\unit_decode/n2841 ) );
  OAI221_X1 U4764 ( .B1(\unit_decode/n1391 ), .B2(n1105), .C1(
        \unit_decode/n1368 ), .C2(n1108), .A(\unit_decode/n2815 ), .ZN(
        \unit_decode/n2812 ) );
  AOI22_X1 U4765 ( .A1(n1111), .A2(\unit_decode/n4077 ), .B1(n1116), .B2(
        \unit_decode/n3807 ), .ZN(\unit_decode/n2815 ) );
  OAI221_X1 U4766 ( .B1(\unit_decode/n1487 ), .B2(n1153), .C1(
        \unit_decode/n1463 ), .C2(n1156), .A(\unit_decode/n2823 ), .ZN(
        \unit_decode/n2820 ) );
  AOI22_X1 U4767 ( .A1(n1159), .A2(\unit_decode/n4075 ), .B1(n1164), .B2(
        \unit_decode/n3987 ), .ZN(\unit_decode/n2823 ) );
  OAI221_X1 U4768 ( .B1(\unit_decode/n1392 ), .B2(n1105), .C1(
        \unit_decode/n1369 ), .C2(n1108), .A(\unit_decode/n2797 ), .ZN(
        \unit_decode/n2794 ) );
  AOI22_X1 U4769 ( .A1(n1111), .A2(\unit_decode/n4073 ), .B1(n1116), .B2(
        \unit_decode/n3801 ), .ZN(\unit_decode/n2797 ) );
  OAI221_X1 U4770 ( .B1(\unit_decode/n1488 ), .B2(n1153), .C1(
        \unit_decode/n1464 ), .C2(n1156), .A(\unit_decode/n2805 ), .ZN(
        \unit_decode/n2802 ) );
  AOI22_X1 U4771 ( .A1(n1159), .A2(\unit_decode/n4071 ), .B1(n1164), .B2(
        \unit_decode/n3981 ), .ZN(\unit_decode/n2805 ) );
  OAI221_X1 U4772 ( .B1(\unit_decode/n1393 ), .B2(n1105), .C1(
        \unit_decode/n1370 ), .C2(n1108), .A(\unit_decode/n2779 ), .ZN(
        \unit_decode/n2776 ) );
  AOI22_X1 U4773 ( .A1(n1111), .A2(\unit_decode/n4069 ), .B1(n1116), .B2(
        \unit_decode/n3795 ), .ZN(\unit_decode/n2779 ) );
  OAI221_X1 U4774 ( .B1(\unit_decode/n1489 ), .B2(n1153), .C1(
        \unit_decode/n1465 ), .C2(n1156), .A(\unit_decode/n2787 ), .ZN(
        \unit_decode/n2784 ) );
  AOI22_X1 U4775 ( .A1(n1159), .A2(\unit_decode/n4067 ), .B1(n1164), .B2(
        \unit_decode/n3975 ), .ZN(\unit_decode/n2787 ) );
  OAI221_X1 U4776 ( .B1(\unit_decode/n1394 ), .B2(n1105), .C1(
        \unit_decode/n1371 ), .C2(n1108), .A(\unit_decode/n2761 ), .ZN(
        \unit_decode/n2758 ) );
  AOI22_X1 U4777 ( .A1(n1111), .A2(\unit_decode/n4065 ), .B1(n1116), .B2(
        \unit_decode/n3789 ), .ZN(\unit_decode/n2761 ) );
  OAI221_X1 U4778 ( .B1(\unit_decode/n1490 ), .B2(n1153), .C1(
        \unit_decode/n1466 ), .C2(n1156), .A(\unit_decode/n2769 ), .ZN(
        \unit_decode/n2766 ) );
  AOI22_X1 U4779 ( .A1(n1159), .A2(\unit_decode/n4063 ), .B1(n1164), .B2(
        \unit_decode/n3969 ), .ZN(\unit_decode/n2769 ) );
  OAI221_X1 U4780 ( .B1(\unit_decode/n1395 ), .B2(n1105), .C1(
        \unit_decode/n1372 ), .C2(n1108), .A(\unit_decode/n2743 ), .ZN(
        \unit_decode/n2740 ) );
  AOI22_X1 U4781 ( .A1(n1111), .A2(\unit_decode/n4061 ), .B1(n1116), .B2(
        \unit_decode/n3783 ), .ZN(\unit_decode/n2743 ) );
  OAI221_X1 U4782 ( .B1(\unit_decode/n1491 ), .B2(n1153), .C1(
        \unit_decode/n1467 ), .C2(n1156), .A(\unit_decode/n2751 ), .ZN(
        \unit_decode/n2748 ) );
  AOI22_X1 U4783 ( .A1(n1159), .A2(\unit_decode/n4059 ), .B1(n1164), .B2(
        \unit_decode/n3963 ), .ZN(\unit_decode/n2751 ) );
  OAI221_X1 U4784 ( .B1(\unit_decode/n1396 ), .B2(n1105), .C1(
        \unit_decode/n1373 ), .C2(n1108), .A(\unit_decode/n2725 ), .ZN(
        \unit_decode/n2722 ) );
  AOI22_X1 U4785 ( .A1(n1111), .A2(\unit_decode/n4057 ), .B1(n1115), .B2(
        \unit_decode/n3777 ), .ZN(\unit_decode/n2725 ) );
  OAI221_X1 U4786 ( .B1(\unit_decode/n1492 ), .B2(n1153), .C1(
        \unit_decode/n1468 ), .C2(n1156), .A(\unit_decode/n2733 ), .ZN(
        \unit_decode/n2730 ) );
  AOI22_X1 U4787 ( .A1(n1159), .A2(\unit_decode/n4055 ), .B1(n1163), .B2(
        \unit_decode/n3957 ), .ZN(\unit_decode/n2733 ) );
  OAI221_X1 U4788 ( .B1(\unit_decode/n1397 ), .B2(n1105), .C1(
        \unit_decode/n1374 ), .C2(n1108), .A(\unit_decode/n2707 ), .ZN(
        \unit_decode/n2704 ) );
  AOI22_X1 U4789 ( .A1(n1111), .A2(\unit_decode/n4053 ), .B1(n1115), .B2(
        \unit_decode/n3771 ), .ZN(\unit_decode/n2707 ) );
  OAI221_X1 U4790 ( .B1(\unit_decode/n1493 ), .B2(n1153), .C1(
        \unit_decode/n1469 ), .C2(n1156), .A(\unit_decode/n2715 ), .ZN(
        \unit_decode/n2712 ) );
  AOI22_X1 U4791 ( .A1(n1159), .A2(\unit_decode/n4051 ), .B1(n1163), .B2(
        \unit_decode/n3951 ), .ZN(\unit_decode/n2715 ) );
  OAI221_X1 U4792 ( .B1(\unit_decode/n1398 ), .B2(n1105), .C1(
        \unit_decode/n1375 ), .C2(n1108), .A(\unit_decode/n2689 ), .ZN(
        \unit_decode/n2686 ) );
  AOI22_X1 U4793 ( .A1(n1111), .A2(\unit_decode/n4049 ), .B1(n1115), .B2(
        \unit_decode/n3765 ), .ZN(\unit_decode/n2689 ) );
  OAI221_X1 U4794 ( .B1(\unit_decode/n1494 ), .B2(n1153), .C1(
        \unit_decode/n1470 ), .C2(n1156), .A(\unit_decode/n2697 ), .ZN(
        \unit_decode/n2694 ) );
  AOI22_X1 U4795 ( .A1(n1159), .A2(\unit_decode/n4047 ), .B1(n1163), .B2(
        \unit_decode/n3945 ), .ZN(\unit_decode/n2697 ) );
  OAI221_X1 U4796 ( .B1(\unit_decode/n1399 ), .B2(n1105), .C1(
        \unit_decode/n1376 ), .C2(n1108), .A(\unit_decode/n2671 ), .ZN(
        \unit_decode/n2668 ) );
  AOI22_X1 U4797 ( .A1(n1111), .A2(\unit_decode/n4045 ), .B1(n1115), .B2(
        \unit_decode/n3759 ), .ZN(\unit_decode/n2671 ) );
  OAI221_X1 U4798 ( .B1(\unit_decode/n1495 ), .B2(n1153), .C1(
        \unit_decode/n1471 ), .C2(n1156), .A(\unit_decode/n2679 ), .ZN(
        \unit_decode/n2676 ) );
  AOI22_X1 U4799 ( .A1(n1159), .A2(\unit_decode/n4043 ), .B1(n1163), .B2(
        \unit_decode/n3939 ), .ZN(\unit_decode/n2679 ) );
  OAI221_X1 U4800 ( .B1(\unit_decode/n1400 ), .B2(n1106), .C1(
        \unit_decode/n1377 ), .C2(n1109), .A(\unit_decode/n2653 ), .ZN(
        \unit_decode/n2650 ) );
  AOI22_X1 U4801 ( .A1(n1112), .A2(\unit_decode/n4041 ), .B1(n1115), .B2(
        \unit_decode/n3753 ), .ZN(\unit_decode/n2653 ) );
  OAI221_X1 U4802 ( .B1(\unit_decode/n1496 ), .B2(n1154), .C1(
        \unit_decode/n1472 ), .C2(n1157), .A(\unit_decode/n2661 ), .ZN(
        \unit_decode/n2658 ) );
  AOI22_X1 U4803 ( .A1(n1160), .A2(\unit_decode/n4039 ), .B1(n1163), .B2(
        \unit_decode/n3933 ), .ZN(\unit_decode/n2661 ) );
  OAI221_X1 U4804 ( .B1(\unit_decode/n1401 ), .B2(n1106), .C1(
        \unit_decode/n1378 ), .C2(n1109), .A(\unit_decode/n2635 ), .ZN(
        \unit_decode/n2632 ) );
  AOI22_X1 U4805 ( .A1(n1112), .A2(\unit_decode/n4037 ), .B1(n1115), .B2(
        \unit_decode/n3747 ), .ZN(\unit_decode/n2635 ) );
  OAI221_X1 U4806 ( .B1(\unit_decode/n1497 ), .B2(n1154), .C1(
        \unit_decode/n1473 ), .C2(n1157), .A(\unit_decode/n2643 ), .ZN(
        \unit_decode/n2640 ) );
  AOI22_X1 U4807 ( .A1(n1160), .A2(\unit_decode/n4035 ), .B1(n1163), .B2(
        \unit_decode/n3927 ), .ZN(\unit_decode/n2643 ) );
  OAI221_X1 U4808 ( .B1(\unit_decode/n1402 ), .B2(n1106), .C1(
        \unit_decode/n1379 ), .C2(n1109), .A(\unit_decode/n2617 ), .ZN(
        \unit_decode/n2614 ) );
  AOI22_X1 U4809 ( .A1(n1112), .A2(\unit_decode/n4033 ), .B1(n1115), .B2(
        \unit_decode/n3741 ), .ZN(\unit_decode/n2617 ) );
  OAI221_X1 U4810 ( .B1(\unit_decode/n1498 ), .B2(n1154), .C1(
        \unit_decode/n1474 ), .C2(n1157), .A(\unit_decode/n2625 ), .ZN(
        \unit_decode/n2622 ) );
  AOI22_X1 U4811 ( .A1(n1160), .A2(\unit_decode/n4031 ), .B1(n1163), .B2(
        \unit_decode/n3921 ), .ZN(\unit_decode/n2625 ) );
  OAI221_X1 U4812 ( .B1(\unit_decode/n1403 ), .B2(n1106), .C1(
        \unit_decode/n1380 ), .C2(n1109), .A(\unit_decode/n2599 ), .ZN(
        \unit_decode/n2596 ) );
  AOI22_X1 U4813 ( .A1(n1112), .A2(\unit_decode/n4029 ), .B1(n1115), .B2(
        \unit_decode/n3735 ), .ZN(\unit_decode/n2599 ) );
  OAI221_X1 U4814 ( .B1(\unit_decode/n1499 ), .B2(n1154), .C1(
        \unit_decode/n1475 ), .C2(n1157), .A(\unit_decode/n2607 ), .ZN(
        \unit_decode/n2604 ) );
  AOI22_X1 U4815 ( .A1(n1160), .A2(\unit_decode/n4027 ), .B1(n1163), .B2(
        \unit_decode/n3915 ), .ZN(\unit_decode/n2607 ) );
  OAI221_X1 U4816 ( .B1(\unit_decode/n1404 ), .B2(n1106), .C1(
        \unit_decode/n1381 ), .C2(n1109), .A(\unit_decode/n2581 ), .ZN(
        \unit_decode/n2578 ) );
  AOI22_X1 U4817 ( .A1(n1112), .A2(\unit_decode/n4025 ), .B1(n1115), .B2(
        \unit_decode/n3729 ), .ZN(\unit_decode/n2581 ) );
  OAI221_X1 U4818 ( .B1(\unit_decode/n1500 ), .B2(n1154), .C1(
        \unit_decode/n1476 ), .C2(n1157), .A(\unit_decode/n2589 ), .ZN(
        \unit_decode/n2586 ) );
  AOI22_X1 U4819 ( .A1(n1160), .A2(\unit_decode/n4023 ), .B1(n1163), .B2(
        \unit_decode/n3909 ), .ZN(\unit_decode/n2589 ) );
  OAI221_X1 U4820 ( .B1(\unit_decode/n1405 ), .B2(n1106), .C1(
        \unit_decode/n1382 ), .C2(n1109), .A(\unit_decode/n2563 ), .ZN(
        \unit_decode/n2560 ) );
  AOI22_X1 U4821 ( .A1(n1112), .A2(\unit_decode/n4021 ), .B1(n1115), .B2(
        \unit_decode/n3723 ), .ZN(\unit_decode/n2563 ) );
  OAI221_X1 U4822 ( .B1(\unit_decode/n1501 ), .B2(n1154), .C1(
        \unit_decode/n1477 ), .C2(n1157), .A(\unit_decode/n2571 ), .ZN(
        \unit_decode/n2568 ) );
  AOI22_X1 U4823 ( .A1(n1160), .A2(\unit_decode/n4019 ), .B1(n1163), .B2(
        \unit_decode/n3903 ), .ZN(\unit_decode/n2571 ) );
  OAI221_X1 U4824 ( .B1(\unit_decode/n1406 ), .B2(n1106), .C1(
        \unit_decode/n1383 ), .C2(n1109), .A(\unit_decode/n2545 ), .ZN(
        \unit_decode/n2542 ) );
  AOI22_X1 U4825 ( .A1(n1112), .A2(\unit_decode/n4137 ), .B1(n1115), .B2(
        \unit_decode/n3717 ), .ZN(\unit_decode/n2545 ) );
  OAI221_X1 U4826 ( .B1(\unit_decode/n1502 ), .B2(n1154), .C1(
        \unit_decode/n1478 ), .C2(n1157), .A(\unit_decode/n2553 ), .ZN(
        \unit_decode/n2550 ) );
  AOI22_X1 U4827 ( .A1(n1160), .A2(\unit_decode/n4135 ), .B1(n1163), .B2(
        \unit_decode/n3897 ), .ZN(\unit_decode/n2553 ) );
  OAI221_X1 U4828 ( .B1(\unit_decode/n1407 ), .B2(n1106), .C1(
        \unit_decode/n1384 ), .C2(n1109), .A(\unit_decode/n2527 ), .ZN(
        \unit_decode/n2524 ) );
  AOI22_X1 U4829 ( .A1(n1112), .A2(\unit_decode/n4133 ), .B1(n1115), .B2(
        \unit_decode/n3711 ), .ZN(\unit_decode/n2527 ) );
  OAI221_X1 U4830 ( .B1(\unit_decode/n1503 ), .B2(n1154), .C1(
        \unit_decode/n1479 ), .C2(n1157), .A(\unit_decode/n2535 ), .ZN(
        \unit_decode/n2532 ) );
  AOI22_X1 U4831 ( .A1(n1160), .A2(\unit_decode/n4131 ), .B1(n1163), .B2(
        \unit_decode/n3891 ), .ZN(\unit_decode/n2535 ) );
  OAI221_X1 U4832 ( .B1(\unit_decode/n1408 ), .B2(n1106), .C1(
        \unit_decode/n1385 ), .C2(n1109), .A(\unit_decode/n2509 ), .ZN(
        \unit_decode/n2506 ) );
  AOI22_X1 U4833 ( .A1(n1112), .A2(\unit_decode/n4129 ), .B1(n1114), .B2(
        \unit_decode/n3705 ), .ZN(\unit_decode/n2509 ) );
  OAI221_X1 U4834 ( .B1(\unit_decode/n1504 ), .B2(n1154), .C1(
        \unit_decode/n1480 ), .C2(n1157), .A(\unit_decode/n2517 ), .ZN(
        \unit_decode/n2514 ) );
  AOI22_X1 U4835 ( .A1(n1160), .A2(\unit_decode/n4127 ), .B1(n1162), .B2(
        \unit_decode/n3885 ), .ZN(\unit_decode/n2517 ) );
  OAI221_X1 U4836 ( .B1(\unit_decode/n1409 ), .B2(n1106), .C1(
        \unit_decode/n1386 ), .C2(n1109), .A(\unit_decode/n2491 ), .ZN(
        \unit_decode/n2488 ) );
  AOI22_X1 U4837 ( .A1(n1112), .A2(\unit_decode/n4125 ), .B1(n1114), .B2(
        \unit_decode/n3699 ), .ZN(\unit_decode/n2491 ) );
  OAI221_X1 U4838 ( .B1(\unit_decode/n1505 ), .B2(n1154), .C1(
        \unit_decode/n1481 ), .C2(n1157), .A(\unit_decode/n2499 ), .ZN(
        \unit_decode/n2496 ) );
  AOI22_X1 U4839 ( .A1(n1160), .A2(\unit_decode/n4123 ), .B1(n1162), .B2(
        \unit_decode/n3879 ), .ZN(\unit_decode/n2499 ) );
  OAI221_X1 U4840 ( .B1(\unit_decode/n1410 ), .B2(n1106), .C1(
        \unit_decode/n1387 ), .C2(n1109), .A(\unit_decode/n2473 ), .ZN(
        \unit_decode/n2470 ) );
  AOI22_X1 U4841 ( .A1(n1112), .A2(\unit_decode/n4121 ), .B1(n1114), .B2(
        \unit_decode/n3693 ), .ZN(\unit_decode/n2473 ) );
  OAI221_X1 U4842 ( .B1(\unit_decode/n1506 ), .B2(n1154), .C1(
        \unit_decode/n1482 ), .C2(n1157), .A(\unit_decode/n2481 ), .ZN(
        \unit_decode/n2478 ) );
  AOI22_X1 U4843 ( .A1(n1160), .A2(\unit_decode/n4119 ), .B1(n1162), .B2(
        \unit_decode/n3873 ), .ZN(\unit_decode/n2481 ) );
  OAI221_X1 U4844 ( .B1(\unit_decode/n1411 ), .B2(n1106), .C1(
        \unit_decode/n2084 ), .C2(n1109), .A(\unit_decode/n2455 ), .ZN(
        \unit_decode/n2452 ) );
  AOI22_X1 U4845 ( .A1(n1112), .A2(\unit_decode/n4117 ), .B1(n1114), .B2(
        \unit_decode/n3687 ), .ZN(\unit_decode/n2455 ) );
  OAI221_X1 U4846 ( .B1(\unit_decode/n1507 ), .B2(n1154), .C1(
        \unit_decode/n1483 ), .C2(n1157), .A(\unit_decode/n2463 ), .ZN(
        \unit_decode/n2460 ) );
  AOI22_X1 U4847 ( .A1(n1160), .A2(\unit_decode/n4115 ), .B1(n1162), .B2(
        \unit_decode/n3867 ), .ZN(\unit_decode/n2463 ) );
  OAI221_X1 U4848 ( .B1(\unit_decode/n1388 ), .B2(n1201), .C1(
        \unit_decode/n1365 ), .C2(n1204), .A(\unit_decode/n3494 ), .ZN(
        \unit_decode/n3486 ) );
  AOI22_X1 U4849 ( .A1(n1207), .A2(\unit_decode/n4089 ), .B1(n1212), .B2(
        \unit_decode/n3825 ), .ZN(\unit_decode/n3494 ) );
  OAI221_X1 U4850 ( .B1(\unit_decode/n1484 ), .B2(n1249), .C1(
        \unit_decode/n1460 ), .C2(n1252), .A(\unit_decode/n3506 ), .ZN(
        \unit_decode/n3502 ) );
  AOI22_X1 U4851 ( .A1(n1255), .A2(\unit_decode/n4087 ), .B1(n1260), .B2(
        \unit_decode/n4005 ), .ZN(\unit_decode/n3506 ) );
  OAI221_X1 U4852 ( .B1(\unit_decode/n1389 ), .B2(n1201), .C1(
        \unit_decode/n1366 ), .C2(n1204), .A(\unit_decode/n3471 ), .ZN(
        \unit_decode/n3468 ) );
  AOI22_X1 U4853 ( .A1(n1207), .A2(\unit_decode/n4085 ), .B1(n1212), .B2(
        \unit_decode/n3819 ), .ZN(\unit_decode/n3471 ) );
  OAI221_X1 U4854 ( .B1(\unit_decode/n1485 ), .B2(n1249), .C1(
        \unit_decode/n1461 ), .C2(n1252), .A(\unit_decode/n3479 ), .ZN(
        \unit_decode/n3476 ) );
  AOI22_X1 U4855 ( .A1(n1255), .A2(\unit_decode/n4083 ), .B1(n1260), .B2(
        \unit_decode/n3999 ), .ZN(\unit_decode/n3479 ) );
  OAI221_X1 U4856 ( .B1(\unit_decode/n1390 ), .B2(n1201), .C1(
        \unit_decode/n1367 ), .C2(n1204), .A(\unit_decode/n3453 ), .ZN(
        \unit_decode/n3450 ) );
  AOI22_X1 U4857 ( .A1(n1207), .A2(\unit_decode/n4081 ), .B1(n1212), .B2(
        \unit_decode/n3813 ), .ZN(\unit_decode/n3453 ) );
  OAI221_X1 U4858 ( .B1(\unit_decode/n1486 ), .B2(n1249), .C1(
        \unit_decode/n1462 ), .C2(n1252), .A(\unit_decode/n3461 ), .ZN(
        \unit_decode/n3458 ) );
  AOI22_X1 U4859 ( .A1(n1255), .A2(\unit_decode/n4079 ), .B1(n1260), .B2(
        \unit_decode/n3993 ), .ZN(\unit_decode/n3461 ) );
  OAI221_X1 U4860 ( .B1(\unit_decode/n1391 ), .B2(n1201), .C1(
        \unit_decode/n1368 ), .C2(n1204), .A(\unit_decode/n3435 ), .ZN(
        \unit_decode/n3432 ) );
  AOI22_X1 U4861 ( .A1(n1207), .A2(\unit_decode/n4077 ), .B1(n1212), .B2(
        \unit_decode/n3807 ), .ZN(\unit_decode/n3435 ) );
  OAI221_X1 U4862 ( .B1(\unit_decode/n1487 ), .B2(n1249), .C1(
        \unit_decode/n1463 ), .C2(n1252), .A(\unit_decode/n3443 ), .ZN(
        \unit_decode/n3440 ) );
  AOI22_X1 U4863 ( .A1(n1255), .A2(\unit_decode/n4075 ), .B1(n1260), .B2(
        \unit_decode/n3987 ), .ZN(\unit_decode/n3443 ) );
  OAI221_X1 U4864 ( .B1(\unit_decode/n1392 ), .B2(n1201), .C1(
        \unit_decode/n1369 ), .C2(n1204), .A(\unit_decode/n3417 ), .ZN(
        \unit_decode/n3414 ) );
  AOI22_X1 U4865 ( .A1(n1207), .A2(\unit_decode/n4073 ), .B1(n1212), .B2(
        \unit_decode/n3801 ), .ZN(\unit_decode/n3417 ) );
  OAI221_X1 U4866 ( .B1(\unit_decode/n1488 ), .B2(n1249), .C1(
        \unit_decode/n1464 ), .C2(n1252), .A(\unit_decode/n3425 ), .ZN(
        \unit_decode/n3422 ) );
  AOI22_X1 U4867 ( .A1(n1255), .A2(\unit_decode/n4071 ), .B1(n1260), .B2(
        \unit_decode/n3981 ), .ZN(\unit_decode/n3425 ) );
  OAI221_X1 U4868 ( .B1(\unit_decode/n1393 ), .B2(n1201), .C1(
        \unit_decode/n1370 ), .C2(n1204), .A(\unit_decode/n3399 ), .ZN(
        \unit_decode/n3396 ) );
  AOI22_X1 U4869 ( .A1(n1207), .A2(\unit_decode/n4069 ), .B1(n1212), .B2(
        \unit_decode/n3795 ), .ZN(\unit_decode/n3399 ) );
  OAI221_X1 U4870 ( .B1(\unit_decode/n1489 ), .B2(n1249), .C1(
        \unit_decode/n1465 ), .C2(n1252), .A(\unit_decode/n3407 ), .ZN(
        \unit_decode/n3404 ) );
  AOI22_X1 U4871 ( .A1(n1255), .A2(\unit_decode/n4067 ), .B1(n1260), .B2(
        \unit_decode/n3975 ), .ZN(\unit_decode/n3407 ) );
  OAI221_X1 U4872 ( .B1(\unit_decode/n1394 ), .B2(n1201), .C1(
        \unit_decode/n1371 ), .C2(n1204), .A(\unit_decode/n3381 ), .ZN(
        \unit_decode/n3378 ) );
  AOI22_X1 U4873 ( .A1(n1207), .A2(\unit_decode/n4065 ), .B1(n1212), .B2(
        \unit_decode/n3789 ), .ZN(\unit_decode/n3381 ) );
  OAI221_X1 U4874 ( .B1(\unit_decode/n1490 ), .B2(n1249), .C1(
        \unit_decode/n1466 ), .C2(n1252), .A(\unit_decode/n3389 ), .ZN(
        \unit_decode/n3386 ) );
  AOI22_X1 U4875 ( .A1(n1255), .A2(\unit_decode/n4063 ), .B1(n1260), .B2(
        \unit_decode/n3969 ), .ZN(\unit_decode/n3389 ) );
  OAI221_X1 U4876 ( .B1(\unit_decode/n1395 ), .B2(n1201), .C1(
        \unit_decode/n1372 ), .C2(n1204), .A(\unit_decode/n3363 ), .ZN(
        \unit_decode/n3360 ) );
  AOI22_X1 U4877 ( .A1(n1207), .A2(\unit_decode/n4061 ), .B1(n1212), .B2(
        \unit_decode/n3783 ), .ZN(\unit_decode/n3363 ) );
  OAI221_X1 U4878 ( .B1(\unit_decode/n1491 ), .B2(n1249), .C1(
        \unit_decode/n1467 ), .C2(n1252), .A(\unit_decode/n3371 ), .ZN(
        \unit_decode/n3368 ) );
  AOI22_X1 U4879 ( .A1(n1255), .A2(\unit_decode/n4059 ), .B1(n1260), .B2(
        \unit_decode/n3963 ), .ZN(\unit_decode/n3371 ) );
  OAI221_X1 U4880 ( .B1(\unit_decode/n1396 ), .B2(n1201), .C1(
        \unit_decode/n1373 ), .C2(n1204), .A(\unit_decode/n3345 ), .ZN(
        \unit_decode/n3342 ) );
  AOI22_X1 U4881 ( .A1(n1207), .A2(\unit_decode/n4057 ), .B1(n1211), .B2(
        \unit_decode/n3777 ), .ZN(\unit_decode/n3345 ) );
  OAI221_X1 U4882 ( .B1(\unit_decode/n1492 ), .B2(n1249), .C1(
        \unit_decode/n1468 ), .C2(n1252), .A(\unit_decode/n3353 ), .ZN(
        \unit_decode/n3350 ) );
  AOI22_X1 U4883 ( .A1(n1255), .A2(\unit_decode/n4055 ), .B1(n1259), .B2(
        \unit_decode/n3957 ), .ZN(\unit_decode/n3353 ) );
  OAI221_X1 U4884 ( .B1(\unit_decode/n1397 ), .B2(n1201), .C1(
        \unit_decode/n1374 ), .C2(n1204), .A(\unit_decode/n3327 ), .ZN(
        \unit_decode/n3324 ) );
  AOI22_X1 U4885 ( .A1(n1207), .A2(\unit_decode/n4053 ), .B1(n1211), .B2(
        \unit_decode/n3771 ), .ZN(\unit_decode/n3327 ) );
  OAI221_X1 U4886 ( .B1(\unit_decode/n1493 ), .B2(n1249), .C1(
        \unit_decode/n1469 ), .C2(n1252), .A(\unit_decode/n3335 ), .ZN(
        \unit_decode/n3332 ) );
  AOI22_X1 U4887 ( .A1(n1255), .A2(\unit_decode/n4051 ), .B1(n1259), .B2(
        \unit_decode/n3951 ), .ZN(\unit_decode/n3335 ) );
  OAI221_X1 U4888 ( .B1(\unit_decode/n1398 ), .B2(n1201), .C1(
        \unit_decode/n1375 ), .C2(n1204), .A(\unit_decode/n3309 ), .ZN(
        \unit_decode/n3306 ) );
  AOI22_X1 U4889 ( .A1(n1207), .A2(\unit_decode/n4049 ), .B1(n1211), .B2(
        \unit_decode/n3765 ), .ZN(\unit_decode/n3309 ) );
  OAI221_X1 U4890 ( .B1(\unit_decode/n1494 ), .B2(n1249), .C1(
        \unit_decode/n1470 ), .C2(n1252), .A(\unit_decode/n3317 ), .ZN(
        \unit_decode/n3314 ) );
  AOI22_X1 U4891 ( .A1(n1255), .A2(\unit_decode/n4047 ), .B1(n1259), .B2(
        \unit_decode/n3945 ), .ZN(\unit_decode/n3317 ) );
  OAI221_X1 U4892 ( .B1(\unit_decode/n1399 ), .B2(n1201), .C1(
        \unit_decode/n1376 ), .C2(n1204), .A(\unit_decode/n3291 ), .ZN(
        \unit_decode/n3288 ) );
  AOI22_X1 U4893 ( .A1(n1207), .A2(\unit_decode/n4045 ), .B1(n1211), .B2(
        \unit_decode/n3759 ), .ZN(\unit_decode/n3291 ) );
  OAI221_X1 U4894 ( .B1(\unit_decode/n1495 ), .B2(n1249), .C1(
        \unit_decode/n1471 ), .C2(n1252), .A(\unit_decode/n3299 ), .ZN(
        \unit_decode/n3296 ) );
  AOI22_X1 U4895 ( .A1(n1255), .A2(\unit_decode/n4043 ), .B1(n1259), .B2(
        \unit_decode/n3939 ), .ZN(\unit_decode/n3299 ) );
  OAI221_X1 U4896 ( .B1(\unit_decode/n1400 ), .B2(n1202), .C1(
        \unit_decode/n1377 ), .C2(n1205), .A(\unit_decode/n3273 ), .ZN(
        \unit_decode/n3270 ) );
  AOI22_X1 U4897 ( .A1(n1208), .A2(\unit_decode/n4041 ), .B1(n1211), .B2(
        \unit_decode/n3753 ), .ZN(\unit_decode/n3273 ) );
  OAI221_X1 U4898 ( .B1(\unit_decode/n1496 ), .B2(n1250), .C1(
        \unit_decode/n1472 ), .C2(n1253), .A(\unit_decode/n3281 ), .ZN(
        \unit_decode/n3278 ) );
  AOI22_X1 U4899 ( .A1(n1256), .A2(\unit_decode/n4039 ), .B1(n1259), .B2(
        \unit_decode/n3933 ), .ZN(\unit_decode/n3281 ) );
  OAI221_X1 U4900 ( .B1(\unit_decode/n1401 ), .B2(n1202), .C1(
        \unit_decode/n1378 ), .C2(n1205), .A(\unit_decode/n3255 ), .ZN(
        \unit_decode/n3252 ) );
  AOI22_X1 U4901 ( .A1(n1208), .A2(\unit_decode/n4037 ), .B1(n1211), .B2(
        \unit_decode/n3747 ), .ZN(\unit_decode/n3255 ) );
  OAI221_X1 U4902 ( .B1(\unit_decode/n1497 ), .B2(n1250), .C1(
        \unit_decode/n1473 ), .C2(n1253), .A(\unit_decode/n3263 ), .ZN(
        \unit_decode/n3260 ) );
  AOI22_X1 U4903 ( .A1(n1256), .A2(\unit_decode/n4035 ), .B1(n1259), .B2(
        \unit_decode/n3927 ), .ZN(\unit_decode/n3263 ) );
  OAI221_X1 U4904 ( .B1(\unit_decode/n1402 ), .B2(n1202), .C1(
        \unit_decode/n1379 ), .C2(n1205), .A(\unit_decode/n3237 ), .ZN(
        \unit_decode/n3234 ) );
  AOI22_X1 U4905 ( .A1(n1208), .A2(\unit_decode/n4033 ), .B1(n1211), .B2(
        \unit_decode/n3741 ), .ZN(\unit_decode/n3237 ) );
  OAI221_X1 U4906 ( .B1(\unit_decode/n1498 ), .B2(n1250), .C1(
        \unit_decode/n1474 ), .C2(n1253), .A(\unit_decode/n3245 ), .ZN(
        \unit_decode/n3242 ) );
  AOI22_X1 U4907 ( .A1(n1256), .A2(\unit_decode/n4031 ), .B1(n1259), .B2(
        \unit_decode/n3921 ), .ZN(\unit_decode/n3245 ) );
  OAI221_X1 U4908 ( .B1(\unit_decode/n1403 ), .B2(n1202), .C1(
        \unit_decode/n1380 ), .C2(n1205), .A(\unit_decode/n3219 ), .ZN(
        \unit_decode/n3216 ) );
  AOI22_X1 U4909 ( .A1(n1208), .A2(\unit_decode/n4029 ), .B1(n1211), .B2(
        \unit_decode/n3735 ), .ZN(\unit_decode/n3219 ) );
  OAI221_X1 U4910 ( .B1(\unit_decode/n1499 ), .B2(n1250), .C1(
        \unit_decode/n1475 ), .C2(n1253), .A(\unit_decode/n3227 ), .ZN(
        \unit_decode/n3224 ) );
  AOI22_X1 U4911 ( .A1(n1256), .A2(\unit_decode/n4027 ), .B1(n1259), .B2(
        \unit_decode/n3915 ), .ZN(\unit_decode/n3227 ) );
  OAI221_X1 U4912 ( .B1(\unit_decode/n1404 ), .B2(n1202), .C1(
        \unit_decode/n1381 ), .C2(n1205), .A(\unit_decode/n3201 ), .ZN(
        \unit_decode/n3198 ) );
  AOI22_X1 U4913 ( .A1(n1208), .A2(\unit_decode/n4025 ), .B1(n1211), .B2(
        \unit_decode/n3729 ), .ZN(\unit_decode/n3201 ) );
  OAI221_X1 U4914 ( .B1(\unit_decode/n1500 ), .B2(n1250), .C1(
        \unit_decode/n1476 ), .C2(n1253), .A(\unit_decode/n3209 ), .ZN(
        \unit_decode/n3206 ) );
  AOI22_X1 U4915 ( .A1(n1256), .A2(\unit_decode/n4023 ), .B1(n1259), .B2(
        \unit_decode/n3909 ), .ZN(\unit_decode/n3209 ) );
  OAI221_X1 U4916 ( .B1(\unit_decode/n1405 ), .B2(n1202), .C1(
        \unit_decode/n1382 ), .C2(n1205), .A(\unit_decode/n3183 ), .ZN(
        \unit_decode/n3180 ) );
  AOI22_X1 U4917 ( .A1(n1208), .A2(\unit_decode/n4021 ), .B1(n1211), .B2(
        \unit_decode/n3723 ), .ZN(\unit_decode/n3183 ) );
  OAI221_X1 U4918 ( .B1(\unit_decode/n1501 ), .B2(n1250), .C1(
        \unit_decode/n1477 ), .C2(n1253), .A(\unit_decode/n3191 ), .ZN(
        \unit_decode/n3188 ) );
  AOI22_X1 U4919 ( .A1(n1256), .A2(\unit_decode/n4019 ), .B1(n1259), .B2(
        \unit_decode/n3903 ), .ZN(\unit_decode/n3191 ) );
  OAI221_X1 U4920 ( .B1(\unit_decode/n1406 ), .B2(n1202), .C1(
        \unit_decode/n1383 ), .C2(n1205), .A(\unit_decode/n3165 ), .ZN(
        \unit_decode/n3162 ) );
  AOI22_X1 U4921 ( .A1(n1208), .A2(\unit_decode/n4137 ), .B1(n1211), .B2(
        \unit_decode/n3717 ), .ZN(\unit_decode/n3165 ) );
  OAI221_X1 U4922 ( .B1(\unit_decode/n1502 ), .B2(n1250), .C1(
        \unit_decode/n1478 ), .C2(n1253), .A(\unit_decode/n3173 ), .ZN(
        \unit_decode/n3170 ) );
  AOI22_X1 U4923 ( .A1(n1256), .A2(\unit_decode/n4135 ), .B1(n1259), .B2(
        \unit_decode/n3897 ), .ZN(\unit_decode/n3173 ) );
  OAI221_X1 U4924 ( .B1(\unit_decode/n1407 ), .B2(n1202), .C1(
        \unit_decode/n1384 ), .C2(n1205), .A(\unit_decode/n3147 ), .ZN(
        \unit_decode/n3144 ) );
  AOI22_X1 U4925 ( .A1(n1208), .A2(\unit_decode/n4133 ), .B1(n1211), .B2(
        \unit_decode/n3711 ), .ZN(\unit_decode/n3147 ) );
  OAI221_X1 U4926 ( .B1(\unit_decode/n1503 ), .B2(n1250), .C1(
        \unit_decode/n1479 ), .C2(n1253), .A(\unit_decode/n3155 ), .ZN(
        \unit_decode/n3152 ) );
  AOI22_X1 U4927 ( .A1(n1256), .A2(\unit_decode/n4131 ), .B1(n1259), .B2(
        \unit_decode/n3891 ), .ZN(\unit_decode/n3155 ) );
  OAI221_X1 U4928 ( .B1(\unit_decode/n1408 ), .B2(n1202), .C1(
        \unit_decode/n1385 ), .C2(n1205), .A(\unit_decode/n3129 ), .ZN(
        \unit_decode/n3126 ) );
  AOI22_X1 U4929 ( .A1(n1208), .A2(\unit_decode/n4129 ), .B1(n1210), .B2(
        \unit_decode/n3705 ), .ZN(\unit_decode/n3129 ) );
  OAI221_X1 U4930 ( .B1(\unit_decode/n1504 ), .B2(n1250), .C1(
        \unit_decode/n1480 ), .C2(n1253), .A(\unit_decode/n3137 ), .ZN(
        \unit_decode/n3134 ) );
  AOI22_X1 U4931 ( .A1(n1256), .A2(\unit_decode/n4127 ), .B1(n1258), .B2(
        \unit_decode/n3885 ), .ZN(\unit_decode/n3137 ) );
  OAI221_X1 U4932 ( .B1(\unit_decode/n1409 ), .B2(n1202), .C1(
        \unit_decode/n1386 ), .C2(n1205), .A(\unit_decode/n3111 ), .ZN(
        \unit_decode/n3108 ) );
  AOI22_X1 U4933 ( .A1(n1208), .A2(\unit_decode/n4125 ), .B1(n1210), .B2(
        \unit_decode/n3699 ), .ZN(\unit_decode/n3111 ) );
  OAI221_X1 U4934 ( .B1(\unit_decode/n1505 ), .B2(n1250), .C1(
        \unit_decode/n1481 ), .C2(n1253), .A(\unit_decode/n3119 ), .ZN(
        \unit_decode/n3116 ) );
  AOI22_X1 U4935 ( .A1(n1256), .A2(\unit_decode/n4123 ), .B1(n1258), .B2(
        \unit_decode/n3879 ), .ZN(\unit_decode/n3119 ) );
  OAI221_X1 U4936 ( .B1(\unit_decode/n1410 ), .B2(n1202), .C1(
        \unit_decode/n1387 ), .C2(n1205), .A(\unit_decode/n3093 ), .ZN(
        \unit_decode/n3090 ) );
  AOI22_X1 U4937 ( .A1(n1208), .A2(\unit_decode/n4121 ), .B1(n1210), .B2(
        \unit_decode/n3693 ), .ZN(\unit_decode/n3093 ) );
  OAI221_X1 U4938 ( .B1(\unit_decode/n1506 ), .B2(n1250), .C1(
        \unit_decode/n1482 ), .C2(n1253), .A(\unit_decode/n3101 ), .ZN(
        \unit_decode/n3098 ) );
  AOI22_X1 U4939 ( .A1(n1256), .A2(\unit_decode/n4119 ), .B1(n1258), .B2(
        \unit_decode/n3873 ), .ZN(\unit_decode/n3101 ) );
  OAI221_X1 U4940 ( .B1(\unit_decode/n1411 ), .B2(n1202), .C1(
        \unit_decode/n2084 ), .C2(n1205), .A(\unit_decode/n3075 ), .ZN(
        \unit_decode/n3072 ) );
  AOI22_X1 U4941 ( .A1(n1208), .A2(\unit_decode/n4117 ), .B1(n1210), .B2(
        \unit_decode/n3687 ), .ZN(\unit_decode/n3075 ) );
  OAI221_X1 U4942 ( .B1(\unit_decode/n1507 ), .B2(n1250), .C1(
        \unit_decode/n1483 ), .C2(n1253), .A(\unit_decode/n3083 ), .ZN(
        \unit_decode/n3080 ) );
  AOI22_X1 U4943 ( .A1(n1256), .A2(\unit_decode/n4115 ), .B1(n1258), .B2(
        \unit_decode/n3867 ), .ZN(\unit_decode/n3083 ) );
  OAI221_X1 U4944 ( .B1(\unit_decode/RegisterFile/n3707 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3739 ), .C2(n1120), .A(\unit_decode/n2876 ), 
        .ZN(\unit_decode/n2865 ) );
  AOI22_X1 U4945 ( .A1(n1123), .A2(\unit_decode/n2011 ), .B1(n1128), .B2(
        \unit_decode/n1987 ), .ZN(\unit_decode/n2876 ) );
  OAI221_X1 U4946 ( .B1(\unit_decode/RegisterFile/n3706 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3738 ), .C2(n1120), .A(\unit_decode/n2852 ), 
        .ZN(\unit_decode/n2847 ) );
  AOI22_X1 U4947 ( .A1(n1123), .A2(\unit_decode/n2010 ), .B1(n1128), .B2(
        \unit_decode/n1986 ), .ZN(\unit_decode/n2852 ) );
  OAI221_X1 U4948 ( .B1(\unit_decode/RegisterFile/n3705 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3737 ), .C2(n1120), .A(\unit_decode/n2834 ), 
        .ZN(\unit_decode/n2829 ) );
  AOI22_X1 U4949 ( .A1(n1123), .A2(\unit_decode/n2009 ), .B1(n1128), .B2(
        \unit_decode/n1985 ), .ZN(\unit_decode/n2834 ) );
  OAI221_X1 U4950 ( .B1(\unit_decode/RegisterFile/n3704 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3736 ), .C2(n1120), .A(\unit_decode/n2816 ), 
        .ZN(\unit_decode/n2811 ) );
  AOI22_X1 U4951 ( .A1(n1123), .A2(\unit_decode/n2008 ), .B1(n1128), .B2(
        \unit_decode/n1984 ), .ZN(\unit_decode/n2816 ) );
  OAI221_X1 U4952 ( .B1(\unit_decode/RegisterFile/n3703 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3735 ), .C2(n1120), .A(\unit_decode/n2798 ), 
        .ZN(\unit_decode/n2793 ) );
  AOI22_X1 U4953 ( .A1(n1123), .A2(\unit_decode/n2007 ), .B1(n1128), .B2(
        \unit_decode/n1983 ), .ZN(\unit_decode/n2798 ) );
  OAI221_X1 U4954 ( .B1(\unit_decode/RegisterFile/n3702 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3734 ), .C2(n1120), .A(\unit_decode/n2780 ), 
        .ZN(\unit_decode/n2775 ) );
  AOI22_X1 U4955 ( .A1(n1123), .A2(\unit_decode/n2006 ), .B1(n1128), .B2(
        \unit_decode/n1982 ), .ZN(\unit_decode/n2780 ) );
  OAI221_X1 U4956 ( .B1(\unit_decode/RegisterFile/n3701 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3733 ), .C2(n1120), .A(\unit_decode/n2762 ), 
        .ZN(\unit_decode/n2757 ) );
  AOI22_X1 U4957 ( .A1(n1123), .A2(\unit_decode/n2005 ), .B1(n1128), .B2(
        \unit_decode/n1981 ), .ZN(\unit_decode/n2762 ) );
  OAI221_X1 U4958 ( .B1(\unit_decode/RegisterFile/n3700 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3732 ), .C2(n1120), .A(\unit_decode/n2744 ), 
        .ZN(\unit_decode/n2739 ) );
  AOI22_X1 U4959 ( .A1(n1123), .A2(\unit_decode/n2004 ), .B1(n1128), .B2(
        \unit_decode/n1980 ), .ZN(\unit_decode/n2744 ) );
  OAI221_X1 U4960 ( .B1(\unit_decode/RegisterFile/n3699 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3731 ), .C2(n1120), .A(\unit_decode/n2726 ), 
        .ZN(\unit_decode/n2721 ) );
  AOI22_X1 U4961 ( .A1(n1123), .A2(\unit_decode/n2003 ), .B1(n1127), .B2(
        \unit_decode/n1979 ), .ZN(\unit_decode/n2726 ) );
  OAI221_X1 U4962 ( .B1(\unit_decode/RegisterFile/n3698 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3730 ), .C2(n1120), .A(\unit_decode/n2708 ), 
        .ZN(\unit_decode/n2703 ) );
  AOI22_X1 U4963 ( .A1(n1123), .A2(\unit_decode/n2002 ), .B1(n1127), .B2(
        \unit_decode/n1978 ), .ZN(\unit_decode/n2708 ) );
  OAI221_X1 U4964 ( .B1(\unit_decode/RegisterFile/n3697 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3729 ), .C2(n1120), .A(\unit_decode/n2690 ), 
        .ZN(\unit_decode/n2685 ) );
  AOI22_X1 U4965 ( .A1(n1123), .A2(\unit_decode/n2001 ), .B1(n1127), .B2(
        \unit_decode/n1977 ), .ZN(\unit_decode/n2690 ) );
  OAI221_X1 U4966 ( .B1(\unit_decode/RegisterFile/n3696 ), .B2(n1117), .C1(
        \unit_decode/RegisterFile/n3728 ), .C2(n1120), .A(\unit_decode/n2672 ), 
        .ZN(\unit_decode/n2667 ) );
  AOI22_X1 U4967 ( .A1(n1123), .A2(\unit_decode/n2000 ), .B1(n1127), .B2(
        \unit_decode/n1976 ), .ZN(\unit_decode/n2672 ) );
  OAI221_X1 U4968 ( .B1(\unit_decode/RegisterFile/n3695 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3727 ), .C2(n1121), .A(\unit_decode/n2654 ), 
        .ZN(\unit_decode/n2649 ) );
  AOI22_X1 U4969 ( .A1(n1124), .A2(\unit_decode/n1999 ), .B1(n1127), .B2(
        \unit_decode/n1975 ), .ZN(\unit_decode/n2654 ) );
  OAI221_X1 U4970 ( .B1(\unit_decode/RegisterFile/n3694 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3726 ), .C2(n1121), .A(\unit_decode/n2636 ), 
        .ZN(\unit_decode/n2631 ) );
  AOI22_X1 U4971 ( .A1(n1124), .A2(\unit_decode/n1998 ), .B1(n1127), .B2(
        \unit_decode/n1974 ), .ZN(\unit_decode/n2636 ) );
  OAI221_X1 U4972 ( .B1(\unit_decode/RegisterFile/n3693 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3725 ), .C2(n1121), .A(\unit_decode/n2618 ), 
        .ZN(\unit_decode/n2613 ) );
  AOI22_X1 U4973 ( .A1(n1124), .A2(\unit_decode/n1997 ), .B1(n1127), .B2(
        \unit_decode/n1973 ), .ZN(\unit_decode/n2618 ) );
  OAI221_X1 U4974 ( .B1(\unit_decode/RegisterFile/n3692 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3724 ), .C2(n1121), .A(\unit_decode/n2600 ), 
        .ZN(\unit_decode/n2595 ) );
  AOI22_X1 U4975 ( .A1(n1124), .A2(\unit_decode/n1996 ), .B1(n1127), .B2(
        \unit_decode/n1972 ), .ZN(\unit_decode/n2600 ) );
  OAI221_X1 U4976 ( .B1(\unit_decode/RegisterFile/n3691 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3723 ), .C2(n1121), .A(\unit_decode/n2582 ), 
        .ZN(\unit_decode/n2577 ) );
  AOI22_X1 U4977 ( .A1(n1124), .A2(\unit_decode/n1995 ), .B1(n1127), .B2(
        \unit_decode/n1971 ), .ZN(\unit_decode/n2582 ) );
  OAI221_X1 U4978 ( .B1(\unit_decode/RegisterFile/n3690 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3722 ), .C2(n1121), .A(\unit_decode/n2564 ), 
        .ZN(\unit_decode/n2559 ) );
  AOI22_X1 U4979 ( .A1(n1124), .A2(\unit_decode/n1994 ), .B1(n1127), .B2(
        \unit_decode/n1970 ), .ZN(\unit_decode/n2564 ) );
  OAI221_X1 U4980 ( .B1(\unit_decode/RegisterFile/n3689 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3721 ), .C2(n1121), .A(\unit_decode/n2546 ), 
        .ZN(\unit_decode/n2541 ) );
  AOI22_X1 U4981 ( .A1(n1124), .A2(\unit_decode/n1993 ), .B1(n1127), .B2(
        \unit_decode/n1969 ), .ZN(\unit_decode/n2546 ) );
  OAI221_X1 U4982 ( .B1(\unit_decode/RegisterFile/n3688 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3720 ), .C2(n1121), .A(\unit_decode/n2528 ), 
        .ZN(\unit_decode/n2523 ) );
  AOI22_X1 U4983 ( .A1(n1124), .A2(\unit_decode/n1992 ), .B1(n1127), .B2(
        \unit_decode/n1968 ), .ZN(\unit_decode/n2528 ) );
  OAI221_X1 U4984 ( .B1(\unit_decode/RegisterFile/n3687 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3719 ), .C2(n1121), .A(\unit_decode/n2510 ), 
        .ZN(\unit_decode/n2505 ) );
  AOI22_X1 U4985 ( .A1(n1124), .A2(\unit_decode/n1991 ), .B1(n1126), .B2(
        \unit_decode/n1967 ), .ZN(\unit_decode/n2510 ) );
  OAI221_X1 U4986 ( .B1(\unit_decode/RegisterFile/n3686 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3718 ), .C2(n1121), .A(\unit_decode/n2492 ), 
        .ZN(\unit_decode/n2487 ) );
  AOI22_X1 U4987 ( .A1(n1124), .A2(\unit_decode/n1990 ), .B1(n1126), .B2(
        \unit_decode/n1966 ), .ZN(\unit_decode/n2492 ) );
  OAI221_X1 U4988 ( .B1(\unit_decode/RegisterFile/n3685 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3717 ), .C2(n1121), .A(\unit_decode/n2474 ), 
        .ZN(\unit_decode/n2469 ) );
  AOI22_X1 U4989 ( .A1(n1124), .A2(\unit_decode/n1989 ), .B1(n1126), .B2(
        \unit_decode/n1965 ), .ZN(\unit_decode/n2474 ) );
  OAI221_X1 U4990 ( .B1(\unit_decode/RegisterFile/n3684 ), .B2(n1118), .C1(
        \unit_decode/RegisterFile/n3716 ), .C2(n1121), .A(\unit_decode/n2456 ), 
        .ZN(\unit_decode/n2451 ) );
  AOI22_X1 U4991 ( .A1(n1124), .A2(\unit_decode/n1988 ), .B1(n1126), .B2(
        \unit_decode/n1964 ), .ZN(\unit_decode/n2456 ) );
  OAI221_X1 U4992 ( .B1(\unit_decode/RegisterFile/n3683 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3715 ), .C2(n1122), .A(\unit_decode/n2438 ), 
        .ZN(\unit_decode/n2433 ) );
  AOI22_X1 U4993 ( .A1(n1125), .A2(\unit_decode/n1763 ), .B1(n1126), .B2(
        \unit_decode/n1755 ), .ZN(\unit_decode/n2438 ) );
  OAI221_X1 U4994 ( .B1(\unit_decode/RegisterFile/n3682 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3714 ), .C2(n1122), .A(\unit_decode/n2420 ), 
        .ZN(\unit_decode/n2415 ) );
  AOI22_X1 U4995 ( .A1(n1125), .A2(\unit_decode/n1762 ), .B1(n1126), .B2(
        \unit_decode/n1754 ), .ZN(\unit_decode/n2420 ) );
  OAI221_X1 U4996 ( .B1(\unit_decode/RegisterFile/n3681 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3713 ), .C2(n1122), .A(\unit_decode/n2402 ), 
        .ZN(\unit_decode/n2397 ) );
  AOI22_X1 U4997 ( .A1(n1125), .A2(\unit_decode/n1761 ), .B1(n1126), .B2(
        \unit_decode/n1753 ), .ZN(\unit_decode/n2402 ) );
  OAI221_X1 U4998 ( .B1(\unit_decode/RegisterFile/n3680 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3712 ), .C2(n1122), .A(\unit_decode/n2384 ), 
        .ZN(\unit_decode/n2379 ) );
  AOI22_X1 U4999 ( .A1(n1125), .A2(\unit_decode/n1760 ), .B1(n1126), .B2(
        \unit_decode/n1752 ), .ZN(\unit_decode/n2384 ) );
  OAI221_X1 U5000 ( .B1(\unit_decode/RegisterFile/n3679 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3711 ), .C2(n1122), .A(\unit_decode/n2366 ), 
        .ZN(\unit_decode/n2361 ) );
  AOI22_X1 U5001 ( .A1(n1125), .A2(\unit_decode/n1759 ), .B1(n1126), .B2(
        \unit_decode/n1751 ), .ZN(\unit_decode/n2366 ) );
  OAI221_X1 U5002 ( .B1(\unit_decode/RegisterFile/n3678 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3710 ), .C2(n1122), .A(\unit_decode/n2348 ), 
        .ZN(\unit_decode/n2343 ) );
  AOI22_X1 U5003 ( .A1(n1125), .A2(\unit_decode/n1758 ), .B1(n1126), .B2(
        \unit_decode/n1750 ), .ZN(\unit_decode/n2348 ) );
  OAI221_X1 U5004 ( .B1(\unit_decode/RegisterFile/n3677 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3709 ), .C2(n1122), .A(\unit_decode/n2330 ), 
        .ZN(\unit_decode/n2325 ) );
  AOI22_X1 U5005 ( .A1(n1125), .A2(\unit_decode/n1757 ), .B1(n1126), .B2(
        \unit_decode/n1749 ), .ZN(\unit_decode/n2330 ) );
  OAI221_X1 U5006 ( .B1(\unit_decode/RegisterFile/n3676 ), .B2(n1119), .C1(
        \unit_decode/RegisterFile/n3708 ), .C2(n1122), .A(\unit_decode/n2290 ), 
        .ZN(\unit_decode/n2275 ) );
  AOI22_X1 U5007 ( .A1(n1125), .A2(\unit_decode/n1756 ), .B1(n1126), .B2(
        \unit_decode/n1748 ), .ZN(\unit_decode/n2290 ) );
  OAI221_X1 U5008 ( .B1(\unit_decode/RegisterFile/n3707 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3739 ), .C2(n1216), .A(\unit_decode/n3496 ), 
        .ZN(\unit_decode/n3485 ) );
  AOI22_X1 U5009 ( .A1(n1219), .A2(\unit_decode/n2011 ), .B1(n1224), .B2(
        \unit_decode/n1987 ), .ZN(\unit_decode/n3496 ) );
  OAI221_X1 U5010 ( .B1(\unit_decode/RegisterFile/n3706 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3738 ), .C2(n1216), .A(\unit_decode/n3472 ), 
        .ZN(\unit_decode/n3467 ) );
  AOI22_X1 U5011 ( .A1(n1219), .A2(\unit_decode/n2010 ), .B1(n1224), .B2(
        \unit_decode/n1986 ), .ZN(\unit_decode/n3472 ) );
  OAI221_X1 U5012 ( .B1(\unit_decode/RegisterFile/n3705 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3737 ), .C2(n1216), .A(\unit_decode/n3454 ), 
        .ZN(\unit_decode/n3449 ) );
  AOI22_X1 U5013 ( .A1(n1219), .A2(\unit_decode/n2009 ), .B1(n1224), .B2(
        \unit_decode/n1985 ), .ZN(\unit_decode/n3454 ) );
  OAI221_X1 U5014 ( .B1(\unit_decode/RegisterFile/n3704 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3736 ), .C2(n1216), .A(\unit_decode/n3436 ), 
        .ZN(\unit_decode/n3431 ) );
  AOI22_X1 U5015 ( .A1(n1219), .A2(\unit_decode/n2008 ), .B1(n1224), .B2(
        \unit_decode/n1984 ), .ZN(\unit_decode/n3436 ) );
  OAI221_X1 U5016 ( .B1(\unit_decode/RegisterFile/n3703 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3735 ), .C2(n1216), .A(\unit_decode/n3418 ), 
        .ZN(\unit_decode/n3413 ) );
  AOI22_X1 U5017 ( .A1(n1219), .A2(\unit_decode/n2007 ), .B1(n1224), .B2(
        \unit_decode/n1983 ), .ZN(\unit_decode/n3418 ) );
  OAI221_X1 U5018 ( .B1(\unit_decode/RegisterFile/n3702 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3734 ), .C2(n1216), .A(\unit_decode/n3400 ), 
        .ZN(\unit_decode/n3395 ) );
  AOI22_X1 U5019 ( .A1(n1219), .A2(\unit_decode/n2006 ), .B1(n1224), .B2(
        \unit_decode/n1982 ), .ZN(\unit_decode/n3400 ) );
  OAI221_X1 U5020 ( .B1(\unit_decode/RegisterFile/n3701 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3733 ), .C2(n1216), .A(\unit_decode/n3382 ), 
        .ZN(\unit_decode/n3377 ) );
  AOI22_X1 U5021 ( .A1(n1219), .A2(\unit_decode/n2005 ), .B1(n1224), .B2(
        \unit_decode/n1981 ), .ZN(\unit_decode/n3382 ) );
  OAI221_X1 U5022 ( .B1(\unit_decode/RegisterFile/n3700 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3732 ), .C2(n1216), .A(\unit_decode/n3364 ), 
        .ZN(\unit_decode/n3359 ) );
  AOI22_X1 U5023 ( .A1(n1219), .A2(\unit_decode/n2004 ), .B1(n1224), .B2(
        \unit_decode/n1980 ), .ZN(\unit_decode/n3364 ) );
  OAI221_X1 U5024 ( .B1(\unit_decode/RegisterFile/n3699 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3731 ), .C2(n1216), .A(\unit_decode/n3346 ), 
        .ZN(\unit_decode/n3341 ) );
  AOI22_X1 U5025 ( .A1(n1219), .A2(\unit_decode/n2003 ), .B1(n1223), .B2(
        \unit_decode/n1979 ), .ZN(\unit_decode/n3346 ) );
  OAI221_X1 U5026 ( .B1(\unit_decode/RegisterFile/n3698 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3730 ), .C2(n1216), .A(\unit_decode/n3328 ), 
        .ZN(\unit_decode/n3323 ) );
  AOI22_X1 U5027 ( .A1(n1219), .A2(\unit_decode/n2002 ), .B1(n1223), .B2(
        \unit_decode/n1978 ), .ZN(\unit_decode/n3328 ) );
  OAI221_X1 U5028 ( .B1(\unit_decode/RegisterFile/n3697 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3729 ), .C2(n1216), .A(\unit_decode/n3310 ), 
        .ZN(\unit_decode/n3305 ) );
  AOI22_X1 U5029 ( .A1(n1219), .A2(\unit_decode/n2001 ), .B1(n1223), .B2(
        \unit_decode/n1977 ), .ZN(\unit_decode/n3310 ) );
  OAI221_X1 U5030 ( .B1(\unit_decode/RegisterFile/n3696 ), .B2(n1213), .C1(
        \unit_decode/RegisterFile/n3728 ), .C2(n1216), .A(\unit_decode/n3292 ), 
        .ZN(\unit_decode/n3287 ) );
  AOI22_X1 U5031 ( .A1(n1219), .A2(\unit_decode/n2000 ), .B1(n1223), .B2(
        \unit_decode/n1976 ), .ZN(\unit_decode/n3292 ) );
  OAI221_X1 U5032 ( .B1(\unit_decode/RegisterFile/n3695 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3727 ), .C2(n1217), .A(\unit_decode/n3274 ), 
        .ZN(\unit_decode/n3269 ) );
  AOI22_X1 U5033 ( .A1(n1220), .A2(\unit_decode/n1999 ), .B1(n1223), .B2(
        \unit_decode/n1975 ), .ZN(\unit_decode/n3274 ) );
  OAI221_X1 U5034 ( .B1(\unit_decode/RegisterFile/n3694 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3726 ), .C2(n1217), .A(\unit_decode/n3256 ), 
        .ZN(\unit_decode/n3251 ) );
  AOI22_X1 U5035 ( .A1(n1220), .A2(\unit_decode/n1998 ), .B1(n1223), .B2(
        \unit_decode/n1974 ), .ZN(\unit_decode/n3256 ) );
  OAI221_X1 U5036 ( .B1(\unit_decode/RegisterFile/n3693 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3725 ), .C2(n1217), .A(\unit_decode/n3238 ), 
        .ZN(\unit_decode/n3233 ) );
  AOI22_X1 U5037 ( .A1(n1220), .A2(\unit_decode/n1997 ), .B1(n1223), .B2(
        \unit_decode/n1973 ), .ZN(\unit_decode/n3238 ) );
  OAI221_X1 U5038 ( .B1(\unit_decode/RegisterFile/n3692 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3724 ), .C2(n1217), .A(\unit_decode/n3220 ), 
        .ZN(\unit_decode/n3215 ) );
  AOI22_X1 U5039 ( .A1(n1220), .A2(\unit_decode/n1996 ), .B1(n1223), .B2(
        \unit_decode/n1972 ), .ZN(\unit_decode/n3220 ) );
  OAI221_X1 U5040 ( .B1(\unit_decode/RegisterFile/n3691 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3723 ), .C2(n1217), .A(\unit_decode/n3202 ), 
        .ZN(\unit_decode/n3197 ) );
  AOI22_X1 U5041 ( .A1(n1220), .A2(\unit_decode/n1995 ), .B1(n1223), .B2(
        \unit_decode/n1971 ), .ZN(\unit_decode/n3202 ) );
  OAI221_X1 U5042 ( .B1(\unit_decode/RegisterFile/n3690 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3722 ), .C2(n1217), .A(\unit_decode/n3184 ), 
        .ZN(\unit_decode/n3179 ) );
  AOI22_X1 U5043 ( .A1(n1220), .A2(\unit_decode/n1994 ), .B1(n1223), .B2(
        \unit_decode/n1970 ), .ZN(\unit_decode/n3184 ) );
  OAI221_X1 U5044 ( .B1(\unit_decode/RegisterFile/n3689 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3721 ), .C2(n1217), .A(\unit_decode/n3166 ), 
        .ZN(\unit_decode/n3161 ) );
  AOI22_X1 U5045 ( .A1(n1220), .A2(\unit_decode/n1993 ), .B1(n1223), .B2(
        \unit_decode/n1969 ), .ZN(\unit_decode/n3166 ) );
  OAI221_X1 U5046 ( .B1(\unit_decode/RegisterFile/n3688 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3720 ), .C2(n1217), .A(\unit_decode/n3148 ), 
        .ZN(\unit_decode/n3143 ) );
  AOI22_X1 U5047 ( .A1(n1220), .A2(\unit_decode/n1992 ), .B1(n1223), .B2(
        \unit_decode/n1968 ), .ZN(\unit_decode/n3148 ) );
  OAI221_X1 U5048 ( .B1(\unit_decode/RegisterFile/n3687 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3719 ), .C2(n1217), .A(\unit_decode/n3130 ), 
        .ZN(\unit_decode/n3125 ) );
  AOI22_X1 U5049 ( .A1(n1220), .A2(\unit_decode/n1991 ), .B1(n1222), .B2(
        \unit_decode/n1967 ), .ZN(\unit_decode/n3130 ) );
  OAI221_X1 U5050 ( .B1(\unit_decode/RegisterFile/n3686 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3718 ), .C2(n1217), .A(\unit_decode/n3112 ), 
        .ZN(\unit_decode/n3107 ) );
  AOI22_X1 U5051 ( .A1(n1220), .A2(\unit_decode/n1990 ), .B1(n1222), .B2(
        \unit_decode/n1966 ), .ZN(\unit_decode/n3112 ) );
  OAI221_X1 U5052 ( .B1(\unit_decode/RegisterFile/n3685 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3717 ), .C2(n1217), .A(\unit_decode/n3094 ), 
        .ZN(\unit_decode/n3089 ) );
  AOI22_X1 U5053 ( .A1(n1220), .A2(\unit_decode/n1989 ), .B1(n1222), .B2(
        \unit_decode/n1965 ), .ZN(\unit_decode/n3094 ) );
  OAI221_X1 U5054 ( .B1(\unit_decode/RegisterFile/n3684 ), .B2(n1214), .C1(
        \unit_decode/RegisterFile/n3716 ), .C2(n1217), .A(\unit_decode/n3076 ), 
        .ZN(\unit_decode/n3071 ) );
  AOI22_X1 U5055 ( .A1(n1220), .A2(\unit_decode/n1988 ), .B1(n1222), .B2(
        \unit_decode/n1964 ), .ZN(\unit_decode/n3076 ) );
  OAI221_X1 U5056 ( .B1(\unit_decode/RegisterFile/n3683 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3715 ), .C2(n1218), .A(\unit_decode/n3058 ), 
        .ZN(\unit_decode/n3053 ) );
  AOI22_X1 U5057 ( .A1(n1221), .A2(\unit_decode/n1763 ), .B1(n1222), .B2(
        \unit_decode/n1755 ), .ZN(\unit_decode/n3058 ) );
  OAI221_X1 U5058 ( .B1(\unit_decode/RegisterFile/n3682 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3714 ), .C2(n1218), .A(\unit_decode/n3040 ), 
        .ZN(\unit_decode/n3035 ) );
  AOI22_X1 U5059 ( .A1(n1221), .A2(\unit_decode/n1762 ), .B1(n1222), .B2(
        \unit_decode/n1754 ), .ZN(\unit_decode/n3040 ) );
  OAI221_X1 U5060 ( .B1(\unit_decode/RegisterFile/n3681 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3713 ), .C2(n1218), .A(\unit_decode/n3022 ), 
        .ZN(\unit_decode/n3017 ) );
  AOI22_X1 U5061 ( .A1(n1221), .A2(\unit_decode/n1761 ), .B1(n1222), .B2(
        \unit_decode/n1753 ), .ZN(\unit_decode/n3022 ) );
  OAI221_X1 U5062 ( .B1(\unit_decode/RegisterFile/n3680 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3712 ), .C2(n1218), .A(\unit_decode/n3004 ), 
        .ZN(\unit_decode/n2999 ) );
  AOI22_X1 U5063 ( .A1(n1221), .A2(\unit_decode/n1760 ), .B1(n1222), .B2(
        \unit_decode/n1752 ), .ZN(\unit_decode/n3004 ) );
  OAI221_X1 U5064 ( .B1(\unit_decode/RegisterFile/n3679 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3711 ), .C2(n1218), .A(\unit_decode/n2986 ), 
        .ZN(\unit_decode/n2981 ) );
  AOI22_X1 U5065 ( .A1(n1221), .A2(\unit_decode/n1759 ), .B1(n1222), .B2(
        \unit_decode/n1751 ), .ZN(\unit_decode/n2986 ) );
  OAI221_X1 U5066 ( .B1(\unit_decode/RegisterFile/n3678 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3710 ), .C2(n1218), .A(\unit_decode/n2968 ), 
        .ZN(\unit_decode/n2963 ) );
  AOI22_X1 U5067 ( .A1(n1221), .A2(\unit_decode/n1758 ), .B1(n1222), .B2(
        \unit_decode/n1750 ), .ZN(\unit_decode/n2968 ) );
  OAI221_X1 U5068 ( .B1(\unit_decode/RegisterFile/n3677 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3709 ), .C2(n1218), .A(\unit_decode/n2950 ), 
        .ZN(\unit_decode/n2945 ) );
  AOI22_X1 U5069 ( .A1(n1221), .A2(\unit_decode/n1757 ), .B1(n1222), .B2(
        \unit_decode/n1749 ), .ZN(\unit_decode/n2950 ) );
  OAI221_X1 U5070 ( .B1(\unit_decode/RegisterFile/n3676 ), .B2(n1215), .C1(
        \unit_decode/RegisterFile/n3708 ), .C2(n1218), .A(\unit_decode/n2910 ), 
        .ZN(\unit_decode/n2895 ) );
  AOI22_X1 U5071 ( .A1(n1221), .A2(\unit_decode/n1756 ), .B1(n1222), .B2(
        \unit_decode/n1748 ), .ZN(\unit_decode/n2910 ) );
  OAI221_X1 U5072 ( .B1(\unit_decode/n1774 ), .B2(n1167), .C1(
        \unit_decode/RegisterFile/n3587 ), .C2(n1170), .A(\unit_decode/n2446 ), 
        .ZN(\unit_decode/n2441 ) );
  AOI22_X1 U5073 ( .A1(n1173), .A2(\unit_decode/RegisterFile/n8 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n40 ), .ZN(\unit_decode/n2446 ) );
  OAI221_X1 U5074 ( .B1(\unit_decode/n1773 ), .B2(n1167), .C1(
        \unit_decode/RegisterFile/n3586 ), .C2(n1170), .A(\unit_decode/n2428 ), 
        .ZN(\unit_decode/n2423 ) );
  AOI22_X1 U5075 ( .A1(n1173), .A2(\unit_decode/RegisterFile/n7 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n39 ), .ZN(\unit_decode/n2428 ) );
  OAI221_X1 U5076 ( .B1(\unit_decode/n1772 ), .B2(n1167), .C1(
        \unit_decode/RegisterFile/n3585 ), .C2(n1170), .A(\unit_decode/n2410 ), 
        .ZN(\unit_decode/n2405 ) );
  AOI22_X1 U5077 ( .A1(n1173), .A2(\unit_decode/RegisterFile/n6 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n38 ), .ZN(\unit_decode/n2410 ) );
  OAI221_X1 U5078 ( .B1(\unit_decode/n1771 ), .B2(n1167), .C1(
        \unit_decode/RegisterFile/n3584 ), .C2(n1170), .A(\unit_decode/n2392 ), 
        .ZN(\unit_decode/n2387 ) );
  AOI22_X1 U5079 ( .A1(n1173), .A2(\unit_decode/RegisterFile/n5 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n37 ), .ZN(\unit_decode/n2392 ) );
  OAI221_X1 U5080 ( .B1(\unit_decode/n1770 ), .B2(n1167), .C1(
        \unit_decode/RegisterFile/n3583 ), .C2(n1170), .A(\unit_decode/n2374 ), 
        .ZN(\unit_decode/n2369 ) );
  AOI22_X1 U5081 ( .A1(n1173), .A2(\unit_decode/RegisterFile/n4 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n36 ), .ZN(\unit_decode/n2374 ) );
  OAI221_X1 U5082 ( .B1(\unit_decode/n1774 ), .B2(n1263), .C1(
        \unit_decode/RegisterFile/n3587 ), .C2(n1266), .A(\unit_decode/n3066 ), 
        .ZN(\unit_decode/n3061 ) );
  AOI22_X1 U5083 ( .A1(n1269), .A2(\unit_decode/RegisterFile/n8 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n40 ), .ZN(\unit_decode/n3066 ) );
  OAI221_X1 U5084 ( .B1(\unit_decode/n1773 ), .B2(n1263), .C1(
        \unit_decode/RegisterFile/n3586 ), .C2(n1266), .A(\unit_decode/n3048 ), 
        .ZN(\unit_decode/n3043 ) );
  AOI22_X1 U5085 ( .A1(n1269), .A2(\unit_decode/RegisterFile/n7 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n39 ), .ZN(\unit_decode/n3048 ) );
  OAI221_X1 U5086 ( .B1(\unit_decode/n1772 ), .B2(n1263), .C1(
        \unit_decode/RegisterFile/n3585 ), .C2(n1266), .A(\unit_decode/n3030 ), 
        .ZN(\unit_decode/n3025 ) );
  AOI22_X1 U5087 ( .A1(n1269), .A2(\unit_decode/RegisterFile/n6 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n38 ), .ZN(\unit_decode/n3030 ) );
  OAI221_X1 U5088 ( .B1(\unit_decode/n1771 ), .B2(n1263), .C1(
        \unit_decode/RegisterFile/n3584 ), .C2(n1266), .A(\unit_decode/n3012 ), 
        .ZN(\unit_decode/n3007 ) );
  AOI22_X1 U5089 ( .A1(n1269), .A2(\unit_decode/RegisterFile/n5 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n37 ), .ZN(\unit_decode/n3012 ) );
  OAI221_X1 U5090 ( .B1(\unit_decode/n1770 ), .B2(n1263), .C1(
        \unit_decode/RegisterFile/n3583 ), .C2(n1266), .A(\unit_decode/n2994 ), 
        .ZN(\unit_decode/n2989 ) );
  AOI22_X1 U5091 ( .A1(n1269), .A2(\unit_decode/RegisterFile/n4 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n36 ), .ZN(\unit_decode/n2994 ) );
  OAI221_X1 U5092 ( .B1(\unit_decode/RegisterFile/n3870 ), .B2(n1131), .C1(
        \unit_decode/n1865 ), .C2(n1134), .A(\unit_decode/n2349 ), .ZN(
        \unit_decode/n2342 ) );
  AOI22_X1 U5093 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n451 ), .B1(n1138), .B2(\unit_decode/n3 ), .ZN(\unit_decode/n2349 ) );
  OAI221_X1 U5094 ( .B1(\unit_decode/RegisterFile/n3869 ), .B2(n1131), .C1(
        \unit_decode/n1864 ), .C2(n1134), .A(\unit_decode/n2331 ), .ZN(
        \unit_decode/n2324 ) );
  AOI22_X1 U5095 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n450 ), .B1(n1138), .B2(\unit_decode/n2 ), .ZN(\unit_decode/n2331 ) );
  OAI221_X1 U5096 ( .B1(\unit_decode/RegisterFile/n3868 ), .B2(n1131), .C1(
        \unit_decode/n1863 ), .C2(n1134), .A(\unit_decode/n2295 ), .ZN(
        \unit_decode/n2274 ) );
  AOI22_X1 U5097 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n449 ), .B1(n1138), .B2(\unit_decode/n1 ), .ZN(\unit_decode/n2295 ) );
  OAI221_X1 U5098 ( .B1(\unit_decode/RegisterFile/n3870 ), .B2(n1227), .C1(
        \unit_decode/n1865 ), .C2(n1230), .A(\unit_decode/n2969 ), .ZN(
        \unit_decode/n2962 ) );
  AOI22_X1 U5099 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n451 ), .B1(n1234), .B2(\unit_decode/n3 ), .ZN(\unit_decode/n2969 ) );
  OAI221_X1 U5100 ( .B1(\unit_decode/RegisterFile/n3869 ), .B2(n1227), .C1(
        \unit_decode/n1864 ), .C2(n1230), .A(\unit_decode/n2951 ), .ZN(
        \unit_decode/n2944 ) );
  AOI22_X1 U5101 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n450 ), .B1(n1234), .B2(\unit_decode/n2 ), .ZN(\unit_decode/n2951 ) );
  OAI221_X1 U5102 ( .B1(\unit_decode/RegisterFile/n3868 ), .B2(n1227), .C1(
        \unit_decode/n1863 ), .C2(n1230), .A(\unit_decode/n2915 ), .ZN(
        \unit_decode/n2894 ) );
  AOI22_X1 U5103 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n449 ), .B1(n1234), .B2(\unit_decode/n1 ), .ZN(\unit_decode/n2915 ) );
  OAI221_X1 U5104 ( .B1(\unit_decode/n1875 ), .B2(n1131), .C1(
        \unit_decode/n1870 ), .C2(n1134), .A(\unit_decode/n2439 ), .ZN(
        \unit_decode/n2432 ) );
  AOI22_X1 U5105 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n456 ), .B1(n1138), .B2(\unit_decode/n8 ), .ZN(\unit_decode/n2439 ) );
  OAI221_X1 U5106 ( .B1(\unit_decode/n1874 ), .B2(n1131), .C1(
        \unit_decode/n1869 ), .C2(n1134), .A(\unit_decode/n2421 ), .ZN(
        \unit_decode/n2414 ) );
  AOI22_X1 U5107 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n455 ), .B1(n1138), .B2(\unit_decode/n7 ), .ZN(\unit_decode/n2421 ) );
  OAI221_X1 U5108 ( .B1(\unit_decode/n1873 ), .B2(n1131), .C1(
        \unit_decode/n1868 ), .C2(n1134), .A(\unit_decode/n2403 ), .ZN(
        \unit_decode/n2396 ) );
  AOI22_X1 U5109 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n454 ), .B1(n1138), .B2(\unit_decode/n6 ), .ZN(\unit_decode/n2403 ) );
  OAI221_X1 U5110 ( .B1(\unit_decode/n1872 ), .B2(n1131), .C1(
        \unit_decode/n1867 ), .C2(n1134), .A(\unit_decode/n2385 ), .ZN(
        \unit_decode/n2378 ) );
  AOI22_X1 U5111 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n453 ), .B1(n1138), .B2(\unit_decode/n5 ), .ZN(\unit_decode/n2385 ) );
  OAI221_X1 U5112 ( .B1(\unit_decode/n1871 ), .B2(n1131), .C1(
        \unit_decode/n1866 ), .C2(n1134), .A(\unit_decode/n2367 ), .ZN(
        \unit_decode/n2360 ) );
  AOI22_X1 U5113 ( .A1(n1137), .A2(\unit_decode/RegisterFile/n452 ), .B1(n1138), .B2(\unit_decode/n4 ), .ZN(\unit_decode/n2367 ) );
  OAI221_X1 U5114 ( .B1(\unit_decode/n1875 ), .B2(n1227), .C1(
        \unit_decode/n1870 ), .C2(n1230), .A(\unit_decode/n3059 ), .ZN(
        \unit_decode/n3052 ) );
  AOI22_X1 U5115 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n456 ), .B1(n1234), .B2(\unit_decode/n8 ), .ZN(\unit_decode/n3059 ) );
  OAI221_X1 U5116 ( .B1(\unit_decode/n1874 ), .B2(n1227), .C1(
        \unit_decode/n1869 ), .C2(n1230), .A(\unit_decode/n3041 ), .ZN(
        \unit_decode/n3034 ) );
  AOI22_X1 U5117 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n455 ), .B1(n1234), .B2(\unit_decode/n7 ), .ZN(\unit_decode/n3041 ) );
  OAI221_X1 U5118 ( .B1(\unit_decode/n1873 ), .B2(n1227), .C1(
        \unit_decode/n1868 ), .C2(n1230), .A(\unit_decode/n3023 ), .ZN(
        \unit_decode/n3016 ) );
  AOI22_X1 U5119 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n454 ), .B1(n1234), .B2(\unit_decode/n6 ), .ZN(\unit_decode/n3023 ) );
  OAI221_X1 U5120 ( .B1(\unit_decode/n1872 ), .B2(n1227), .C1(
        \unit_decode/n1867 ), .C2(n1230), .A(\unit_decode/n3005 ), .ZN(
        \unit_decode/n2998 ) );
  AOI22_X1 U5121 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n453 ), .B1(n1234), .B2(\unit_decode/n5 ), .ZN(\unit_decode/n3005 ) );
  OAI221_X1 U5122 ( .B1(\unit_decode/n1871 ), .B2(n1227), .C1(
        \unit_decode/n1866 ), .C2(n1230), .A(\unit_decode/n2987 ), .ZN(
        \unit_decode/n2980 ) );
  AOI22_X1 U5123 ( .A1(n1233), .A2(\unit_decode/RegisterFile/n452 ), .B1(n1234), .B2(\unit_decode/n4 ), .ZN(\unit_decode/n2987 ) );
  OAI221_X1 U5124 ( .B1(\unit_memory/DRAM/n2615 ), .B2(n248), .C1(
        \unit_memory/DRAM/n2871 ), .C2(n235), .A(\unit_memory/DRAM/n2218 ), 
        .ZN(\unit_memory/DRAM/n2217 ) );
  AOI22_X1 U5125 ( .A1(n209), .A2(\unit_memory/DRAM/n249 ), .B1(n222), .B2(
        \unit_memory/DRAM/n505 ), .ZN(\unit_memory/DRAM/n2218 ) );
  OAI221_X1 U5126 ( .B1(\unit_memory/DRAM/n2497 ), .B2(n248), .C1(
        \unit_memory/DRAM/n2753 ), .C2(n235), .A(\unit_memory/DRAM/n873 ), 
        .ZN(\unit_memory/DRAM/n872 ) );
  AOI22_X1 U5127 ( .A1(n209), .A2(\unit_memory/DRAM/n131 ), .B1(n222), .B2(
        \unit_memory/DRAM/n387 ), .ZN(\unit_memory/DRAM/n873 ) );
  OAI221_X1 U5128 ( .B1(\unit_memory/DRAM/n2498 ), .B2(n248), .C1(
        \unit_memory/DRAM/n2754 ), .C2(n235), .A(\unit_memory/DRAM/n894 ), 
        .ZN(\unit_memory/DRAM/n893 ) );
  AOI22_X1 U5129 ( .A1(n209), .A2(\unit_memory/DRAM/n132 ), .B1(n222), .B2(
        \unit_memory/DRAM/n388 ), .ZN(\unit_memory/DRAM/n894 ) );
  OAI221_X1 U5130 ( .B1(\unit_decode/n2035 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3611 ), .C2(n1168), .A(\unit_decode/n2888 ), 
        .ZN(\unit_decode/n2881 ) );
  AOI22_X1 U5131 ( .A1(n1171), .A2(\unit_decode/n2083 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n64 ), .ZN(\unit_decode/n2888 ) );
  OAI221_X1 U5132 ( .B1(\unit_decode/n2034 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3610 ), .C2(n1168), .A(\unit_decode/n2860 ), 
        .ZN(\unit_decode/n2855 ) );
  AOI22_X1 U5133 ( .A1(n1171), .A2(\unit_decode/n2082 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n63 ), .ZN(\unit_decode/n2860 ) );
  OAI221_X1 U5134 ( .B1(\unit_decode/n2033 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3609 ), .C2(n1168), .A(\unit_decode/n2842 ), 
        .ZN(\unit_decode/n2837 ) );
  AOI22_X1 U5135 ( .A1(n1171), .A2(\unit_decode/n2081 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n62 ), .ZN(\unit_decode/n2842 ) );
  OAI221_X1 U5136 ( .B1(\unit_decode/n2032 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3608 ), .C2(n1168), .A(\unit_decode/n2824 ), 
        .ZN(\unit_decode/n2819 ) );
  AOI22_X1 U5137 ( .A1(n1171), .A2(\unit_decode/n2080 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n61 ), .ZN(\unit_decode/n2824 ) );
  OAI221_X1 U5138 ( .B1(\unit_decode/n2031 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3607 ), .C2(n1168), .A(\unit_decode/n2806 ), 
        .ZN(\unit_decode/n2801 ) );
  AOI22_X1 U5139 ( .A1(n1171), .A2(\unit_decode/n2079 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n60 ), .ZN(\unit_decode/n2806 ) );
  OAI221_X1 U5140 ( .B1(\unit_decode/n2030 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3606 ), .C2(n1168), .A(\unit_decode/n2788 ), 
        .ZN(\unit_decode/n2783 ) );
  AOI22_X1 U5141 ( .A1(n1171), .A2(\unit_decode/n2078 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n59 ), .ZN(\unit_decode/n2788 ) );
  OAI221_X1 U5142 ( .B1(\unit_decode/n2029 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3605 ), .C2(n1168), .A(\unit_decode/n2770 ), 
        .ZN(\unit_decode/n2765 ) );
  AOI22_X1 U5143 ( .A1(n1171), .A2(\unit_decode/n2077 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n58 ), .ZN(\unit_decode/n2770 ) );
  OAI221_X1 U5144 ( .B1(\unit_decode/n2028 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3604 ), .C2(n1168), .A(\unit_decode/n2752 ), 
        .ZN(\unit_decode/n2747 ) );
  AOI22_X1 U5145 ( .A1(n1171), .A2(\unit_decode/n2076 ), .B1(n1176), .B2(
        \unit_decode/RegisterFile/n57 ), .ZN(\unit_decode/n2752 ) );
  OAI221_X1 U5146 ( .B1(\unit_decode/n2027 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3603 ), .C2(n1168), .A(\unit_decode/n2734 ), 
        .ZN(\unit_decode/n2729 ) );
  AOI22_X1 U5147 ( .A1(n1171), .A2(\unit_decode/n2075 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n56 ), .ZN(\unit_decode/n2734 ) );
  OAI221_X1 U5148 ( .B1(\unit_decode/n2026 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3602 ), .C2(n1168), .A(\unit_decode/n2716 ), 
        .ZN(\unit_decode/n2711 ) );
  AOI22_X1 U5149 ( .A1(n1171), .A2(\unit_decode/n2074 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n55 ), .ZN(\unit_decode/n2716 ) );
  OAI221_X1 U5150 ( .B1(\unit_decode/n2025 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3601 ), .C2(n1168), .A(\unit_decode/n2698 ), 
        .ZN(\unit_decode/n2693 ) );
  AOI22_X1 U5151 ( .A1(n1171), .A2(\unit_decode/n2073 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n54 ), .ZN(\unit_decode/n2698 ) );
  OAI221_X1 U5152 ( .B1(\unit_decode/n2024 ), .B2(n1165), .C1(
        \unit_decode/RegisterFile/n3600 ), .C2(n1168), .A(\unit_decode/n2680 ), 
        .ZN(\unit_decode/n2675 ) );
  AOI22_X1 U5153 ( .A1(n1171), .A2(\unit_decode/n2072 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n53 ), .ZN(\unit_decode/n2680 ) );
  OAI221_X1 U5154 ( .B1(\unit_decode/n2023 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3599 ), .C2(n1169), .A(\unit_decode/n2662 ), 
        .ZN(\unit_decode/n2657 ) );
  AOI22_X1 U5155 ( .A1(n1172), .A2(\unit_decode/n2071 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n52 ), .ZN(\unit_decode/n2662 ) );
  OAI221_X1 U5156 ( .B1(\unit_decode/n2022 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3598 ), .C2(n1169), .A(\unit_decode/n2644 ), 
        .ZN(\unit_decode/n2639 ) );
  AOI22_X1 U5157 ( .A1(n1172), .A2(\unit_decode/n2070 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n51 ), .ZN(\unit_decode/n2644 ) );
  OAI221_X1 U5158 ( .B1(\unit_decode/n2021 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3597 ), .C2(n1169), .A(\unit_decode/n2626 ), 
        .ZN(\unit_decode/n2621 ) );
  AOI22_X1 U5159 ( .A1(n1172), .A2(\unit_decode/n2069 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n50 ), .ZN(\unit_decode/n2626 ) );
  OAI221_X1 U5160 ( .B1(\unit_decode/n2020 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3596 ), .C2(n1169), .A(\unit_decode/n2608 ), 
        .ZN(\unit_decode/n2603 ) );
  AOI22_X1 U5161 ( .A1(n1172), .A2(\unit_decode/n2068 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n49 ), .ZN(\unit_decode/n2608 ) );
  OAI221_X1 U5162 ( .B1(\unit_decode/n2019 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3595 ), .C2(n1169), .A(\unit_decode/n2590 ), 
        .ZN(\unit_decode/n2585 ) );
  AOI22_X1 U5163 ( .A1(n1172), .A2(\unit_decode/n2067 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n48 ), .ZN(\unit_decode/n2590 ) );
  OAI221_X1 U5164 ( .B1(\unit_decode/n2018 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3594 ), .C2(n1169), .A(\unit_decode/n2572 ), 
        .ZN(\unit_decode/n2567 ) );
  AOI22_X1 U5165 ( .A1(n1172), .A2(\unit_decode/n2066 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n47 ), .ZN(\unit_decode/n2572 ) );
  OAI221_X1 U5166 ( .B1(\unit_decode/n2017 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3593 ), .C2(n1169), .A(\unit_decode/n2554 ), 
        .ZN(\unit_decode/n2549 ) );
  AOI22_X1 U5167 ( .A1(n1172), .A2(\unit_decode/n2065 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n46 ), .ZN(\unit_decode/n2554 ) );
  OAI221_X1 U5168 ( .B1(\unit_decode/n2016 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3592 ), .C2(n1169), .A(\unit_decode/n2536 ), 
        .ZN(\unit_decode/n2531 ) );
  AOI22_X1 U5169 ( .A1(n1172), .A2(\unit_decode/n2064 ), .B1(n1175), .B2(
        \unit_decode/RegisterFile/n45 ), .ZN(\unit_decode/n2536 ) );
  OAI221_X1 U5170 ( .B1(\unit_decode/n2015 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3591 ), .C2(n1169), .A(\unit_decode/n2518 ), 
        .ZN(\unit_decode/n2513 ) );
  AOI22_X1 U5171 ( .A1(n1172), .A2(\unit_decode/n2063 ), .B1(n1174), .B2(
        \unit_decode/RegisterFile/n44 ), .ZN(\unit_decode/n2518 ) );
  OAI221_X1 U5172 ( .B1(\unit_decode/n2014 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3590 ), .C2(n1169), .A(\unit_decode/n2500 ), 
        .ZN(\unit_decode/n2495 ) );
  AOI22_X1 U5173 ( .A1(n1172), .A2(\unit_decode/n2062 ), .B1(n1174), .B2(
        \unit_decode/RegisterFile/n43 ), .ZN(\unit_decode/n2500 ) );
  OAI221_X1 U5174 ( .B1(\unit_decode/n2013 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3589 ), .C2(n1169), .A(\unit_decode/n2482 ), 
        .ZN(\unit_decode/n2477 ) );
  AOI22_X1 U5175 ( .A1(n1172), .A2(\unit_decode/n2061 ), .B1(n1174), .B2(
        \unit_decode/RegisterFile/n42 ), .ZN(\unit_decode/n2482 ) );
  OAI221_X1 U5176 ( .B1(\unit_decode/n2012 ), .B2(n1166), .C1(
        \unit_decode/RegisterFile/n3588 ), .C2(n1169), .A(\unit_decode/n2464 ), 
        .ZN(\unit_decode/n2459 ) );
  AOI22_X1 U5177 ( .A1(n1172), .A2(\unit_decode/RegisterFile/n9 ), .B1(n1174), 
        .B2(\unit_decode/RegisterFile/n41 ), .ZN(\unit_decode/n2464 ) );
  OAI221_X1 U5178 ( .B1(\unit_decode/n2035 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3611 ), .C2(n1264), .A(\unit_decode/n3508 ), 
        .ZN(\unit_decode/n3501 ) );
  AOI22_X1 U5179 ( .A1(n1267), .A2(\unit_decode/n2083 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n64 ), .ZN(\unit_decode/n3508 ) );
  OAI221_X1 U5180 ( .B1(\unit_decode/n2034 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3610 ), .C2(n1264), .A(\unit_decode/n3480 ), 
        .ZN(\unit_decode/n3475 ) );
  AOI22_X1 U5181 ( .A1(n1267), .A2(\unit_decode/n2082 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n63 ), .ZN(\unit_decode/n3480 ) );
  OAI221_X1 U5182 ( .B1(\unit_decode/n2033 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3609 ), .C2(n1264), .A(\unit_decode/n3462 ), 
        .ZN(\unit_decode/n3457 ) );
  AOI22_X1 U5183 ( .A1(n1267), .A2(\unit_decode/n2081 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n62 ), .ZN(\unit_decode/n3462 ) );
  OAI221_X1 U5184 ( .B1(\unit_decode/n2032 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3608 ), .C2(n1264), .A(\unit_decode/n3444 ), 
        .ZN(\unit_decode/n3439 ) );
  AOI22_X1 U5185 ( .A1(n1267), .A2(\unit_decode/n2080 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n61 ), .ZN(\unit_decode/n3444 ) );
  OAI221_X1 U5186 ( .B1(\unit_decode/n2031 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3607 ), .C2(n1264), .A(\unit_decode/n3426 ), 
        .ZN(\unit_decode/n3421 ) );
  AOI22_X1 U5187 ( .A1(n1267), .A2(\unit_decode/n2079 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n60 ), .ZN(\unit_decode/n3426 ) );
  OAI221_X1 U5188 ( .B1(\unit_decode/n2030 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3606 ), .C2(n1264), .A(\unit_decode/n3408 ), 
        .ZN(\unit_decode/n3403 ) );
  AOI22_X1 U5189 ( .A1(n1267), .A2(\unit_decode/n2078 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n59 ), .ZN(\unit_decode/n3408 ) );
  OAI221_X1 U5190 ( .B1(\unit_decode/n2029 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3605 ), .C2(n1264), .A(\unit_decode/n3390 ), 
        .ZN(\unit_decode/n3385 ) );
  AOI22_X1 U5191 ( .A1(n1267), .A2(\unit_decode/n2077 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n58 ), .ZN(\unit_decode/n3390 ) );
  OAI221_X1 U5192 ( .B1(\unit_decode/n2028 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3604 ), .C2(n1264), .A(\unit_decode/n3372 ), 
        .ZN(\unit_decode/n3367 ) );
  AOI22_X1 U5193 ( .A1(n1267), .A2(\unit_decode/n2076 ), .B1(n1272), .B2(
        \unit_decode/RegisterFile/n57 ), .ZN(\unit_decode/n3372 ) );
  OAI221_X1 U5194 ( .B1(\unit_decode/n2027 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3603 ), .C2(n1264), .A(\unit_decode/n3354 ), 
        .ZN(\unit_decode/n3349 ) );
  AOI22_X1 U5195 ( .A1(n1267), .A2(\unit_decode/n2075 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n56 ), .ZN(\unit_decode/n3354 ) );
  OAI221_X1 U5196 ( .B1(\unit_decode/n2026 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3602 ), .C2(n1264), .A(\unit_decode/n3336 ), 
        .ZN(\unit_decode/n3331 ) );
  AOI22_X1 U5197 ( .A1(n1267), .A2(\unit_decode/n2074 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n55 ), .ZN(\unit_decode/n3336 ) );
  OAI221_X1 U5198 ( .B1(\unit_decode/n2025 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3601 ), .C2(n1264), .A(\unit_decode/n3318 ), 
        .ZN(\unit_decode/n3313 ) );
  AOI22_X1 U5199 ( .A1(n1267), .A2(\unit_decode/n2073 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n54 ), .ZN(\unit_decode/n3318 ) );
  OAI221_X1 U5200 ( .B1(\unit_decode/n2024 ), .B2(n1261), .C1(
        \unit_decode/RegisterFile/n3600 ), .C2(n1264), .A(\unit_decode/n3300 ), 
        .ZN(\unit_decode/n3295 ) );
  AOI22_X1 U5201 ( .A1(n1267), .A2(\unit_decode/n2072 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n53 ), .ZN(\unit_decode/n3300 ) );
  OAI221_X1 U5202 ( .B1(\unit_decode/n2023 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3599 ), .C2(n1265), .A(\unit_decode/n3282 ), 
        .ZN(\unit_decode/n3277 ) );
  AOI22_X1 U5203 ( .A1(n1268), .A2(\unit_decode/n2071 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n52 ), .ZN(\unit_decode/n3282 ) );
  OAI221_X1 U5204 ( .B1(\unit_decode/n2022 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3598 ), .C2(n1265), .A(\unit_decode/n3264 ), 
        .ZN(\unit_decode/n3259 ) );
  AOI22_X1 U5205 ( .A1(n1268), .A2(\unit_decode/n2070 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n51 ), .ZN(\unit_decode/n3264 ) );
  OAI221_X1 U5206 ( .B1(\unit_decode/n2021 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3597 ), .C2(n1265), .A(\unit_decode/n3246 ), 
        .ZN(\unit_decode/n3241 ) );
  AOI22_X1 U5207 ( .A1(n1268), .A2(\unit_decode/n2069 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n50 ), .ZN(\unit_decode/n3246 ) );
  OAI221_X1 U5208 ( .B1(\unit_decode/n2020 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3596 ), .C2(n1265), .A(\unit_decode/n3228 ), 
        .ZN(\unit_decode/n3223 ) );
  AOI22_X1 U5209 ( .A1(n1268), .A2(\unit_decode/n2068 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n49 ), .ZN(\unit_decode/n3228 ) );
  OAI221_X1 U5210 ( .B1(\unit_decode/n2019 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3595 ), .C2(n1265), .A(\unit_decode/n3210 ), 
        .ZN(\unit_decode/n3205 ) );
  AOI22_X1 U5211 ( .A1(n1268), .A2(\unit_decode/n2067 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n48 ), .ZN(\unit_decode/n3210 ) );
  OAI221_X1 U5212 ( .B1(\unit_decode/n2018 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3594 ), .C2(n1265), .A(\unit_decode/n3192 ), 
        .ZN(\unit_decode/n3187 ) );
  AOI22_X1 U5213 ( .A1(n1268), .A2(\unit_decode/n2066 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n47 ), .ZN(\unit_decode/n3192 ) );
  OAI221_X1 U5214 ( .B1(\unit_decode/n2017 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3593 ), .C2(n1265), .A(\unit_decode/n3174 ), 
        .ZN(\unit_decode/n3169 ) );
  AOI22_X1 U5215 ( .A1(n1268), .A2(\unit_decode/n2065 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n46 ), .ZN(\unit_decode/n3174 ) );
  OAI221_X1 U5216 ( .B1(\unit_decode/n2016 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3592 ), .C2(n1265), .A(\unit_decode/n3156 ), 
        .ZN(\unit_decode/n3151 ) );
  AOI22_X1 U5217 ( .A1(n1268), .A2(\unit_decode/n2064 ), .B1(n1271), .B2(
        \unit_decode/RegisterFile/n45 ), .ZN(\unit_decode/n3156 ) );
  OAI221_X1 U5218 ( .B1(\unit_decode/n2015 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3591 ), .C2(n1265), .A(\unit_decode/n3138 ), 
        .ZN(\unit_decode/n3133 ) );
  AOI22_X1 U5219 ( .A1(n1268), .A2(\unit_decode/n2063 ), .B1(n1270), .B2(
        \unit_decode/RegisterFile/n44 ), .ZN(\unit_decode/n3138 ) );
  OAI221_X1 U5220 ( .B1(\unit_decode/n2014 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3590 ), .C2(n1265), .A(\unit_decode/n3120 ), 
        .ZN(\unit_decode/n3115 ) );
  AOI22_X1 U5221 ( .A1(n1268), .A2(\unit_decode/n2062 ), .B1(n1270), .B2(
        \unit_decode/RegisterFile/n43 ), .ZN(\unit_decode/n3120 ) );
  OAI221_X1 U5222 ( .B1(\unit_decode/n2013 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3589 ), .C2(n1265), .A(\unit_decode/n3102 ), 
        .ZN(\unit_decode/n3097 ) );
  AOI22_X1 U5223 ( .A1(n1268), .A2(\unit_decode/n2061 ), .B1(n1270), .B2(
        \unit_decode/RegisterFile/n42 ), .ZN(\unit_decode/n3102 ) );
  OAI221_X1 U5224 ( .B1(\unit_decode/n2012 ), .B2(n1262), .C1(
        \unit_decode/RegisterFile/n3588 ), .C2(n1265), .A(\unit_decode/n3084 ), 
        .ZN(\unit_decode/n3079 ) );
  AOI22_X1 U5225 ( .A1(n1268), .A2(\unit_decode/RegisterFile/n9 ), .B1(n1270), 
        .B2(\unit_decode/RegisterFile/n41 ), .ZN(\unit_decode/n3084 ) );
  OAI221_X1 U5226 ( .B1(\unit_decode/n1245 ), .B2(n1129), .C1(
        \unit_decode/n1221 ), .C2(n1132), .A(\unit_decode/n2878 ), .ZN(
        \unit_decode/n2864 ) );
  AOI22_X1 U5227 ( .A1(n1135), .A2(\unit_decode/n96 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n512 ), .ZN(\unit_decode/n2878 ) );
  OAI221_X1 U5228 ( .B1(\unit_decode/n1246 ), .B2(n1129), .C1(
        \unit_decode/n1222 ), .C2(n1132), .A(\unit_decode/n2853 ), .ZN(
        \unit_decode/n2846 ) );
  AOI22_X1 U5229 ( .A1(n1135), .A2(\unit_decode/n94 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n511 ), .ZN(\unit_decode/n2853 ) );
  OAI221_X1 U5230 ( .B1(\unit_decode/n1247 ), .B2(n1129), .C1(
        \unit_decode/n1223 ), .C2(n1132), .A(\unit_decode/n2835 ), .ZN(
        \unit_decode/n2828 ) );
  AOI22_X1 U5231 ( .A1(n1135), .A2(\unit_decode/n92 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n510 ), .ZN(\unit_decode/n2835 ) );
  OAI221_X1 U5232 ( .B1(\unit_decode/n1248 ), .B2(n1129), .C1(
        \unit_decode/n1224 ), .C2(n1132), .A(\unit_decode/n2817 ), .ZN(
        \unit_decode/n2810 ) );
  AOI22_X1 U5233 ( .A1(n1135), .A2(\unit_decode/n90 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n509 ), .ZN(\unit_decode/n2817 ) );
  OAI221_X1 U5234 ( .B1(\unit_decode/n1249 ), .B2(n1129), .C1(
        \unit_decode/n1225 ), .C2(n1132), .A(\unit_decode/n2799 ), .ZN(
        \unit_decode/n2792 ) );
  AOI22_X1 U5235 ( .A1(n1135), .A2(\unit_decode/n88 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n508 ), .ZN(\unit_decode/n2799 ) );
  OAI221_X1 U5236 ( .B1(\unit_decode/n1250 ), .B2(n1129), .C1(
        \unit_decode/n1226 ), .C2(n1132), .A(\unit_decode/n2781 ), .ZN(
        \unit_decode/n2774 ) );
  AOI22_X1 U5237 ( .A1(n1135), .A2(\unit_decode/n86 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n507 ), .ZN(\unit_decode/n2781 ) );
  OAI221_X1 U5238 ( .B1(\unit_decode/n1251 ), .B2(n1129), .C1(
        \unit_decode/n1227 ), .C2(n1132), .A(\unit_decode/n2763 ), .ZN(
        \unit_decode/n2756 ) );
  AOI22_X1 U5239 ( .A1(n1135), .A2(\unit_decode/n84 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n506 ), .ZN(\unit_decode/n2763 ) );
  OAI221_X1 U5240 ( .B1(\unit_decode/n1252 ), .B2(n1129), .C1(
        \unit_decode/n1228 ), .C2(n1132), .A(\unit_decode/n2745 ), .ZN(
        \unit_decode/n2738 ) );
  AOI22_X1 U5241 ( .A1(n1135), .A2(\unit_decode/n82 ), .B1(n1140), .B2(
        \unit_decode/RegisterFile/n505 ), .ZN(\unit_decode/n2745 ) );
  OAI221_X1 U5242 ( .B1(\unit_decode/n1253 ), .B2(n1129), .C1(
        \unit_decode/n1229 ), .C2(n1132), .A(\unit_decode/n2727 ), .ZN(
        \unit_decode/n2720 ) );
  AOI22_X1 U5243 ( .A1(n1135), .A2(\unit_decode/n80 ), .B1(n1139), .B2(
        \unit_decode/n24 ), .ZN(\unit_decode/n2727 ) );
  OAI221_X1 U5244 ( .B1(\unit_decode/n1254 ), .B2(n1129), .C1(
        \unit_decode/n1230 ), .C2(n1132), .A(\unit_decode/n2709 ), .ZN(
        \unit_decode/n2702 ) );
  AOI22_X1 U5245 ( .A1(n1135), .A2(\unit_decode/n78 ), .B1(n1139), .B2(
        \unit_decode/n23 ), .ZN(\unit_decode/n2709 ) );
  OAI221_X1 U5246 ( .B1(\unit_decode/n1255 ), .B2(n1129), .C1(
        \unit_decode/n1231 ), .C2(n1132), .A(\unit_decode/n2691 ), .ZN(
        \unit_decode/n2684 ) );
  AOI22_X1 U5247 ( .A1(n1135), .A2(\unit_decode/n76 ), .B1(n1139), .B2(
        \unit_decode/n22 ), .ZN(\unit_decode/n2691 ) );
  OAI221_X1 U5248 ( .B1(\unit_decode/n1256 ), .B2(n1129), .C1(
        \unit_decode/n1232 ), .C2(n1132), .A(\unit_decode/n2673 ), .ZN(
        \unit_decode/n2666 ) );
  AOI22_X1 U5249 ( .A1(n1135), .A2(\unit_decode/n74 ), .B1(n1139), .B2(
        \unit_decode/n21 ), .ZN(\unit_decode/n2673 ) );
  OAI221_X1 U5250 ( .B1(\unit_decode/n1257 ), .B2(n1130), .C1(
        \unit_decode/n1233 ), .C2(n1133), .A(\unit_decode/n2655 ), .ZN(
        \unit_decode/n2648 ) );
  AOI22_X1 U5251 ( .A1(n1136), .A2(\unit_decode/n72 ), .B1(n1139), .B2(
        \unit_decode/n20 ), .ZN(\unit_decode/n2655 ) );
  OAI221_X1 U5252 ( .B1(\unit_decode/n1258 ), .B2(n1130), .C1(
        \unit_decode/n1234 ), .C2(n1133), .A(\unit_decode/n2637 ), .ZN(
        \unit_decode/n2630 ) );
  AOI22_X1 U5253 ( .A1(n1136), .A2(\unit_decode/n70 ), .B1(n1139), .B2(
        \unit_decode/n19 ), .ZN(\unit_decode/n2637 ) );
  OAI221_X1 U5254 ( .B1(\unit_decode/n1259 ), .B2(n1130), .C1(
        \unit_decode/n1235 ), .C2(n1133), .A(\unit_decode/n2619 ), .ZN(
        \unit_decode/n2612 ) );
  AOI22_X1 U5255 ( .A1(n1136), .A2(\unit_decode/n68 ), .B1(n1139), .B2(
        \unit_decode/n18 ), .ZN(\unit_decode/n2619 ) );
  OAI221_X1 U5256 ( .B1(\unit_decode/n1260 ), .B2(n1130), .C1(
        \unit_decode/n1236 ), .C2(n1133), .A(\unit_decode/n2601 ), .ZN(
        \unit_decode/n2594 ) );
  AOI22_X1 U5257 ( .A1(n1136), .A2(\unit_decode/n66 ), .B1(n1139), .B2(
        \unit_decode/n17 ), .ZN(\unit_decode/n2601 ) );
  OAI221_X1 U5258 ( .B1(\unit_decode/n1261 ), .B2(n1130), .C1(
        \unit_decode/n1237 ), .C2(n1133), .A(\unit_decode/n2583 ), .ZN(
        \unit_decode/n2576 ) );
  AOI22_X1 U5259 ( .A1(n1136), .A2(\unit_decode/n64 ), .B1(n1139), .B2(
        \unit_decode/n16 ), .ZN(\unit_decode/n2583 ) );
  OAI221_X1 U5260 ( .B1(\unit_decode/n1262 ), .B2(n1130), .C1(
        \unit_decode/n1238 ), .C2(n1133), .A(\unit_decode/n2565 ), .ZN(
        \unit_decode/n2558 ) );
  AOI22_X1 U5261 ( .A1(n1136), .A2(\unit_decode/n62 ), .B1(n1139), .B2(
        \unit_decode/n15 ), .ZN(\unit_decode/n2565 ) );
  OAI221_X1 U5262 ( .B1(\unit_decode/n1263 ), .B2(n1130), .C1(
        \unit_decode/n1239 ), .C2(n1133), .A(\unit_decode/n2547 ), .ZN(
        \unit_decode/n2540 ) );
  AOI22_X1 U5263 ( .A1(n1136), .A2(\unit_decode/n60 ), .B1(n1139), .B2(
        \unit_decode/n14 ), .ZN(\unit_decode/n2547 ) );
  OAI221_X1 U5264 ( .B1(\unit_decode/n1264 ), .B2(n1130), .C1(
        \unit_decode/n1240 ), .C2(n1133), .A(\unit_decode/n2529 ), .ZN(
        \unit_decode/n2522 ) );
  AOI22_X1 U5265 ( .A1(n1136), .A2(\unit_decode/n58 ), .B1(n1139), .B2(
        \unit_decode/n13 ), .ZN(\unit_decode/n2529 ) );
  OAI221_X1 U5266 ( .B1(\unit_decode/n1265 ), .B2(n1130), .C1(
        \unit_decode/n1241 ), .C2(n1133), .A(\unit_decode/n2511 ), .ZN(
        \unit_decode/n2504 ) );
  AOI22_X1 U5267 ( .A1(n1136), .A2(\unit_decode/n56 ), .B1(n1138), .B2(
        \unit_decode/n12 ), .ZN(\unit_decode/n2511 ) );
  OAI221_X1 U5268 ( .B1(\unit_decode/n1266 ), .B2(n1130), .C1(
        \unit_decode/n1242 ), .C2(n1133), .A(\unit_decode/n2493 ), .ZN(
        \unit_decode/n2486 ) );
  AOI22_X1 U5269 ( .A1(n1136), .A2(\unit_decode/n54 ), .B1(n1138), .B2(
        \unit_decode/n11 ), .ZN(\unit_decode/n2493 ) );
  OAI221_X1 U5270 ( .B1(\unit_decode/n1267 ), .B2(n1130), .C1(
        \unit_decode/n1243 ), .C2(n1133), .A(\unit_decode/n2475 ), .ZN(
        \unit_decode/n2468 ) );
  AOI22_X1 U5271 ( .A1(n1136), .A2(\unit_decode/n52 ), .B1(n1138), .B2(
        \unit_decode/n10 ), .ZN(\unit_decode/n2475 ) );
  OAI221_X1 U5272 ( .B1(\unit_decode/n1268 ), .B2(n1130), .C1(
        \unit_decode/n1244 ), .C2(n1133), .A(\unit_decode/n2457 ), .ZN(
        \unit_decode/n2450 ) );
  AOI22_X1 U5273 ( .A1(n1136), .A2(\unit_decode/n50 ), .B1(n1138), .B2(
        \unit_decode/n9 ), .ZN(\unit_decode/n2457 ) );
  OAI221_X1 U5274 ( .B1(\unit_decode/n1245 ), .B2(n1225), .C1(
        \unit_decode/n1221 ), .C2(n1228), .A(\unit_decode/n3498 ), .ZN(
        \unit_decode/n3484 ) );
  AOI22_X1 U5275 ( .A1(n1231), .A2(\unit_decode/n96 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n512 ), .ZN(\unit_decode/n3498 ) );
  OAI221_X1 U5276 ( .B1(\unit_decode/n1246 ), .B2(n1225), .C1(
        \unit_decode/n1222 ), .C2(n1228), .A(\unit_decode/n3473 ), .ZN(
        \unit_decode/n3466 ) );
  AOI22_X1 U5277 ( .A1(n1231), .A2(\unit_decode/n94 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n511 ), .ZN(\unit_decode/n3473 ) );
  OAI221_X1 U5278 ( .B1(\unit_decode/n1247 ), .B2(n1225), .C1(
        \unit_decode/n1223 ), .C2(n1228), .A(\unit_decode/n3455 ), .ZN(
        \unit_decode/n3448 ) );
  AOI22_X1 U5279 ( .A1(n1231), .A2(\unit_decode/n92 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n510 ), .ZN(\unit_decode/n3455 ) );
  OAI221_X1 U5280 ( .B1(\unit_decode/n1248 ), .B2(n1225), .C1(
        \unit_decode/n1224 ), .C2(n1228), .A(\unit_decode/n3437 ), .ZN(
        \unit_decode/n3430 ) );
  AOI22_X1 U5281 ( .A1(n1231), .A2(\unit_decode/n90 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n509 ), .ZN(\unit_decode/n3437 ) );
  OAI221_X1 U5282 ( .B1(\unit_decode/n1249 ), .B2(n1225), .C1(
        \unit_decode/n1225 ), .C2(n1228), .A(\unit_decode/n3419 ), .ZN(
        \unit_decode/n3412 ) );
  AOI22_X1 U5283 ( .A1(n1231), .A2(\unit_decode/n88 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n508 ), .ZN(\unit_decode/n3419 ) );
  OAI221_X1 U5284 ( .B1(\unit_decode/n1250 ), .B2(n1225), .C1(
        \unit_decode/n1226 ), .C2(n1228), .A(\unit_decode/n3401 ), .ZN(
        \unit_decode/n3394 ) );
  AOI22_X1 U5285 ( .A1(n1231), .A2(\unit_decode/n86 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n507 ), .ZN(\unit_decode/n3401 ) );
  OAI221_X1 U5286 ( .B1(\unit_decode/n1251 ), .B2(n1225), .C1(
        \unit_decode/n1227 ), .C2(n1228), .A(\unit_decode/n3383 ), .ZN(
        \unit_decode/n3376 ) );
  AOI22_X1 U5287 ( .A1(n1231), .A2(\unit_decode/n84 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n506 ), .ZN(\unit_decode/n3383 ) );
  OAI221_X1 U5288 ( .B1(\unit_decode/n1252 ), .B2(n1225), .C1(
        \unit_decode/n1228 ), .C2(n1228), .A(\unit_decode/n3365 ), .ZN(
        \unit_decode/n3358 ) );
  AOI22_X1 U5289 ( .A1(n1231), .A2(\unit_decode/n82 ), .B1(n1236), .B2(
        \unit_decode/RegisterFile/n505 ), .ZN(\unit_decode/n3365 ) );
  OAI221_X1 U5290 ( .B1(\unit_decode/n1253 ), .B2(n1225), .C1(
        \unit_decode/n1229 ), .C2(n1228), .A(\unit_decode/n3347 ), .ZN(
        \unit_decode/n3340 ) );
  AOI22_X1 U5291 ( .A1(n1231), .A2(\unit_decode/n80 ), .B1(n1235), .B2(
        \unit_decode/n24 ), .ZN(\unit_decode/n3347 ) );
  OAI221_X1 U5292 ( .B1(\unit_decode/n1254 ), .B2(n1225), .C1(
        \unit_decode/n1230 ), .C2(n1228), .A(\unit_decode/n3329 ), .ZN(
        \unit_decode/n3322 ) );
  AOI22_X1 U5293 ( .A1(n1231), .A2(\unit_decode/n78 ), .B1(n1235), .B2(
        \unit_decode/n23 ), .ZN(\unit_decode/n3329 ) );
  OAI221_X1 U5294 ( .B1(\unit_decode/n1255 ), .B2(n1225), .C1(
        \unit_decode/n1231 ), .C2(n1228), .A(\unit_decode/n3311 ), .ZN(
        \unit_decode/n3304 ) );
  AOI22_X1 U5295 ( .A1(n1231), .A2(\unit_decode/n76 ), .B1(n1235), .B2(
        \unit_decode/n22 ), .ZN(\unit_decode/n3311 ) );
  OAI221_X1 U5296 ( .B1(\unit_decode/n1256 ), .B2(n1225), .C1(
        \unit_decode/n1232 ), .C2(n1228), .A(\unit_decode/n3293 ), .ZN(
        \unit_decode/n3286 ) );
  AOI22_X1 U5297 ( .A1(n1231), .A2(\unit_decode/n74 ), .B1(n1235), .B2(
        \unit_decode/n21 ), .ZN(\unit_decode/n3293 ) );
  OAI221_X1 U5298 ( .B1(\unit_decode/n1257 ), .B2(n1226), .C1(
        \unit_decode/n1233 ), .C2(n1229), .A(\unit_decode/n3275 ), .ZN(
        \unit_decode/n3268 ) );
  AOI22_X1 U5299 ( .A1(n1232), .A2(\unit_decode/n72 ), .B1(n1235), .B2(
        \unit_decode/n20 ), .ZN(\unit_decode/n3275 ) );
  OAI221_X1 U5300 ( .B1(\unit_decode/n1258 ), .B2(n1226), .C1(
        \unit_decode/n1234 ), .C2(n1229), .A(\unit_decode/n3257 ), .ZN(
        \unit_decode/n3250 ) );
  AOI22_X1 U5301 ( .A1(n1232), .A2(\unit_decode/n70 ), .B1(n1235), .B2(
        \unit_decode/n19 ), .ZN(\unit_decode/n3257 ) );
  OAI221_X1 U5302 ( .B1(\unit_decode/n1259 ), .B2(n1226), .C1(
        \unit_decode/n1235 ), .C2(n1229), .A(\unit_decode/n3239 ), .ZN(
        \unit_decode/n3232 ) );
  AOI22_X1 U5303 ( .A1(n1232), .A2(\unit_decode/n68 ), .B1(n1235), .B2(
        \unit_decode/n18 ), .ZN(\unit_decode/n3239 ) );
  OAI221_X1 U5304 ( .B1(\unit_decode/n1260 ), .B2(n1226), .C1(
        \unit_decode/n1236 ), .C2(n1229), .A(\unit_decode/n3221 ), .ZN(
        \unit_decode/n3214 ) );
  AOI22_X1 U5305 ( .A1(n1232), .A2(\unit_decode/n66 ), .B1(n1235), .B2(
        \unit_decode/n17 ), .ZN(\unit_decode/n3221 ) );
  OAI221_X1 U5306 ( .B1(\unit_decode/n1261 ), .B2(n1226), .C1(
        \unit_decode/n1237 ), .C2(n1229), .A(\unit_decode/n3203 ), .ZN(
        \unit_decode/n3196 ) );
  AOI22_X1 U5307 ( .A1(n1232), .A2(\unit_decode/n64 ), .B1(n1235), .B2(
        \unit_decode/n16 ), .ZN(\unit_decode/n3203 ) );
  OAI221_X1 U5308 ( .B1(\unit_decode/n1262 ), .B2(n1226), .C1(
        \unit_decode/n1238 ), .C2(n1229), .A(\unit_decode/n3185 ), .ZN(
        \unit_decode/n3178 ) );
  AOI22_X1 U5309 ( .A1(n1232), .A2(\unit_decode/n62 ), .B1(n1235), .B2(
        \unit_decode/n15 ), .ZN(\unit_decode/n3185 ) );
  OAI221_X1 U5310 ( .B1(\unit_decode/n1263 ), .B2(n1226), .C1(
        \unit_decode/n1239 ), .C2(n1229), .A(\unit_decode/n3167 ), .ZN(
        \unit_decode/n3160 ) );
  AOI22_X1 U5311 ( .A1(n1232), .A2(\unit_decode/n60 ), .B1(n1235), .B2(
        \unit_decode/n14 ), .ZN(\unit_decode/n3167 ) );
  OAI221_X1 U5312 ( .B1(\unit_decode/n1264 ), .B2(n1226), .C1(
        \unit_decode/n1240 ), .C2(n1229), .A(\unit_decode/n3149 ), .ZN(
        \unit_decode/n3142 ) );
  AOI22_X1 U5313 ( .A1(n1232), .A2(\unit_decode/n58 ), .B1(n1235), .B2(
        \unit_decode/n13 ), .ZN(\unit_decode/n3149 ) );
  OAI221_X1 U5314 ( .B1(\unit_decode/n1265 ), .B2(n1226), .C1(
        \unit_decode/n1241 ), .C2(n1229), .A(\unit_decode/n3131 ), .ZN(
        \unit_decode/n3124 ) );
  AOI22_X1 U5315 ( .A1(n1232), .A2(\unit_decode/n56 ), .B1(n1234), .B2(
        \unit_decode/n12 ), .ZN(\unit_decode/n3131 ) );
  OAI221_X1 U5316 ( .B1(\unit_decode/n1266 ), .B2(n1226), .C1(
        \unit_decode/n1242 ), .C2(n1229), .A(\unit_decode/n3113 ), .ZN(
        \unit_decode/n3106 ) );
  AOI22_X1 U5317 ( .A1(n1232), .A2(\unit_decode/n54 ), .B1(n1234), .B2(
        \unit_decode/n11 ), .ZN(\unit_decode/n3113 ) );
  OAI221_X1 U5318 ( .B1(\unit_decode/n1267 ), .B2(n1226), .C1(
        \unit_decode/n1243 ), .C2(n1229), .A(\unit_decode/n3095 ), .ZN(
        \unit_decode/n3088 ) );
  AOI22_X1 U5319 ( .A1(n1232), .A2(\unit_decode/n52 ), .B1(n1234), .B2(
        \unit_decode/n10 ), .ZN(\unit_decode/n3095 ) );
  OAI221_X1 U5320 ( .B1(\unit_decode/n1268 ), .B2(n1226), .C1(
        \unit_decode/n1244 ), .C2(n1229), .A(\unit_decode/n3077 ), .ZN(
        \unit_decode/n3070 ) );
  AOI22_X1 U5321 ( .A1(n1232), .A2(\unit_decode/n50 ), .B1(n1234), .B2(
        \unit_decode/n9 ), .ZN(\unit_decode/n3077 ) );
  OAI221_X1 U5322 ( .B1(\unit_memory/DRAM/n2543 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2799 ), .C2(n231), .A(\unit_memory/DRAM/n1149 ), 
        .ZN(\unit_memory/DRAM/n1147 ) );
  AOI22_X1 U5323 ( .A1(n205), .A2(\unit_memory/DRAM/n177 ), .B1(n218), .B2(
        \unit_memory/DRAM/n433 ), .ZN(\unit_memory/DRAM/n1149 ) );
  OAI221_X1 U5324 ( .B1(\unit_memory/DRAM/n2575 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2831 ), .C2(n233), .A(\unit_memory/DRAM/n1153 ), 
        .ZN(\unit_memory/DRAM/n1152 ) );
  AOI22_X1 U5325 ( .A1(n207), .A2(\unit_memory/DRAM/n209 ), .B1(n220), .B2(
        \unit_memory/DRAM/n465 ), .ZN(\unit_memory/DRAM/n1153 ) );
  OAI221_X1 U5326 ( .B1(\unit_memory/DRAM/n2607 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2863 ), .C2(n233), .A(\unit_memory/DRAM/n2181 ), 
        .ZN(\unit_memory/DRAM/n1156 ) );
  AOI22_X1 U5327 ( .A1(n207), .A2(\unit_memory/DRAM/n241 ), .B1(n220), .B2(
        \unit_memory/DRAM/n497 ), .ZN(\unit_memory/DRAM/n2181 ) );
  OAI221_X1 U5328 ( .B1(\unit_memory/DRAM/n2551 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2807 ), .C2(n234), .A(\unit_memory/DRAM/n2210 ), 
        .ZN(\unit_memory/DRAM/n2209 ) );
  AOI22_X1 U5329 ( .A1(n208), .A2(\unit_memory/DRAM/n185 ), .B1(n221), .B2(
        \unit_memory/DRAM/n441 ), .ZN(\unit_memory/DRAM/n2210 ) );
  OAI221_X1 U5330 ( .B1(\unit_memory/DRAM/n2495 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2751 ), .C2(n235), .A(\unit_memory/DRAM/n830 ), 
        .ZN(\unit_memory/DRAM/n828 ) );
  AOI22_X1 U5331 ( .A1(n209), .A2(\unit_memory/DRAM/n129 ), .B1(n222), .B2(
        \unit_memory/DRAM/n385 ), .ZN(\unit_memory/DRAM/n830 ) );
  OAI221_X1 U5332 ( .B1(\unit_memory/DRAM/n2527 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2783 ), .C2(n234), .A(\unit_memory/DRAM/n835 ), 
        .ZN(\unit_memory/DRAM/n833 ) );
  AOI22_X1 U5333 ( .A1(n208), .A2(\unit_memory/DRAM/n161 ), .B1(n221), .B2(
        \unit_memory/DRAM/n417 ), .ZN(\unit_memory/DRAM/n835 ) );
  OAI221_X1 U5334 ( .B1(\unit_memory/DRAM/n2496 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2752 ), .C2(n234), .A(\unit_memory/DRAM/n852 ), 
        .ZN(\unit_memory/DRAM/n851 ) );
  AOI22_X1 U5335 ( .A1(n208), .A2(\unit_memory/DRAM/n130 ), .B1(n221), .B2(
        \unit_memory/DRAM/n386 ), .ZN(\unit_memory/DRAM/n852 ) );
  OAI221_X1 U5336 ( .B1(\unit_memory/DRAM/n2528 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2784 ), .C2(n235), .A(\unit_memory/DRAM/n856 ), 
        .ZN(\unit_memory/DRAM/n855 ) );
  AOI22_X1 U5337 ( .A1(n209), .A2(\unit_memory/DRAM/n162 ), .B1(n222), .B2(
        \unit_memory/DRAM/n418 ), .ZN(\unit_memory/DRAM/n856 ) );
  OAI221_X1 U5338 ( .B1(\unit_memory/DRAM/n2529 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2785 ), .C2(n234), .A(\unit_memory/DRAM/n877 ), 
        .ZN(\unit_memory/DRAM/n876 ) );
  AOI22_X1 U5339 ( .A1(n208), .A2(\unit_memory/DRAM/n163 ), .B1(n221), .B2(
        \unit_memory/DRAM/n419 ), .ZN(\unit_memory/DRAM/n877 ) );
  OAI221_X1 U5340 ( .B1(\unit_memory/DRAM/n2530 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2786 ), .C2(n233), .A(\unit_memory/DRAM/n898 ), 
        .ZN(\unit_memory/DRAM/n897 ) );
  AOI22_X1 U5341 ( .A1(n207), .A2(\unit_memory/DRAM/n164 ), .B1(n220), .B2(
        \unit_memory/DRAM/n420 ), .ZN(\unit_memory/DRAM/n898 ) );
  OAI221_X1 U5342 ( .B1(\unit_memory/DRAM/n2499 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2755 ), .C2(n233), .A(\unit_memory/DRAM/n915 ), 
        .ZN(\unit_memory/DRAM/n914 ) );
  AOI22_X1 U5343 ( .A1(n207), .A2(\unit_memory/DRAM/n133 ), .B1(n220), .B2(
        \unit_memory/DRAM/n389 ), .ZN(\unit_memory/DRAM/n915 ) );
  OAI221_X1 U5344 ( .B1(\unit_memory/DRAM/n2531 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2787 ), .C2(n232), .A(\unit_memory/DRAM/n919 ), 
        .ZN(\unit_memory/DRAM/n918 ) );
  AOI22_X1 U5345 ( .A1(n206), .A2(\unit_memory/DRAM/n165 ), .B1(n219), .B2(
        \unit_memory/DRAM/n421 ), .ZN(\unit_memory/DRAM/n919 ) );
  OAI221_X1 U5346 ( .B1(\unit_memory/DRAM/n2500 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2756 ), .C2(n232), .A(\unit_memory/DRAM/n936 ), 
        .ZN(\unit_memory/DRAM/n935 ) );
  AOI22_X1 U5347 ( .A1(n206), .A2(\unit_memory/DRAM/n134 ), .B1(n219), .B2(
        \unit_memory/DRAM/n390 ), .ZN(\unit_memory/DRAM/n936 ) );
  OAI221_X1 U5348 ( .B1(\unit_memory/DRAM/n2532 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2788 ), .C2(n234), .A(\unit_memory/DRAM/n940 ), 
        .ZN(\unit_memory/DRAM/n939 ) );
  AOI22_X1 U5349 ( .A1(n208), .A2(\unit_memory/DRAM/n166 ), .B1(n221), .B2(
        \unit_memory/DRAM/n422 ), .ZN(\unit_memory/DRAM/n940 ) );
  OAI221_X1 U5350 ( .B1(\unit_memory/DRAM/n2501 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2757 ), .C2(n234), .A(\unit_memory/DRAM/n957 ), 
        .ZN(\unit_memory/DRAM/n956 ) );
  AOI22_X1 U5351 ( .A1(n208), .A2(\unit_memory/DRAM/n135 ), .B1(n221), .B2(
        \unit_memory/DRAM/n391 ), .ZN(\unit_memory/DRAM/n957 ) );
  OAI221_X1 U5352 ( .B1(\unit_memory/DRAM/n2533 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2789 ), .C2(n232), .A(\unit_memory/DRAM/n961 ), 
        .ZN(\unit_memory/DRAM/n960 ) );
  AOI22_X1 U5353 ( .A1(n206), .A2(\unit_memory/DRAM/n167 ), .B1(n219), .B2(
        \unit_memory/DRAM/n423 ), .ZN(\unit_memory/DRAM/n961 ) );
  OAI221_X1 U5354 ( .B1(\unit_memory/DRAM/n2502 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2758 ), .C2(n232), .A(\unit_memory/DRAM/n978 ), 
        .ZN(\unit_memory/DRAM/n977 ) );
  AOI22_X1 U5355 ( .A1(n206), .A2(\unit_memory/DRAM/n136 ), .B1(n219), .B2(
        \unit_memory/DRAM/n392 ), .ZN(\unit_memory/DRAM/n978 ) );
  OAI221_X1 U5356 ( .B1(\unit_memory/DRAM/n2534 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2790 ), .C2(n232), .A(\unit_memory/DRAM/n982 ), 
        .ZN(\unit_memory/DRAM/n981 ) );
  AOI22_X1 U5357 ( .A1(n206), .A2(\unit_memory/DRAM/n168 ), .B1(n219), .B2(
        \unit_memory/DRAM/n424 ), .ZN(\unit_memory/DRAM/n982 ) );
  OAI221_X1 U5358 ( .B1(\unit_memory/DRAM/n2503 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2759 ), .C2(n231), .A(\unit_memory/DRAM/n999 ), 
        .ZN(\unit_memory/DRAM/n998 ) );
  AOI22_X1 U5359 ( .A1(n205), .A2(\unit_memory/DRAM/n137 ), .B1(n218), .B2(
        \unit_memory/DRAM/n393 ), .ZN(\unit_memory/DRAM/n999 ) );
  OAI221_X1 U5360 ( .B1(\unit_memory/DRAM/n2535 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2791 ), .C2(n234), .A(\unit_memory/DRAM/n1003 ), 
        .ZN(\unit_memory/DRAM/n1002 ) );
  AOI22_X1 U5361 ( .A1(n208), .A2(\unit_memory/DRAM/n169 ), .B1(n221), .B2(
        \unit_memory/DRAM/n425 ), .ZN(\unit_memory/DRAM/n1003 ) );
  OAI221_X1 U5362 ( .B1(\unit_memory/DRAM/n2504 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2760 ), .C2(n233), .A(\unit_memory/DRAM/n1020 ), 
        .ZN(\unit_memory/DRAM/n1019 ) );
  AOI22_X1 U5363 ( .A1(n207), .A2(\unit_memory/DRAM/n138 ), .B1(n220), .B2(
        \unit_memory/DRAM/n394 ), .ZN(\unit_memory/DRAM/n1020 ) );
  OAI221_X1 U5364 ( .B1(\unit_memory/DRAM/n2536 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2792 ), .C2(n231), .A(\unit_memory/DRAM/n1024 ), 
        .ZN(\unit_memory/DRAM/n1023 ) );
  AOI22_X1 U5365 ( .A1(n205), .A2(\unit_memory/DRAM/n170 ), .B1(n218), .B2(
        \unit_memory/DRAM/n426 ), .ZN(\unit_memory/DRAM/n1024 ) );
  OAI221_X1 U5366 ( .B1(\unit_memory/DRAM/n2505 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2761 ), .C2(n232), .A(\unit_memory/DRAM/n1041 ), 
        .ZN(\unit_memory/DRAM/n1040 ) );
  AOI22_X1 U5367 ( .A1(n206), .A2(\unit_memory/DRAM/n139 ), .B1(n219), .B2(
        \unit_memory/DRAM/n395 ), .ZN(\unit_memory/DRAM/n1041 ) );
  OAI221_X1 U5368 ( .B1(\unit_memory/DRAM/n2537 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2793 ), .C2(n231), .A(\unit_memory/DRAM/n1045 ), 
        .ZN(\unit_memory/DRAM/n1044 ) );
  AOI22_X1 U5369 ( .A1(n205), .A2(\unit_memory/DRAM/n171 ), .B1(n218), .B2(
        \unit_memory/DRAM/n427 ), .ZN(\unit_memory/DRAM/n1045 ) );
  OAI221_X1 U5370 ( .B1(\unit_memory/DRAM/n2506 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2762 ), .C2(n231), .A(\unit_memory/DRAM/n1062 ), 
        .ZN(\unit_memory/DRAM/n1061 ) );
  AOI22_X1 U5371 ( .A1(n205), .A2(\unit_memory/DRAM/n140 ), .B1(n218), .B2(
        \unit_memory/DRAM/n396 ), .ZN(\unit_memory/DRAM/n1062 ) );
  OAI221_X1 U5372 ( .B1(\unit_memory/DRAM/n2538 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2794 ), .C2(n232), .A(\unit_memory/DRAM/n1066 ), 
        .ZN(\unit_memory/DRAM/n1065 ) );
  AOI22_X1 U5373 ( .A1(n206), .A2(\unit_memory/DRAM/n172 ), .B1(n219), .B2(
        \unit_memory/DRAM/n428 ), .ZN(\unit_memory/DRAM/n1066 ) );
  OAI221_X1 U5374 ( .B1(\unit_memory/DRAM/n2507 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2763 ), .C2(n232), .A(\unit_memory/DRAM/n1083 ), 
        .ZN(\unit_memory/DRAM/n1082 ) );
  AOI22_X1 U5375 ( .A1(n206), .A2(\unit_memory/DRAM/n141 ), .B1(n219), .B2(
        \unit_memory/DRAM/n397 ), .ZN(\unit_memory/DRAM/n1083 ) );
  OAI221_X1 U5376 ( .B1(\unit_memory/DRAM/n2539 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2795 ), .C2(n231), .A(\unit_memory/DRAM/n1087 ), 
        .ZN(\unit_memory/DRAM/n1086 ) );
  AOI22_X1 U5377 ( .A1(n205), .A2(\unit_memory/DRAM/n173 ), .B1(n218), .B2(
        \unit_memory/DRAM/n429 ), .ZN(\unit_memory/DRAM/n1087 ) );
  OAI221_X1 U5378 ( .B1(\unit_memory/DRAM/n2508 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2764 ), .C2(n231), .A(\unit_memory/DRAM/n1104 ), 
        .ZN(\unit_memory/DRAM/n1103 ) );
  AOI22_X1 U5379 ( .A1(n205), .A2(\unit_memory/DRAM/n142 ), .B1(n218), .B2(
        \unit_memory/DRAM/n398 ), .ZN(\unit_memory/DRAM/n1104 ) );
  OAI221_X1 U5380 ( .B1(\unit_memory/DRAM/n2540 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2796 ), .C2(n231), .A(\unit_memory/DRAM/n1108 ), 
        .ZN(\unit_memory/DRAM/n1107 ) );
  AOI22_X1 U5381 ( .A1(n205), .A2(\unit_memory/DRAM/n174 ), .B1(n218), .B2(
        \unit_memory/DRAM/n430 ), .ZN(\unit_memory/DRAM/n1108 ) );
  OAI221_X1 U5382 ( .B1(\unit_memory/DRAM/n2509 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2765 ), .C2(n233), .A(\unit_memory/DRAM/n1125 ), 
        .ZN(\unit_memory/DRAM/n1124 ) );
  AOI22_X1 U5383 ( .A1(n207), .A2(\unit_memory/DRAM/n143 ), .B1(n220), .B2(
        \unit_memory/DRAM/n399 ), .ZN(\unit_memory/DRAM/n1125 ) );
  OAI221_X1 U5384 ( .B1(\unit_memory/DRAM/n2541 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2797 ), .C2(n232), .A(\unit_memory/DRAM/n1129 ), 
        .ZN(\unit_memory/DRAM/n1128 ) );
  AOI22_X1 U5385 ( .A1(n206), .A2(\unit_memory/DRAM/n175 ), .B1(n219), .B2(
        \unit_memory/DRAM/n431 ), .ZN(\unit_memory/DRAM/n1129 ) );
  OAI221_X1 U5386 ( .B1(\unit_memory/DRAM/n2510 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2766 ), .C2(n233), .A(\unit_memory/DRAM/n2193 ), 
        .ZN(\unit_memory/DRAM/n2192 ) );
  AOI22_X1 U5387 ( .A1(n207), .A2(\unit_memory/DRAM/n144 ), .B1(n220), .B2(
        \unit_memory/DRAM/n400 ), .ZN(\unit_memory/DRAM/n2193 ) );
  OAI221_X1 U5388 ( .B1(\unit_memory/DRAM/n2542 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2798 ), .C2(n233), .A(\unit_memory/DRAM/n2197 ), 
        .ZN(\unit_memory/DRAM/n2196 ) );
  AOI22_X1 U5389 ( .A1(n207), .A2(\unit_memory/DRAM/n176 ), .B1(n220), .B2(
        \unit_memory/DRAM/n432 ), .ZN(\unit_memory/DRAM/n2197 ) );
  OAI221_X1 U5390 ( .B1(\unit_memory/DRAM/n2487 ), .B2(n196), .C1(
        \unit_memory/DRAM/n2743 ), .C2(n183), .A(\unit_memory/DRAM/n2219 ), 
        .ZN(\unit_memory/DRAM/n2216 ) );
  AOI22_X1 U5391 ( .A1(n157), .A2(\unit_memory/DRAM/n121 ), .B1(n170), .B2(
        \unit_memory/DRAM/n377 ), .ZN(\unit_memory/DRAM/n2219 ) );
  OAI221_X1 U5392 ( .B1(\unit_memory/DRAM/n2369 ), .B2(n196), .C1(
        \unit_memory/DRAM/n2625 ), .C2(n183), .A(\unit_memory/DRAM/n874 ), 
        .ZN(\unit_memory/DRAM/n871 ) );
  AOI22_X1 U5393 ( .A1(n157), .A2(\unit_memory/DRAM/n3 ), .B1(n170), .B2(
        \unit_memory/DRAM/n259 ), .ZN(\unit_memory/DRAM/n874 ) );
  OAI221_X1 U5394 ( .B1(\unit_memory/DRAM/n2370 ), .B2(n196), .C1(
        \unit_memory/DRAM/n2626 ), .C2(n183), .A(\unit_memory/DRAM/n895 ), 
        .ZN(\unit_memory/DRAM/n892 ) );
  AOI22_X1 U5395 ( .A1(n157), .A2(\unit_memory/DRAM/n4 ), .B1(n170), .B2(
        \unit_memory/DRAM/n260 ), .ZN(\unit_memory/DRAM/n895 ) );
  OAI221_X1 U5396 ( .B1(\unit_memory/DRAM/n2415 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2671 ), .C2(n179), .A(\unit_memory/DRAM/n1150 ), 
        .ZN(\unit_memory/DRAM/n1146 ) );
  AOI22_X1 U5397 ( .A1(n153), .A2(\unit_memory/DRAM/n49 ), .B1(n166), .B2(
        \unit_memory/DRAM/n305 ), .ZN(\unit_memory/DRAM/n1150 ) );
  OAI221_X1 U5398 ( .B1(\unit_memory/DRAM/n2447 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2703 ), .C2(n181), .A(\unit_memory/DRAM/n1154 ), 
        .ZN(\unit_memory/DRAM/n1151 ) );
  AOI22_X1 U5399 ( .A1(n155), .A2(\unit_memory/DRAM/n81 ), .B1(n168), .B2(
        \unit_memory/DRAM/n337 ), .ZN(\unit_memory/DRAM/n1154 ) );
  OAI221_X1 U5400 ( .B1(\unit_memory/DRAM/n2479 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2735 ), .C2(n181), .A(\unit_memory/DRAM/n2182 ), 
        .ZN(\unit_memory/DRAM/n1155 ) );
  AOI22_X1 U5401 ( .A1(n155), .A2(\unit_memory/DRAM/n113 ), .B1(n168), .B2(
        \unit_memory/DRAM/n369 ), .ZN(\unit_memory/DRAM/n2182 ) );
  OAI221_X1 U5402 ( .B1(\unit_memory/DRAM/n2423 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2679 ), .C2(n182), .A(\unit_memory/DRAM/n2211 ), 
        .ZN(\unit_memory/DRAM/n2208 ) );
  AOI22_X1 U5403 ( .A1(n156), .A2(\unit_memory/DRAM/n57 ), .B1(n169), .B2(
        \unit_memory/DRAM/n313 ), .ZN(\unit_memory/DRAM/n2211 ) );
  OAI221_X1 U5404 ( .B1(\unit_memory/DRAM/n2367 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2623 ), .C2(n183), .A(\unit_memory/DRAM/n831 ), 
        .ZN(\unit_memory/DRAM/n827 ) );
  AOI22_X1 U5405 ( .A1(n157), .A2(\unit_memory/DRAM/n1 ), .B1(n170), .B2(
        \unit_memory/DRAM/n257 ), .ZN(\unit_memory/DRAM/n831 ) );
  OAI221_X1 U5406 ( .B1(\unit_memory/DRAM/n2399 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2655 ), .C2(n182), .A(\unit_memory/DRAM/n836 ), 
        .ZN(\unit_memory/DRAM/n832 ) );
  AOI22_X1 U5407 ( .A1(n156), .A2(\unit_memory/DRAM/n33 ), .B1(n169), .B2(
        \unit_memory/DRAM/n289 ), .ZN(\unit_memory/DRAM/n836 ) );
  OAI221_X1 U5408 ( .B1(\unit_memory/DRAM/n2368 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2624 ), .C2(n182), .A(\unit_memory/DRAM/n853 ), 
        .ZN(\unit_memory/DRAM/n850 ) );
  AOI22_X1 U5409 ( .A1(n156), .A2(\unit_memory/DRAM/n2 ), .B1(n169), .B2(
        \unit_memory/DRAM/n258 ), .ZN(\unit_memory/DRAM/n853 ) );
  OAI221_X1 U5410 ( .B1(\unit_memory/DRAM/n2400 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2656 ), .C2(n183), .A(\unit_memory/DRAM/n857 ), 
        .ZN(\unit_memory/DRAM/n854 ) );
  AOI22_X1 U5411 ( .A1(n157), .A2(\unit_memory/DRAM/n34 ), .B1(n170), .B2(
        \unit_memory/DRAM/n290 ), .ZN(\unit_memory/DRAM/n857 ) );
  OAI221_X1 U5412 ( .B1(\unit_memory/DRAM/n2401 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2657 ), .C2(n182), .A(\unit_memory/DRAM/n878 ), 
        .ZN(\unit_memory/DRAM/n875 ) );
  AOI22_X1 U5413 ( .A1(n156), .A2(\unit_memory/DRAM/n35 ), .B1(n169), .B2(
        \unit_memory/DRAM/n291 ), .ZN(\unit_memory/DRAM/n878 ) );
  OAI221_X1 U5414 ( .B1(\unit_memory/DRAM/n2402 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2658 ), .C2(n181), .A(\unit_memory/DRAM/n899 ), 
        .ZN(\unit_memory/DRAM/n896 ) );
  AOI22_X1 U5415 ( .A1(n155), .A2(\unit_memory/DRAM/n36 ), .B1(n168), .B2(
        \unit_memory/DRAM/n292 ), .ZN(\unit_memory/DRAM/n899 ) );
  OAI221_X1 U5416 ( .B1(\unit_memory/DRAM/n2371 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2627 ), .C2(n181), .A(\unit_memory/DRAM/n916 ), 
        .ZN(\unit_memory/DRAM/n913 ) );
  AOI22_X1 U5417 ( .A1(n155), .A2(\unit_memory/DRAM/n5 ), .B1(n168), .B2(
        \unit_memory/DRAM/n261 ), .ZN(\unit_memory/DRAM/n916 ) );
  OAI221_X1 U5418 ( .B1(\unit_memory/DRAM/n2403 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2659 ), .C2(n180), .A(\unit_memory/DRAM/n920 ), 
        .ZN(\unit_memory/DRAM/n917 ) );
  AOI22_X1 U5419 ( .A1(n154), .A2(\unit_memory/DRAM/n37 ), .B1(n167), .B2(
        \unit_memory/DRAM/n293 ), .ZN(\unit_memory/DRAM/n920 ) );
  OAI221_X1 U5420 ( .B1(\unit_memory/DRAM/n2372 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2628 ), .C2(n180), .A(\unit_memory/DRAM/n937 ), 
        .ZN(\unit_memory/DRAM/n934 ) );
  AOI22_X1 U5421 ( .A1(n154), .A2(\unit_memory/DRAM/n6 ), .B1(n167), .B2(
        \unit_memory/DRAM/n262 ), .ZN(\unit_memory/DRAM/n937 ) );
  OAI221_X1 U5422 ( .B1(\unit_memory/DRAM/n2404 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2660 ), .C2(n182), .A(\unit_memory/DRAM/n941 ), 
        .ZN(\unit_memory/DRAM/n938 ) );
  AOI22_X1 U5423 ( .A1(n156), .A2(\unit_memory/DRAM/n38 ), .B1(n169), .B2(
        \unit_memory/DRAM/n294 ), .ZN(\unit_memory/DRAM/n941 ) );
  OAI221_X1 U5424 ( .B1(\unit_memory/DRAM/n2373 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2629 ), .C2(n182), .A(\unit_memory/DRAM/n958 ), 
        .ZN(\unit_memory/DRAM/n955 ) );
  AOI22_X1 U5425 ( .A1(n156), .A2(\unit_memory/DRAM/n7 ), .B1(n169), .B2(
        \unit_memory/DRAM/n263 ), .ZN(\unit_memory/DRAM/n958 ) );
  OAI221_X1 U5426 ( .B1(\unit_memory/DRAM/n2405 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2661 ), .C2(n180), .A(\unit_memory/DRAM/n962 ), 
        .ZN(\unit_memory/DRAM/n959 ) );
  AOI22_X1 U5427 ( .A1(n154), .A2(\unit_memory/DRAM/n39 ), .B1(n167), .B2(
        \unit_memory/DRAM/n295 ), .ZN(\unit_memory/DRAM/n962 ) );
  OAI221_X1 U5428 ( .B1(\unit_memory/DRAM/n2374 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2630 ), .C2(n180), .A(\unit_memory/DRAM/n979 ), 
        .ZN(\unit_memory/DRAM/n976 ) );
  AOI22_X1 U5429 ( .A1(n154), .A2(\unit_memory/DRAM/n8 ), .B1(n167), .B2(
        \unit_memory/DRAM/n264 ), .ZN(\unit_memory/DRAM/n979 ) );
  OAI221_X1 U5430 ( .B1(\unit_memory/DRAM/n2406 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2662 ), .C2(n180), .A(\unit_memory/DRAM/n983 ), 
        .ZN(\unit_memory/DRAM/n980 ) );
  AOI22_X1 U5431 ( .A1(n154), .A2(\unit_memory/DRAM/n40 ), .B1(n167), .B2(
        \unit_memory/DRAM/n296 ), .ZN(\unit_memory/DRAM/n983 ) );
  OAI221_X1 U5432 ( .B1(\unit_memory/DRAM/n2375 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2631 ), .C2(n179), .A(\unit_memory/DRAM/n1000 ), 
        .ZN(\unit_memory/DRAM/n997 ) );
  AOI22_X1 U5433 ( .A1(n153), .A2(\unit_memory/DRAM/n9 ), .B1(n166), .B2(
        \unit_memory/DRAM/n265 ), .ZN(\unit_memory/DRAM/n1000 ) );
  OAI221_X1 U5434 ( .B1(\unit_memory/DRAM/n2407 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2663 ), .C2(n182), .A(\unit_memory/DRAM/n1004 ), 
        .ZN(\unit_memory/DRAM/n1001 ) );
  AOI22_X1 U5435 ( .A1(n156), .A2(\unit_memory/DRAM/n41 ), .B1(n169), .B2(
        \unit_memory/DRAM/n297 ), .ZN(\unit_memory/DRAM/n1004 ) );
  OAI221_X1 U5436 ( .B1(\unit_memory/DRAM/n2376 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2632 ), .C2(n181), .A(\unit_memory/DRAM/n1021 ), 
        .ZN(\unit_memory/DRAM/n1018 ) );
  AOI22_X1 U5437 ( .A1(n155), .A2(\unit_memory/DRAM/n10 ), .B1(n168), .B2(
        \unit_memory/DRAM/n266 ), .ZN(\unit_memory/DRAM/n1021 ) );
  OAI221_X1 U5438 ( .B1(\unit_memory/DRAM/n2408 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2664 ), .C2(n179), .A(\unit_memory/DRAM/n1025 ), 
        .ZN(\unit_memory/DRAM/n1022 ) );
  AOI22_X1 U5439 ( .A1(n153), .A2(\unit_memory/DRAM/n42 ), .B1(n166), .B2(
        \unit_memory/DRAM/n298 ), .ZN(\unit_memory/DRAM/n1025 ) );
  OAI221_X1 U5440 ( .B1(\unit_memory/DRAM/n2377 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2633 ), .C2(n180), .A(\unit_memory/DRAM/n1042 ), 
        .ZN(\unit_memory/DRAM/n1039 ) );
  AOI22_X1 U5441 ( .A1(n154), .A2(\unit_memory/DRAM/n11 ), .B1(n167), .B2(
        \unit_memory/DRAM/n267 ), .ZN(\unit_memory/DRAM/n1042 ) );
  OAI221_X1 U5442 ( .B1(\unit_memory/DRAM/n2409 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2665 ), .C2(n179), .A(\unit_memory/DRAM/n1046 ), 
        .ZN(\unit_memory/DRAM/n1043 ) );
  AOI22_X1 U5443 ( .A1(n153), .A2(\unit_memory/DRAM/n43 ), .B1(n166), .B2(
        \unit_memory/DRAM/n299 ), .ZN(\unit_memory/DRAM/n1046 ) );
  OAI221_X1 U5444 ( .B1(\unit_memory/DRAM/n2378 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2634 ), .C2(n179), .A(\unit_memory/DRAM/n1063 ), 
        .ZN(\unit_memory/DRAM/n1060 ) );
  AOI22_X1 U5445 ( .A1(n153), .A2(\unit_memory/DRAM/n12 ), .B1(n166), .B2(
        \unit_memory/DRAM/n268 ), .ZN(\unit_memory/DRAM/n1063 ) );
  OAI221_X1 U5446 ( .B1(\unit_memory/DRAM/n2410 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2666 ), .C2(n180), .A(\unit_memory/DRAM/n1067 ), 
        .ZN(\unit_memory/DRAM/n1064 ) );
  AOI22_X1 U5447 ( .A1(n154), .A2(\unit_memory/DRAM/n44 ), .B1(n167), .B2(
        \unit_memory/DRAM/n300 ), .ZN(\unit_memory/DRAM/n1067 ) );
  OAI221_X1 U5448 ( .B1(\unit_memory/DRAM/n2379 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2635 ), .C2(n180), .A(\unit_memory/DRAM/n1084 ), 
        .ZN(\unit_memory/DRAM/n1081 ) );
  AOI22_X1 U5449 ( .A1(n154), .A2(\unit_memory/DRAM/n13 ), .B1(n167), .B2(
        \unit_memory/DRAM/n269 ), .ZN(\unit_memory/DRAM/n1084 ) );
  OAI221_X1 U5450 ( .B1(\unit_memory/DRAM/n2411 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2667 ), .C2(n179), .A(\unit_memory/DRAM/n1088 ), 
        .ZN(\unit_memory/DRAM/n1085 ) );
  AOI22_X1 U5451 ( .A1(n153), .A2(\unit_memory/DRAM/n45 ), .B1(n166), .B2(
        \unit_memory/DRAM/n301 ), .ZN(\unit_memory/DRAM/n1088 ) );
  OAI221_X1 U5452 ( .B1(\unit_memory/DRAM/n2380 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2636 ), .C2(n179), .A(\unit_memory/DRAM/n1105 ), 
        .ZN(\unit_memory/DRAM/n1102 ) );
  AOI22_X1 U5453 ( .A1(n153), .A2(\unit_memory/DRAM/n14 ), .B1(n166), .B2(
        \unit_memory/DRAM/n270 ), .ZN(\unit_memory/DRAM/n1105 ) );
  OAI221_X1 U5454 ( .B1(\unit_memory/DRAM/n2412 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2668 ), .C2(n179), .A(\unit_memory/DRAM/n1109 ), 
        .ZN(\unit_memory/DRAM/n1106 ) );
  AOI22_X1 U5455 ( .A1(n153), .A2(\unit_memory/DRAM/n46 ), .B1(n166), .B2(
        \unit_memory/DRAM/n302 ), .ZN(\unit_memory/DRAM/n1109 ) );
  OAI221_X1 U5456 ( .B1(\unit_memory/DRAM/n2381 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2637 ), .C2(n181), .A(\unit_memory/DRAM/n1126 ), 
        .ZN(\unit_memory/DRAM/n1123 ) );
  AOI22_X1 U5457 ( .A1(n155), .A2(\unit_memory/DRAM/n15 ), .B1(n168), .B2(
        \unit_memory/DRAM/n271 ), .ZN(\unit_memory/DRAM/n1126 ) );
  OAI221_X1 U5458 ( .B1(\unit_memory/DRAM/n2413 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2669 ), .C2(n180), .A(\unit_memory/DRAM/n1130 ), 
        .ZN(\unit_memory/DRAM/n1127 ) );
  AOI22_X1 U5459 ( .A1(n154), .A2(\unit_memory/DRAM/n47 ), .B1(n167), .B2(
        \unit_memory/DRAM/n303 ), .ZN(\unit_memory/DRAM/n1130 ) );
  OAI221_X1 U5460 ( .B1(\unit_memory/DRAM/n2382 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2638 ), .C2(n181), .A(\unit_memory/DRAM/n2194 ), 
        .ZN(\unit_memory/DRAM/n2191 ) );
  AOI22_X1 U5461 ( .A1(n155), .A2(\unit_memory/DRAM/n16 ), .B1(n168), .B2(
        \unit_memory/DRAM/n272 ), .ZN(\unit_memory/DRAM/n2194 ) );
  OAI221_X1 U5462 ( .B1(\unit_memory/DRAM/n2414 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2670 ), .C2(n181), .A(\unit_memory/DRAM/n2198 ), 
        .ZN(\unit_memory/DRAM/n2195 ) );
  AOI22_X1 U5463 ( .A1(n155), .A2(\unit_memory/DRAM/n48 ), .B1(n168), .B2(
        \unit_memory/DRAM/n304 ), .ZN(\unit_memory/DRAM/n2198 ) );
  OAI22_X1 U5464 ( .A1(\unit_memory/DRAM/n2719 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2463 ), .B2(n188), .ZN(\unit_memory/DRAM/n820 ) );
  OAI22_X1 U5465 ( .A1(\unit_memory/DRAM/n2847 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2591 ), .B2(n240), .ZN(\unit_memory/DRAM/n821 ) );
  OAI22_X1 U5466 ( .A1(\unit_memory/DRAM/n2720 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2464 ), .B2(n188), .ZN(\unit_memory/DRAM/n844 ) );
  OAI22_X1 U5467 ( .A1(\unit_memory/DRAM/n2848 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2592 ), .B2(n240), .ZN(\unit_memory/DRAM/n845 ) );
  OAI22_X1 U5468 ( .A1(\unit_memory/DRAM/n2721 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2465 ), .B2(n188), .ZN(\unit_memory/DRAM/n865 ) );
  OAI22_X1 U5469 ( .A1(\unit_memory/DRAM/n2849 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2593 ), .B2(n240), .ZN(\unit_memory/DRAM/n866 ) );
  OAI22_X1 U5470 ( .A1(\unit_memory/DRAM/n2722 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2466 ), .B2(n188), .ZN(\unit_memory/DRAM/n886 ) );
  OAI22_X1 U5471 ( .A1(\unit_memory/DRAM/n2850 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2594 ), .B2(n240), .ZN(\unit_memory/DRAM/n887 ) );
  OAI22_X1 U5472 ( .A1(\unit_memory/DRAM/n2723 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2467 ), .B2(n188), .ZN(\unit_memory/DRAM/n907 ) );
  OAI22_X1 U5473 ( .A1(\unit_memory/DRAM/n2851 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2595 ), .B2(n240), .ZN(\unit_memory/DRAM/n908 ) );
  OAI22_X1 U5474 ( .A1(\unit_memory/DRAM/n2724 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2468 ), .B2(n188), .ZN(\unit_memory/DRAM/n928 ) );
  OAI22_X1 U5475 ( .A1(\unit_memory/DRAM/n2852 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2596 ), .B2(n240), .ZN(\unit_memory/DRAM/n929 ) );
  OAI22_X1 U5476 ( .A1(\unit_memory/DRAM/n2725 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2469 ), .B2(n188), .ZN(\unit_memory/DRAM/n949 ) );
  OAI22_X1 U5477 ( .A1(\unit_memory/DRAM/n2853 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2597 ), .B2(n240), .ZN(\unit_memory/DRAM/n950 ) );
  OAI22_X1 U5478 ( .A1(\unit_memory/DRAM/n2726 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2470 ), .B2(n188), .ZN(\unit_memory/DRAM/n970 ) );
  OAI22_X1 U5479 ( .A1(\unit_memory/DRAM/n2854 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2598 ), .B2(n240), .ZN(\unit_memory/DRAM/n971 ) );
  OAI22_X1 U5480 ( .A1(\unit_memory/DRAM/n2727 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2471 ), .B2(n189), .ZN(\unit_memory/DRAM/n991 ) );
  OAI22_X1 U5481 ( .A1(\unit_memory/DRAM/n2855 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2599 ), .B2(n241), .ZN(\unit_memory/DRAM/n992 ) );
  OAI22_X1 U5482 ( .A1(\unit_memory/DRAM/n2728 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2472 ), .B2(n189), .ZN(\unit_memory/DRAM/n1012 ) );
  OAI22_X1 U5483 ( .A1(\unit_memory/DRAM/n2856 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2600 ), .B2(n241), .ZN(\unit_memory/DRAM/n1013 ) );
  OAI22_X1 U5484 ( .A1(\unit_memory/DRAM/n2729 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2473 ), .B2(n189), .ZN(\unit_memory/DRAM/n1033 ) );
  OAI22_X1 U5485 ( .A1(\unit_memory/DRAM/n2857 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2601 ), .B2(n241), .ZN(\unit_memory/DRAM/n1034 ) );
  OAI22_X1 U5486 ( .A1(\unit_memory/DRAM/n2730 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2474 ), .B2(n189), .ZN(\unit_memory/DRAM/n1054 ) );
  OAI22_X1 U5487 ( .A1(\unit_memory/DRAM/n2858 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2602 ), .B2(n241), .ZN(\unit_memory/DRAM/n1055 ) );
  OAI22_X1 U5488 ( .A1(\unit_memory/DRAM/n2731 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2475 ), .B2(n189), .ZN(\unit_memory/DRAM/n1075 ) );
  OAI22_X1 U5489 ( .A1(\unit_memory/DRAM/n2859 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2603 ), .B2(n241), .ZN(\unit_memory/DRAM/n1076 ) );
  OAI22_X1 U5490 ( .A1(\unit_memory/DRAM/n2732 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2476 ), .B2(n189), .ZN(\unit_memory/DRAM/n1096 ) );
  OAI22_X1 U5491 ( .A1(\unit_memory/DRAM/n2860 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2604 ), .B2(n241), .ZN(\unit_memory/DRAM/n1097 ) );
  OAI22_X1 U5492 ( .A1(\unit_memory/DRAM/n2733 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2477 ), .B2(n189), .ZN(\unit_memory/DRAM/n1117 ) );
  OAI22_X1 U5493 ( .A1(\unit_memory/DRAM/n2861 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2605 ), .B2(n241), .ZN(\unit_memory/DRAM/n1118 ) );
  OAI22_X1 U5494 ( .A1(\unit_memory/DRAM/n2734 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2478 ), .B2(n190), .ZN(\unit_memory/DRAM/n2185 ) );
  OAI22_X1 U5495 ( .A1(\unit_memory/DRAM/n2862 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2606 ), .B2(n242), .ZN(\unit_memory/DRAM/n2186 ) );
  OAI22_X1 U5496 ( .A1(\unit_memory/DRAM/n2736 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2480 ), .B2(n189), .ZN(\unit_memory/DRAM/n573 ) );
  OAI22_X1 U5497 ( .A1(\unit_memory/DRAM/n2864 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2608 ), .B2(n241), .ZN(\unit_memory/DRAM/n578 ) );
  OAI22_X1 U5498 ( .A1(\unit_memory/DRAM/n2704 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2448 ), .B2(n186), .ZN(\unit_memory/DRAM/n584 ) );
  OAI22_X1 U5499 ( .A1(\unit_memory/DRAM/n2832 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2576 ), .B2(n238), .ZN(\unit_memory/DRAM/n585 ) );
  OAI22_X1 U5500 ( .A1(\unit_memory/DRAM/n2737 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2481 ), .B2(n186), .ZN(\unit_memory/DRAM/n601 ) );
  OAI22_X1 U5501 ( .A1(\unit_memory/DRAM/n2865 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2609 ), .B2(n238), .ZN(\unit_memory/DRAM/n602 ) );
  OAI22_X1 U5502 ( .A1(\unit_memory/DRAM/n2705 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2449 ), .B2(n186), .ZN(\unit_memory/DRAM/n605 ) );
  OAI22_X1 U5503 ( .A1(\unit_memory/DRAM/n2833 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2577 ), .B2(n238), .ZN(\unit_memory/DRAM/n606 ) );
  OAI22_X1 U5504 ( .A1(\unit_memory/DRAM/n2738 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2482 ), .B2(n186), .ZN(\unit_memory/DRAM/n622 ) );
  OAI22_X1 U5505 ( .A1(\unit_memory/DRAM/n2866 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2610 ), .B2(n238), .ZN(\unit_memory/DRAM/n623 ) );
  OAI22_X1 U5506 ( .A1(\unit_memory/DRAM/n2706 ), .A2(n173), .B1(
        \unit_memory/DRAM/n2450 ), .B2(n186), .ZN(\unit_memory/DRAM/n626 ) );
  OAI22_X1 U5507 ( .A1(\unit_memory/DRAM/n2834 ), .A2(n225), .B1(
        \unit_memory/DRAM/n2578 ), .B2(n238), .ZN(\unit_memory/DRAM/n627 ) );
  OAI22_X1 U5508 ( .A1(\unit_memory/DRAM/n2739 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2483 ), .B2(n187), .ZN(\unit_memory/DRAM/n643 ) );
  OAI22_X1 U5509 ( .A1(\unit_memory/DRAM/n2867 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2611 ), .B2(n239), .ZN(\unit_memory/DRAM/n644 ) );
  OAI22_X1 U5510 ( .A1(\unit_memory/DRAM/n2707 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2451 ), .B2(n187), .ZN(\unit_memory/DRAM/n647 ) );
  OAI22_X1 U5511 ( .A1(\unit_memory/DRAM/n2835 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2579 ), .B2(n239), .ZN(\unit_memory/DRAM/n648 ) );
  OAI22_X1 U5512 ( .A1(\unit_memory/DRAM/n2740 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2484 ), .B2(n187), .ZN(\unit_memory/DRAM/n664 ) );
  OAI22_X1 U5513 ( .A1(\unit_memory/DRAM/n2868 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2612 ), .B2(n239), .ZN(\unit_memory/DRAM/n665 ) );
  OAI22_X1 U5514 ( .A1(\unit_memory/DRAM/n2708 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2452 ), .B2(n187), .ZN(\unit_memory/DRAM/n668 ) );
  OAI22_X1 U5515 ( .A1(\unit_memory/DRAM/n2836 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2580 ), .B2(n239), .ZN(\unit_memory/DRAM/n669 ) );
  OAI22_X1 U5516 ( .A1(\unit_memory/DRAM/n2741 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2485 ), .B2(n187), .ZN(\unit_memory/DRAM/n685 ) );
  OAI22_X1 U5517 ( .A1(\unit_memory/DRAM/n2869 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2613 ), .B2(n239), .ZN(\unit_memory/DRAM/n686 ) );
  OAI22_X1 U5518 ( .A1(\unit_memory/DRAM/n2709 ), .A2(n174), .B1(
        \unit_memory/DRAM/n2453 ), .B2(n187), .ZN(\unit_memory/DRAM/n689 ) );
  OAI22_X1 U5519 ( .A1(\unit_memory/DRAM/n2837 ), .A2(n226), .B1(
        \unit_memory/DRAM/n2581 ), .B2(n239), .ZN(\unit_memory/DRAM/n690 ) );
  OAI22_X1 U5520 ( .A1(\unit_memory/DRAM/n2742 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2486 ), .B2(n188), .ZN(\unit_memory/DRAM/n706 ) );
  OAI22_X1 U5521 ( .A1(\unit_memory/DRAM/n2870 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2614 ), .B2(n240), .ZN(\unit_memory/DRAM/n707 ) );
  OAI22_X1 U5522 ( .A1(\unit_memory/DRAM/n2710 ), .A2(n175), .B1(
        \unit_memory/DRAM/n2454 ), .B2(n188), .ZN(\unit_memory/DRAM/n710 ) );
  OAI22_X1 U5523 ( .A1(\unit_memory/DRAM/n2838 ), .A2(n227), .B1(
        \unit_memory/DRAM/n2582 ), .B2(n240), .ZN(\unit_memory/DRAM/n711 ) );
  OAI22_X1 U5524 ( .A1(\unit_memory/DRAM/n2744 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2488 ), .B2(n190), .ZN(\unit_memory/DRAM/n2227 ) );
  OAI22_X1 U5525 ( .A1(\unit_memory/DRAM/n2872 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2616 ), .B2(n242), .ZN(\unit_memory/DRAM/n2228 ) );
  OAI22_X1 U5526 ( .A1(\unit_memory/DRAM/n2712 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2456 ), .B2(n190), .ZN(\unit_memory/DRAM/n2231 ) );
  OAI22_X1 U5527 ( .A1(\unit_memory/DRAM/n2840 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2584 ), .B2(n242), .ZN(\unit_memory/DRAM/n2232 ) );
  OAI22_X1 U5528 ( .A1(\unit_memory/DRAM/n2745 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2489 ), .B2(n191), .ZN(\unit_memory/DRAM/n2248 ) );
  OAI22_X1 U5529 ( .A1(\unit_memory/DRAM/n2873 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2617 ), .B2(n243), .ZN(\unit_memory/DRAM/n2249 ) );
  OAI22_X1 U5530 ( .A1(\unit_memory/DRAM/n2713 ), .A2(n176), .B1(
        \unit_memory/DRAM/n2457 ), .B2(n189), .ZN(\unit_memory/DRAM/n2252 ) );
  OAI22_X1 U5531 ( .A1(\unit_memory/DRAM/n2841 ), .A2(n228), .B1(
        \unit_memory/DRAM/n2585 ), .B2(n241), .ZN(\unit_memory/DRAM/n2253 ) );
  OAI22_X1 U5532 ( .A1(\unit_memory/DRAM/n2746 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2490 ), .B2(n190), .ZN(\unit_memory/DRAM/n2269 ) );
  OAI22_X1 U5533 ( .A1(\unit_memory/DRAM/n2874 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2618 ), .B2(n242), .ZN(\unit_memory/DRAM/n2270 ) );
  OAI22_X1 U5534 ( .A1(\unit_memory/DRAM/n2714 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2458 ), .B2(n190), .ZN(\unit_memory/DRAM/n2273 ) );
  OAI22_X1 U5535 ( .A1(\unit_memory/DRAM/n2842 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2586 ), .B2(n242), .ZN(\unit_memory/DRAM/n2274 ) );
  OAI22_X1 U5536 ( .A1(\unit_memory/DRAM/n2747 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2491 ), .B2(n190), .ZN(\unit_memory/DRAM/n2290 ) );
  OAI22_X1 U5537 ( .A1(\unit_memory/DRAM/n2875 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2619 ), .B2(n242), .ZN(\unit_memory/DRAM/n2291 ) );
  OAI22_X1 U5538 ( .A1(\unit_memory/DRAM/n2715 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2459 ), .B2(n191), .ZN(\unit_memory/DRAM/n2294 ) );
  OAI22_X1 U5539 ( .A1(\unit_memory/DRAM/n2843 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2587 ), .B2(n243), .ZN(\unit_memory/DRAM/n2295 ) );
  OAI22_X1 U5540 ( .A1(\unit_memory/DRAM/n2748 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2492 ), .B2(n191), .ZN(\unit_memory/DRAM/n2311 ) );
  OAI22_X1 U5541 ( .A1(\unit_memory/DRAM/n2876 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2620 ), .B2(n243), .ZN(\unit_memory/DRAM/n2312 ) );
  OAI22_X1 U5542 ( .A1(\unit_memory/DRAM/n2716 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2460 ), .B2(n190), .ZN(\unit_memory/DRAM/n2315 ) );
  OAI22_X1 U5543 ( .A1(\unit_memory/DRAM/n2844 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2588 ), .B2(n242), .ZN(\unit_memory/DRAM/n2316 ) );
  OAI22_X1 U5544 ( .A1(\unit_memory/DRAM/n2749 ), .A2(n177), .B1(
        \unit_memory/DRAM/n2493 ), .B2(n190), .ZN(\unit_memory/DRAM/n2332 ) );
  OAI22_X1 U5545 ( .A1(\unit_memory/DRAM/n2877 ), .A2(n229), .B1(
        \unit_memory/DRAM/n2621 ), .B2(n242), .ZN(\unit_memory/DRAM/n2333 ) );
  OAI22_X1 U5546 ( .A1(\unit_memory/DRAM/n2717 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2461 ), .B2(n191), .ZN(\unit_memory/DRAM/n2336 ) );
  OAI22_X1 U5547 ( .A1(\unit_memory/DRAM/n2845 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2589 ), .B2(n243), .ZN(\unit_memory/DRAM/n2337 ) );
  OAI22_X1 U5548 ( .A1(\unit_memory/DRAM/n2750 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2494 ), .B2(n191), .ZN(\unit_memory/DRAM/n2353 ) );
  OAI22_X1 U5549 ( .A1(\unit_memory/DRAM/n2878 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2622 ), .B2(n243), .ZN(\unit_memory/DRAM/n2354 ) );
  OAI22_X1 U5550 ( .A1(\unit_memory/DRAM/n2718 ), .A2(n178), .B1(
        \unit_memory/DRAM/n2462 ), .B2(n191), .ZN(\unit_memory/DRAM/n2357 ) );
  OAI22_X1 U5551 ( .A1(\unit_memory/DRAM/n2846 ), .A2(n230), .B1(
        \unit_memory/DRAM/n2590 ), .B2(n243), .ZN(\unit_memory/DRAM/n2358 ) );
  AOI22_X1 U5552 ( .A1(n209), .A2(\unit_memory/DRAM/n153 ), .B1(n222), .B2(
        \unit_memory/DRAM/n409 ), .ZN(\unit_memory/DRAM/n2206 ) );
  AOI22_X1 U5553 ( .A1(n209), .A2(\unit_memory/DRAM/n217 ), .B1(n222), .B2(
        \unit_memory/DRAM/n473 ), .ZN(\unit_memory/DRAM/n2214 ) );
  AOI22_X1 U5554 ( .A1(n209), .A2(\unit_memory/DRAM/n194 ), .B1(n222), .B2(
        \unit_memory/DRAM/n450 ), .ZN(\unit_memory/DRAM/n848 ) );
  AOI22_X1 U5555 ( .A1(n208), .A2(\unit_memory/DRAM/n145 ), .B1(n221), .B2(
        \unit_memory/DRAM/n401 ), .ZN(\unit_memory/DRAM/n1144 ) );
  AOI22_X1 U5556 ( .A1(n208), .A2(\unit_memory/DRAM/n193 ), .B1(n221), .B2(
        \unit_memory/DRAM/n449 ), .ZN(\unit_memory/DRAM/n825 ) );
  AOI22_X1 U5557 ( .A1(n207), .A2(\unit_memory/DRAM/n195 ), .B1(n220), .B2(
        \unit_memory/DRAM/n451 ), .ZN(\unit_memory/DRAM/n869 ) );
  AOI22_X1 U5558 ( .A1(n207), .A2(\unit_memory/DRAM/n196 ), .B1(n220), .B2(
        \unit_memory/DRAM/n452 ), .ZN(\unit_memory/DRAM/n890 ) );
  AOI22_X1 U5559 ( .A1(n208), .A2(\unit_memory/DRAM/n197 ), .B1(n221), .B2(
        \unit_memory/DRAM/n453 ), .ZN(\unit_memory/DRAM/n911 ) );
  AOI22_X1 U5560 ( .A1(n208), .A2(\unit_memory/DRAM/n198 ), .B1(n221), .B2(
        \unit_memory/DRAM/n454 ), .ZN(\unit_memory/DRAM/n932 ) );
  AOI22_X1 U5561 ( .A1(n206), .A2(\unit_memory/DRAM/n199 ), .B1(n219), .B2(
        \unit_memory/DRAM/n455 ), .ZN(\unit_memory/DRAM/n953 ) );
  AOI22_X1 U5562 ( .A1(n207), .A2(\unit_memory/DRAM/n200 ), .B1(n220), .B2(
        \unit_memory/DRAM/n456 ), .ZN(\unit_memory/DRAM/n974 ) );
  AOI22_X1 U5563 ( .A1(n205), .A2(\unit_memory/DRAM/n201 ), .B1(n218), .B2(
        \unit_memory/DRAM/n457 ), .ZN(\unit_memory/DRAM/n995 ) );
  AOI22_X1 U5564 ( .A1(n205), .A2(\unit_memory/DRAM/n202 ), .B1(n218), .B2(
        \unit_memory/DRAM/n458 ), .ZN(\unit_memory/DRAM/n1016 ) );
  AOI22_X1 U5565 ( .A1(n207), .A2(\unit_memory/DRAM/n203 ), .B1(n220), .B2(
        \unit_memory/DRAM/n459 ), .ZN(\unit_memory/DRAM/n1037 ) );
  AOI22_X1 U5566 ( .A1(n205), .A2(\unit_memory/DRAM/n204 ), .B1(n218), .B2(
        \unit_memory/DRAM/n460 ), .ZN(\unit_memory/DRAM/n1058 ) );
  AOI22_X1 U5567 ( .A1(n206), .A2(\unit_memory/DRAM/n205 ), .B1(n219), .B2(
        \unit_memory/DRAM/n461 ), .ZN(\unit_memory/DRAM/n1079 ) );
  AOI22_X1 U5568 ( .A1(n206), .A2(\unit_memory/DRAM/n206 ), .B1(n219), .B2(
        \unit_memory/DRAM/n462 ), .ZN(\unit_memory/DRAM/n1100 ) );
  AOI22_X1 U5569 ( .A1(n205), .A2(\unit_memory/DRAM/n207 ), .B1(n218), .B2(
        \unit_memory/DRAM/n463 ), .ZN(\unit_memory/DRAM/n1121 ) );
  AOI22_X1 U5570 ( .A1(n208), .A2(\unit_memory/DRAM/n208 ), .B1(n221), .B2(
        \unit_memory/DRAM/n464 ), .ZN(\unit_memory/DRAM/n2189 ) );
  AOI22_X1 U5571 ( .A1(n1183), .A2(\unit_decode/n186 ), .B1(n1188), .B2(
        \unit_decode/n166 ), .ZN(\unit_decode/n2890 ) );
  AOI22_X1 U5572 ( .A1(n1183), .A2(\unit_decode/n185 ), .B1(n1188), .B2(
        \unit_decode/n163 ), .ZN(\unit_decode/n2861 ) );
  AOI22_X1 U5573 ( .A1(n1183), .A2(\unit_decode/n184 ), .B1(n1188), .B2(
        \unit_decode/n160 ), .ZN(\unit_decode/n2843 ) );
  AOI22_X1 U5574 ( .A1(n1183), .A2(\unit_decode/n183 ), .B1(n1188), .B2(
        \unit_decode/n157 ), .ZN(\unit_decode/n2825 ) );
  AOI22_X1 U5575 ( .A1(n1183), .A2(\unit_decode/n182 ), .B1(n1188), .B2(
        \unit_decode/n154 ), .ZN(\unit_decode/n2807 ) );
  AOI22_X1 U5576 ( .A1(n1183), .A2(\unit_decode/n181 ), .B1(n1188), .B2(
        \unit_decode/n151 ), .ZN(\unit_decode/n2789 ) );
  AOI22_X1 U5577 ( .A1(n1183), .A2(\unit_decode/n180 ), .B1(n1188), .B2(
        \unit_decode/n148 ), .ZN(\unit_decode/n2771 ) );
  AOI22_X1 U5578 ( .A1(n1183), .A2(\unit_decode/n179 ), .B1(n1188), .B2(
        \unit_decode/n145 ), .ZN(\unit_decode/n2753 ) );
  AOI22_X1 U5579 ( .A1(n1183), .A2(\unit_decode/n178 ), .B1(n1187), .B2(
        \unit_decode/n142 ), .ZN(\unit_decode/n2735 ) );
  AOI22_X1 U5580 ( .A1(n1183), .A2(\unit_decode/n177 ), .B1(n1187), .B2(
        \unit_decode/n139 ), .ZN(\unit_decode/n2717 ) );
  AOI22_X1 U5581 ( .A1(n1183), .A2(\unit_decode/n176 ), .B1(n1187), .B2(
        \unit_decode/n136 ), .ZN(\unit_decode/n2699 ) );
  AOI22_X1 U5582 ( .A1(n1183), .A2(\unit_decode/n175 ), .B1(n1187), .B2(
        \unit_decode/n133 ), .ZN(\unit_decode/n2681 ) );
  AOI22_X1 U5583 ( .A1(n1184), .A2(\unit_decode/n174 ), .B1(n1187), .B2(
        \unit_decode/n130 ), .ZN(\unit_decode/n2663 ) );
  AOI22_X1 U5584 ( .A1(n1184), .A2(\unit_decode/n173 ), .B1(n1187), .B2(
        \unit_decode/n127 ), .ZN(\unit_decode/n2645 ) );
  AOI22_X1 U5585 ( .A1(n1184), .A2(\unit_decode/n172 ), .B1(n1187), .B2(
        \unit_decode/n124 ), .ZN(\unit_decode/n2627 ) );
  AOI22_X1 U5586 ( .A1(n1184), .A2(\unit_decode/n171 ), .B1(n1187), .B2(
        \unit_decode/n121 ), .ZN(\unit_decode/n2609 ) );
  AOI22_X1 U5587 ( .A1(n1184), .A2(\unit_decode/n170 ), .B1(n1187), .B2(
        \unit_decode/n118 ), .ZN(\unit_decode/n2591 ) );
  AOI22_X1 U5588 ( .A1(n1184), .A2(\unit_decode/n169 ), .B1(n1187), .B2(
        \unit_decode/n115 ), .ZN(\unit_decode/n2573 ) );
  AOI22_X1 U5589 ( .A1(n1184), .A2(\unit_decode/n192 ), .B1(n1187), .B2(
        \unit_decode/n112 ), .ZN(\unit_decode/n2555 ) );
  AOI22_X1 U5590 ( .A1(n1184), .A2(\unit_decode/n191 ), .B1(n1187), .B2(
        \unit_decode/n109 ), .ZN(\unit_decode/n2537 ) );
  AOI22_X1 U5591 ( .A1(n1184), .A2(\unit_decode/n190 ), .B1(n1186), .B2(
        \unit_decode/n106 ), .ZN(\unit_decode/n2519 ) );
  AOI22_X1 U5592 ( .A1(n1184), .A2(\unit_decode/n189 ), .B1(n1186), .B2(
        \unit_decode/n103 ), .ZN(\unit_decode/n2501 ) );
  AOI22_X1 U5593 ( .A1(n1184), .A2(\unit_decode/n188 ), .B1(n1186), .B2(
        \unit_decode/n100 ), .ZN(\unit_decode/n2483 ) );
  AOI22_X1 U5594 ( .A1(n1184), .A2(\unit_decode/n187 ), .B1(n1186), .B2(
        \unit_decode/n97 ), .ZN(\unit_decode/n2465 ) );
  AOI22_X1 U5595 ( .A1(n1279), .A2(\unit_decode/n186 ), .B1(n1284), .B2(
        \unit_decode/n166 ), .ZN(\unit_decode/n3510 ) );
  AOI22_X1 U5596 ( .A1(n1279), .A2(\unit_decode/n185 ), .B1(n1284), .B2(
        \unit_decode/n163 ), .ZN(\unit_decode/n3481 ) );
  AOI22_X1 U5597 ( .A1(n1279), .A2(\unit_decode/n184 ), .B1(n1284), .B2(
        \unit_decode/n160 ), .ZN(\unit_decode/n3463 ) );
  AOI22_X1 U5598 ( .A1(n1279), .A2(\unit_decode/n183 ), .B1(n1284), .B2(
        \unit_decode/n157 ), .ZN(\unit_decode/n3445 ) );
  AOI22_X1 U5599 ( .A1(n1279), .A2(\unit_decode/n182 ), .B1(n1284), .B2(
        \unit_decode/n154 ), .ZN(\unit_decode/n3427 ) );
  AOI22_X1 U5600 ( .A1(n1279), .A2(\unit_decode/n181 ), .B1(n1284), .B2(
        \unit_decode/n151 ), .ZN(\unit_decode/n3409 ) );
  AOI22_X1 U5601 ( .A1(n1279), .A2(\unit_decode/n180 ), .B1(n1284), .B2(
        \unit_decode/n148 ), .ZN(\unit_decode/n3391 ) );
  AOI22_X1 U5602 ( .A1(n1279), .A2(\unit_decode/n179 ), .B1(n1284), .B2(
        \unit_decode/n145 ), .ZN(\unit_decode/n3373 ) );
  AOI22_X1 U5603 ( .A1(n1279), .A2(\unit_decode/n178 ), .B1(n1283), .B2(
        \unit_decode/n142 ), .ZN(\unit_decode/n3355 ) );
  AOI22_X1 U5604 ( .A1(n1279), .A2(\unit_decode/n177 ), .B1(n1283), .B2(
        \unit_decode/n139 ), .ZN(\unit_decode/n3337 ) );
  AOI22_X1 U5605 ( .A1(n1279), .A2(\unit_decode/n176 ), .B1(n1283), .B2(
        \unit_decode/n136 ), .ZN(\unit_decode/n3319 ) );
  AOI22_X1 U5606 ( .A1(n1279), .A2(\unit_decode/n175 ), .B1(n1283), .B2(
        \unit_decode/n133 ), .ZN(\unit_decode/n3301 ) );
  AOI22_X1 U5607 ( .A1(n1280), .A2(\unit_decode/n174 ), .B1(n1283), .B2(
        \unit_decode/n130 ), .ZN(\unit_decode/n3283 ) );
  AOI22_X1 U5608 ( .A1(n1280), .A2(\unit_decode/n173 ), .B1(n1283), .B2(
        \unit_decode/n127 ), .ZN(\unit_decode/n3265 ) );
  AOI22_X1 U5609 ( .A1(n1280), .A2(\unit_decode/n172 ), .B1(n1283), .B2(
        \unit_decode/n124 ), .ZN(\unit_decode/n3247 ) );
  AOI22_X1 U5610 ( .A1(n1280), .A2(\unit_decode/n171 ), .B1(n1283), .B2(
        \unit_decode/n121 ), .ZN(\unit_decode/n3229 ) );
  AOI22_X1 U5611 ( .A1(n1280), .A2(\unit_decode/n170 ), .B1(n1283), .B2(
        \unit_decode/n118 ), .ZN(\unit_decode/n3211 ) );
  AOI22_X1 U5612 ( .A1(n1280), .A2(\unit_decode/n169 ), .B1(n1283), .B2(
        \unit_decode/n115 ), .ZN(\unit_decode/n3193 ) );
  AOI22_X1 U5613 ( .A1(n1280), .A2(\unit_decode/n192 ), .B1(n1283), .B2(
        \unit_decode/n112 ), .ZN(\unit_decode/n3175 ) );
  AOI22_X1 U5614 ( .A1(n1280), .A2(\unit_decode/n191 ), .B1(n1283), .B2(
        \unit_decode/n109 ), .ZN(\unit_decode/n3157 ) );
  AOI22_X1 U5615 ( .A1(n1280), .A2(\unit_decode/n190 ), .B1(n1282), .B2(
        \unit_decode/n106 ), .ZN(\unit_decode/n3139 ) );
  AOI22_X1 U5616 ( .A1(n1280), .A2(\unit_decode/n189 ), .B1(n1282), .B2(
        \unit_decode/n103 ), .ZN(\unit_decode/n3121 ) );
  AOI22_X1 U5617 ( .A1(n1280), .A2(\unit_decode/n188 ), .B1(n1282), .B2(
        \unit_decode/n100 ), .ZN(\unit_decode/n3103 ) );
  AOI22_X1 U5618 ( .A1(n1280), .A2(\unit_decode/n187 ), .B1(n1282), .B2(
        \unit_decode/n97 ), .ZN(\unit_decode/n3085 ) );
  AOI21_X1 U5619 ( .B1(\unit_memory/DRAM/n817 ), .B2(\unit_memory/DRAM/n818 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n815 ) );
  AOI221_X1 U5620 ( .B1(n201), .B2(\unit_memory/DRAM/n225 ), .C1(n214), .C2(
        \unit_memory/DRAM/n481 ), .A(\unit_memory/DRAM/n821 ), .ZN(
        \unit_memory/DRAM/n817 ) );
  AOI221_X1 U5621 ( .B1(n149), .B2(\unit_memory/DRAM/n97 ), .C1(n162), .C2(
        \unit_memory/DRAM/n353 ), .A(\unit_memory/DRAM/n820 ), .ZN(
        \unit_memory/DRAM/n818 ) );
  AOI21_X1 U5622 ( .B1(\unit_memory/DRAM/n842 ), .B2(\unit_memory/DRAM/n843 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n841 ) );
  AOI221_X1 U5623 ( .B1(n201), .B2(\unit_memory/DRAM/n226 ), .C1(n214), .C2(
        \unit_memory/DRAM/n482 ), .A(\unit_memory/DRAM/n845 ), .ZN(
        \unit_memory/DRAM/n842 ) );
  AOI221_X1 U5624 ( .B1(n149), .B2(\unit_memory/DRAM/n98 ), .C1(n162), .C2(
        \unit_memory/DRAM/n354 ), .A(\unit_memory/DRAM/n844 ), .ZN(
        \unit_memory/DRAM/n843 ) );
  AOI21_X1 U5625 ( .B1(\unit_memory/DRAM/n863 ), .B2(\unit_memory/DRAM/n864 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n862 ) );
  AOI221_X1 U5626 ( .B1(n201), .B2(\unit_memory/DRAM/n227 ), .C1(n214), .C2(
        \unit_memory/DRAM/n483 ), .A(\unit_memory/DRAM/n866 ), .ZN(
        \unit_memory/DRAM/n863 ) );
  AOI221_X1 U5627 ( .B1(n149), .B2(\unit_memory/DRAM/n99 ), .C1(n162), .C2(
        \unit_memory/DRAM/n355 ), .A(\unit_memory/DRAM/n865 ), .ZN(
        \unit_memory/DRAM/n864 ) );
  AOI21_X1 U5628 ( .B1(\unit_memory/DRAM/n884 ), .B2(\unit_memory/DRAM/n885 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n883 ) );
  AOI221_X1 U5629 ( .B1(n201), .B2(\unit_memory/DRAM/n228 ), .C1(n214), .C2(
        \unit_memory/DRAM/n484 ), .A(\unit_memory/DRAM/n887 ), .ZN(
        \unit_memory/DRAM/n884 ) );
  AOI221_X1 U5630 ( .B1(n149), .B2(\unit_memory/DRAM/n100 ), .C1(n162), .C2(
        \unit_memory/DRAM/n356 ), .A(\unit_memory/DRAM/n886 ), .ZN(
        \unit_memory/DRAM/n885 ) );
  AOI21_X1 U5631 ( .B1(\unit_memory/DRAM/n905 ), .B2(\unit_memory/DRAM/n906 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n904 ) );
  AOI221_X1 U5632 ( .B1(n201), .B2(\unit_memory/DRAM/n229 ), .C1(n214), .C2(
        \unit_memory/DRAM/n485 ), .A(\unit_memory/DRAM/n908 ), .ZN(
        \unit_memory/DRAM/n905 ) );
  AOI221_X1 U5633 ( .B1(n149), .B2(\unit_memory/DRAM/n101 ), .C1(n162), .C2(
        \unit_memory/DRAM/n357 ), .A(\unit_memory/DRAM/n907 ), .ZN(
        \unit_memory/DRAM/n906 ) );
  AOI21_X1 U5634 ( .B1(\unit_memory/DRAM/n926 ), .B2(\unit_memory/DRAM/n927 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n925 ) );
  AOI221_X1 U5635 ( .B1(n201), .B2(\unit_memory/DRAM/n230 ), .C1(n214), .C2(
        \unit_memory/DRAM/n486 ), .A(\unit_memory/DRAM/n929 ), .ZN(
        \unit_memory/DRAM/n926 ) );
  AOI221_X1 U5636 ( .B1(n149), .B2(\unit_memory/DRAM/n102 ), .C1(n162), .C2(
        \unit_memory/DRAM/n358 ), .A(\unit_memory/DRAM/n928 ), .ZN(
        \unit_memory/DRAM/n927 ) );
  AOI21_X1 U5637 ( .B1(\unit_memory/DRAM/n947 ), .B2(\unit_memory/DRAM/n948 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n946 ) );
  AOI221_X1 U5638 ( .B1(n201), .B2(\unit_memory/DRAM/n231 ), .C1(n214), .C2(
        \unit_memory/DRAM/n487 ), .A(\unit_memory/DRAM/n950 ), .ZN(
        \unit_memory/DRAM/n947 ) );
  AOI221_X1 U5639 ( .B1(n149), .B2(\unit_memory/DRAM/n103 ), .C1(n162), .C2(
        \unit_memory/DRAM/n359 ), .A(\unit_memory/DRAM/n949 ), .ZN(
        \unit_memory/DRAM/n948 ) );
  AOI21_X1 U5640 ( .B1(\unit_memory/DRAM/n968 ), .B2(\unit_memory/DRAM/n969 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n967 ) );
  AOI221_X1 U5641 ( .B1(n201), .B2(\unit_memory/DRAM/n232 ), .C1(n214), .C2(
        \unit_memory/DRAM/n488 ), .A(\unit_memory/DRAM/n971 ), .ZN(
        \unit_memory/DRAM/n968 ) );
  AOI221_X1 U5642 ( .B1(n149), .B2(\unit_memory/DRAM/n104 ), .C1(n162), .C2(
        \unit_memory/DRAM/n360 ), .A(\unit_memory/DRAM/n970 ), .ZN(
        \unit_memory/DRAM/n969 ) );
  AOI21_X1 U5643 ( .B1(\unit_memory/DRAM/n989 ), .B2(\unit_memory/DRAM/n990 ), 
        .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n988 ) );
  AOI221_X1 U5644 ( .B1(n202), .B2(\unit_memory/DRAM/n233 ), .C1(n215), .C2(
        \unit_memory/DRAM/n489 ), .A(\unit_memory/DRAM/n992 ), .ZN(
        \unit_memory/DRAM/n989 ) );
  AOI221_X1 U5645 ( .B1(n150), .B2(\unit_memory/DRAM/n105 ), .C1(n163), .C2(
        \unit_memory/DRAM/n361 ), .A(\unit_memory/DRAM/n991 ), .ZN(
        \unit_memory/DRAM/n990 ) );
  AOI21_X1 U5646 ( .B1(\unit_memory/DRAM/n1010 ), .B2(\unit_memory/DRAM/n1011 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1009 ) );
  AOI221_X1 U5647 ( .B1(n202), .B2(\unit_memory/DRAM/n234 ), .C1(n215), .C2(
        \unit_memory/DRAM/n490 ), .A(\unit_memory/DRAM/n1013 ), .ZN(
        \unit_memory/DRAM/n1010 ) );
  AOI221_X1 U5648 ( .B1(n150), .B2(\unit_memory/DRAM/n106 ), .C1(n163), .C2(
        \unit_memory/DRAM/n362 ), .A(\unit_memory/DRAM/n1012 ), .ZN(
        \unit_memory/DRAM/n1011 ) );
  AOI21_X1 U5649 ( .B1(\unit_memory/DRAM/n1031 ), .B2(\unit_memory/DRAM/n1032 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1030 ) );
  AOI221_X1 U5650 ( .B1(n202), .B2(\unit_memory/DRAM/n235 ), .C1(n215), .C2(
        \unit_memory/DRAM/n491 ), .A(\unit_memory/DRAM/n1034 ), .ZN(
        \unit_memory/DRAM/n1031 ) );
  AOI221_X1 U5651 ( .B1(n150), .B2(\unit_memory/DRAM/n107 ), .C1(n163), .C2(
        \unit_memory/DRAM/n363 ), .A(\unit_memory/DRAM/n1033 ), .ZN(
        \unit_memory/DRAM/n1032 ) );
  AOI21_X1 U5652 ( .B1(\unit_memory/DRAM/n1052 ), .B2(\unit_memory/DRAM/n1053 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1051 ) );
  AOI221_X1 U5653 ( .B1(n202), .B2(\unit_memory/DRAM/n236 ), .C1(n215), .C2(
        \unit_memory/DRAM/n492 ), .A(\unit_memory/DRAM/n1055 ), .ZN(
        \unit_memory/DRAM/n1052 ) );
  AOI221_X1 U5654 ( .B1(n150), .B2(\unit_memory/DRAM/n108 ), .C1(n163), .C2(
        \unit_memory/DRAM/n364 ), .A(\unit_memory/DRAM/n1054 ), .ZN(
        \unit_memory/DRAM/n1053 ) );
  AOI21_X1 U5655 ( .B1(\unit_memory/DRAM/n1073 ), .B2(\unit_memory/DRAM/n1074 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1072 ) );
  AOI221_X1 U5656 ( .B1(n202), .B2(\unit_memory/DRAM/n237 ), .C1(n215), .C2(
        \unit_memory/DRAM/n493 ), .A(\unit_memory/DRAM/n1076 ), .ZN(
        \unit_memory/DRAM/n1073 ) );
  AOI221_X1 U5657 ( .B1(n150), .B2(\unit_memory/DRAM/n109 ), .C1(n163), .C2(
        \unit_memory/DRAM/n365 ), .A(\unit_memory/DRAM/n1075 ), .ZN(
        \unit_memory/DRAM/n1074 ) );
  AOI21_X1 U5658 ( .B1(\unit_memory/DRAM/n1094 ), .B2(\unit_memory/DRAM/n1095 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1093 ) );
  AOI221_X1 U5659 ( .B1(n202), .B2(\unit_memory/DRAM/n238 ), .C1(n215), .C2(
        \unit_memory/DRAM/n494 ), .A(\unit_memory/DRAM/n1097 ), .ZN(
        \unit_memory/DRAM/n1094 ) );
  AOI221_X1 U5660 ( .B1(n150), .B2(\unit_memory/DRAM/n110 ), .C1(n163), .C2(
        \unit_memory/DRAM/n366 ), .A(\unit_memory/DRAM/n1096 ), .ZN(
        \unit_memory/DRAM/n1095 ) );
  AOI21_X1 U5661 ( .B1(\unit_memory/DRAM/n1115 ), .B2(\unit_memory/DRAM/n1116 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1114 ) );
  AOI221_X1 U5662 ( .B1(n202), .B2(\unit_memory/DRAM/n239 ), .C1(n215), .C2(
        \unit_memory/DRAM/n495 ), .A(\unit_memory/DRAM/n1118 ), .ZN(
        \unit_memory/DRAM/n1115 ) );
  AOI221_X1 U5663 ( .B1(n150), .B2(\unit_memory/DRAM/n111 ), .C1(n163), .C2(
        \unit_memory/DRAM/n367 ), .A(\unit_memory/DRAM/n1117 ), .ZN(
        \unit_memory/DRAM/n1116 ) );
  AOI21_X1 U5664 ( .B1(\unit_memory/DRAM/n2183 ), .B2(\unit_memory/DRAM/n2184 ), .A(\unit_memory/DRAM/n819 ), .ZN(\unit_memory/DRAM/n1135 ) );
  AOI221_X1 U5665 ( .B1(n203), .B2(\unit_memory/DRAM/n240 ), .C1(n216), .C2(
        \unit_memory/DRAM/n496 ), .A(\unit_memory/DRAM/n2186 ), .ZN(
        \unit_memory/DRAM/n2183 ) );
  AOI221_X1 U5666 ( .B1(n151), .B2(\unit_memory/DRAM/n112 ), .C1(n164), .C2(
        \unit_memory/DRAM/n368 ), .A(\unit_memory/DRAM/n2185 ), .ZN(
        \unit_memory/DRAM/n2184 ) );
  OAI21_X1 U5667 ( .B1(\unit_memory/DRAM/n822 ), .B2(\unit_memory/DRAM/n823 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n813 ) );
  OAI221_X1 U5668 ( .B1(\unit_memory/DRAM/n2431 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2687 ), .C2(n182), .A(\unit_memory/DRAM/n826 ), 
        .ZN(\unit_memory/DRAM/n822 ) );
  OAI221_X1 U5669 ( .B1(\unit_memory/DRAM/n2559 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2815 ), .C2(n234), .A(\unit_memory/DRAM/n825 ), 
        .ZN(\unit_memory/DRAM/n823 ) );
  AOI22_X1 U5670 ( .A1(n156), .A2(\unit_memory/DRAM/n65 ), .B1(n169), .B2(
        \unit_memory/DRAM/n321 ), .ZN(\unit_memory/DRAM/n826 ) );
  OAI21_X1 U5671 ( .B1(\unit_memory/DRAM/n846 ), .B2(\unit_memory/DRAM/n847 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n839 ) );
  OAI221_X1 U5672 ( .B1(\unit_memory/DRAM/n2432 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2688 ), .C2(n183), .A(\unit_memory/DRAM/n849 ), 
        .ZN(\unit_memory/DRAM/n846 ) );
  OAI221_X1 U5673 ( .B1(\unit_memory/DRAM/n2560 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2816 ), .C2(n235), .A(\unit_memory/DRAM/n848 ), 
        .ZN(\unit_memory/DRAM/n847 ) );
  AOI22_X1 U5674 ( .A1(n157), .A2(\unit_memory/DRAM/n66 ), .B1(n170), .B2(
        \unit_memory/DRAM/n322 ), .ZN(\unit_memory/DRAM/n849 ) );
  OAI21_X1 U5675 ( .B1(\unit_memory/DRAM/n867 ), .B2(\unit_memory/DRAM/n868 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n860 ) );
  OAI221_X1 U5676 ( .B1(\unit_memory/DRAM/n2433 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2689 ), .C2(n181), .A(\unit_memory/DRAM/n870 ), 
        .ZN(\unit_memory/DRAM/n867 ) );
  OAI221_X1 U5677 ( .B1(\unit_memory/DRAM/n2561 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2817 ), .C2(n233), .A(\unit_memory/DRAM/n869 ), 
        .ZN(\unit_memory/DRAM/n868 ) );
  AOI22_X1 U5678 ( .A1(n155), .A2(\unit_memory/DRAM/n67 ), .B1(n168), .B2(
        \unit_memory/DRAM/n323 ), .ZN(\unit_memory/DRAM/n870 ) );
  OAI21_X1 U5679 ( .B1(\unit_memory/DRAM/n888 ), .B2(\unit_memory/DRAM/n889 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n881 ) );
  OAI221_X1 U5680 ( .B1(\unit_memory/DRAM/n2434 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2690 ), .C2(n181), .A(\unit_memory/DRAM/n891 ), 
        .ZN(\unit_memory/DRAM/n888 ) );
  OAI221_X1 U5681 ( .B1(\unit_memory/DRAM/n2562 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2818 ), .C2(n233), .A(\unit_memory/DRAM/n890 ), 
        .ZN(\unit_memory/DRAM/n889 ) );
  AOI22_X1 U5682 ( .A1(n155), .A2(\unit_memory/DRAM/n68 ), .B1(n168), .B2(
        \unit_memory/DRAM/n324 ), .ZN(\unit_memory/DRAM/n891 ) );
  OAI21_X1 U5683 ( .B1(\unit_memory/DRAM/n909 ), .B2(\unit_memory/DRAM/n910 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n902 ) );
  OAI221_X1 U5684 ( .B1(\unit_memory/DRAM/n2435 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2691 ), .C2(n182), .A(\unit_memory/DRAM/n912 ), 
        .ZN(\unit_memory/DRAM/n909 ) );
  OAI221_X1 U5685 ( .B1(\unit_memory/DRAM/n2563 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2819 ), .C2(n234), .A(\unit_memory/DRAM/n911 ), 
        .ZN(\unit_memory/DRAM/n910 ) );
  AOI22_X1 U5686 ( .A1(n156), .A2(\unit_memory/DRAM/n69 ), .B1(n169), .B2(
        \unit_memory/DRAM/n325 ), .ZN(\unit_memory/DRAM/n912 ) );
  OAI21_X1 U5687 ( .B1(\unit_memory/DRAM/n930 ), .B2(\unit_memory/DRAM/n931 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n923 ) );
  OAI221_X1 U5688 ( .B1(\unit_memory/DRAM/n2436 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2692 ), .C2(n182), .A(\unit_memory/DRAM/n933 ), 
        .ZN(\unit_memory/DRAM/n930 ) );
  OAI221_X1 U5689 ( .B1(\unit_memory/DRAM/n2564 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2820 ), .C2(n234), .A(\unit_memory/DRAM/n932 ), 
        .ZN(\unit_memory/DRAM/n931 ) );
  AOI22_X1 U5690 ( .A1(n156), .A2(\unit_memory/DRAM/n70 ), .B1(n169), .B2(
        \unit_memory/DRAM/n326 ), .ZN(\unit_memory/DRAM/n933 ) );
  OAI21_X1 U5691 ( .B1(\unit_memory/DRAM/n951 ), .B2(\unit_memory/DRAM/n952 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n944 ) );
  OAI221_X1 U5692 ( .B1(\unit_memory/DRAM/n2437 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2693 ), .C2(n180), .A(\unit_memory/DRAM/n954 ), 
        .ZN(\unit_memory/DRAM/n951 ) );
  OAI221_X1 U5693 ( .B1(\unit_memory/DRAM/n2565 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2821 ), .C2(n232), .A(\unit_memory/DRAM/n953 ), 
        .ZN(\unit_memory/DRAM/n952 ) );
  AOI22_X1 U5694 ( .A1(n154), .A2(\unit_memory/DRAM/n71 ), .B1(n167), .B2(
        \unit_memory/DRAM/n327 ), .ZN(\unit_memory/DRAM/n954 ) );
  OAI21_X1 U5695 ( .B1(\unit_memory/DRAM/n972 ), .B2(\unit_memory/DRAM/n973 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n965 ) );
  OAI221_X1 U5696 ( .B1(\unit_memory/DRAM/n2438 ), .B2(n194), .C1(
        \unit_memory/DRAM/n2694 ), .C2(n181), .A(\unit_memory/DRAM/n975 ), 
        .ZN(\unit_memory/DRAM/n972 ) );
  OAI221_X1 U5697 ( .B1(\unit_memory/DRAM/n2566 ), .B2(n246), .C1(
        \unit_memory/DRAM/n2822 ), .C2(n233), .A(\unit_memory/DRAM/n974 ), 
        .ZN(\unit_memory/DRAM/n973 ) );
  AOI22_X1 U5698 ( .A1(n155), .A2(\unit_memory/DRAM/n72 ), .B1(n168), .B2(
        \unit_memory/DRAM/n328 ), .ZN(\unit_memory/DRAM/n975 ) );
  OAI21_X1 U5699 ( .B1(\unit_memory/DRAM/n993 ), .B2(\unit_memory/DRAM/n994 ), 
        .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n986 ) );
  OAI221_X1 U5700 ( .B1(\unit_memory/DRAM/n2439 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2695 ), .C2(n179), .A(\unit_memory/DRAM/n996 ), 
        .ZN(\unit_memory/DRAM/n993 ) );
  OAI221_X1 U5701 ( .B1(\unit_memory/DRAM/n2567 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2823 ), .C2(n231), .A(\unit_memory/DRAM/n995 ), 
        .ZN(\unit_memory/DRAM/n994 ) );
  AOI22_X1 U5702 ( .A1(n153), .A2(\unit_memory/DRAM/n73 ), .B1(n166), .B2(
        \unit_memory/DRAM/n329 ), .ZN(\unit_memory/DRAM/n996 ) );
  OAI21_X1 U5703 ( .B1(\unit_memory/DRAM/n1014 ), .B2(\unit_memory/DRAM/n1015 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1007 ) );
  OAI221_X1 U5704 ( .B1(\unit_memory/DRAM/n2440 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2696 ), .C2(n179), .A(\unit_memory/DRAM/n1017 ), 
        .ZN(\unit_memory/DRAM/n1014 ) );
  OAI221_X1 U5705 ( .B1(\unit_memory/DRAM/n2568 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2824 ), .C2(n231), .A(\unit_memory/DRAM/n1016 ), 
        .ZN(\unit_memory/DRAM/n1015 ) );
  AOI22_X1 U5706 ( .A1(n153), .A2(\unit_memory/DRAM/n74 ), .B1(n166), .B2(
        \unit_memory/DRAM/n330 ), .ZN(\unit_memory/DRAM/n1017 ) );
  OAI21_X1 U5707 ( .B1(\unit_memory/DRAM/n1035 ), .B2(\unit_memory/DRAM/n1036 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1028 ) );
  OAI221_X1 U5708 ( .B1(\unit_memory/DRAM/n2441 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2697 ), .C2(n181), .A(\unit_memory/DRAM/n1038 ), 
        .ZN(\unit_memory/DRAM/n1035 ) );
  OAI221_X1 U5709 ( .B1(\unit_memory/DRAM/n2569 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2825 ), .C2(n233), .A(\unit_memory/DRAM/n1037 ), 
        .ZN(\unit_memory/DRAM/n1036 ) );
  AOI22_X1 U5710 ( .A1(n155), .A2(\unit_memory/DRAM/n75 ), .B1(n168), .B2(
        \unit_memory/DRAM/n331 ), .ZN(\unit_memory/DRAM/n1038 ) );
  OAI21_X1 U5711 ( .B1(\unit_memory/DRAM/n1056 ), .B2(\unit_memory/DRAM/n1057 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1049 ) );
  OAI221_X1 U5712 ( .B1(\unit_memory/DRAM/n2442 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2698 ), .C2(n179), .A(\unit_memory/DRAM/n1059 ), 
        .ZN(\unit_memory/DRAM/n1056 ) );
  OAI221_X1 U5713 ( .B1(\unit_memory/DRAM/n2570 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2826 ), .C2(n231), .A(\unit_memory/DRAM/n1058 ), 
        .ZN(\unit_memory/DRAM/n1057 ) );
  AOI22_X1 U5714 ( .A1(n153), .A2(\unit_memory/DRAM/n76 ), .B1(n166), .B2(
        \unit_memory/DRAM/n332 ), .ZN(\unit_memory/DRAM/n1059 ) );
  OAI21_X1 U5715 ( .B1(\unit_memory/DRAM/n1077 ), .B2(\unit_memory/DRAM/n1078 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1070 ) );
  OAI221_X1 U5716 ( .B1(\unit_memory/DRAM/n2443 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2699 ), .C2(n180), .A(\unit_memory/DRAM/n1080 ), 
        .ZN(\unit_memory/DRAM/n1077 ) );
  OAI221_X1 U5717 ( .B1(\unit_memory/DRAM/n2571 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2827 ), .C2(n232), .A(\unit_memory/DRAM/n1079 ), 
        .ZN(\unit_memory/DRAM/n1078 ) );
  AOI22_X1 U5718 ( .A1(n154), .A2(\unit_memory/DRAM/n77 ), .B1(n167), .B2(
        \unit_memory/DRAM/n333 ), .ZN(\unit_memory/DRAM/n1080 ) );
  OAI21_X1 U5719 ( .B1(\unit_memory/DRAM/n1098 ), .B2(\unit_memory/DRAM/n1099 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1091 ) );
  OAI221_X1 U5720 ( .B1(\unit_memory/DRAM/n2444 ), .B2(n193), .C1(
        \unit_memory/DRAM/n2700 ), .C2(n180), .A(\unit_memory/DRAM/n1101 ), 
        .ZN(\unit_memory/DRAM/n1098 ) );
  OAI221_X1 U5721 ( .B1(\unit_memory/DRAM/n2572 ), .B2(n245), .C1(
        \unit_memory/DRAM/n2828 ), .C2(n232), .A(\unit_memory/DRAM/n1100 ), 
        .ZN(\unit_memory/DRAM/n1099 ) );
  AOI22_X1 U5722 ( .A1(n154), .A2(\unit_memory/DRAM/n78 ), .B1(n167), .B2(
        \unit_memory/DRAM/n334 ), .ZN(\unit_memory/DRAM/n1101 ) );
  OAI21_X1 U5723 ( .B1(\unit_memory/DRAM/n1119 ), .B2(\unit_memory/DRAM/n1120 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1112 ) );
  OAI221_X1 U5724 ( .B1(\unit_memory/DRAM/n2445 ), .B2(n192), .C1(
        \unit_memory/DRAM/n2701 ), .C2(n179), .A(\unit_memory/DRAM/n1122 ), 
        .ZN(\unit_memory/DRAM/n1119 ) );
  OAI221_X1 U5725 ( .B1(\unit_memory/DRAM/n2573 ), .B2(n244), .C1(
        \unit_memory/DRAM/n2829 ), .C2(n231), .A(\unit_memory/DRAM/n1121 ), 
        .ZN(\unit_memory/DRAM/n1120 ) );
  AOI22_X1 U5726 ( .A1(n153), .A2(\unit_memory/DRAM/n79 ), .B1(n166), .B2(
        \unit_memory/DRAM/n335 ), .ZN(\unit_memory/DRAM/n1122 ) );
  OAI21_X1 U5727 ( .B1(\unit_memory/DRAM/n2187 ), .B2(\unit_memory/DRAM/n2188 ), .A(\unit_memory/DRAM/n824 ), .ZN(\unit_memory/DRAM/n1133 ) );
  OAI221_X1 U5728 ( .B1(\unit_memory/DRAM/n2446 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2702 ), .C2(n182), .A(\unit_memory/DRAM/n2190 ), 
        .ZN(\unit_memory/DRAM/n2187 ) );
  OAI221_X1 U5729 ( .B1(\unit_memory/DRAM/n2574 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2830 ), .C2(n234), .A(\unit_memory/DRAM/n2189 ), 
        .ZN(\unit_memory/DRAM/n2188 ) );
  AOI22_X1 U5730 ( .A1(n156), .A2(\unit_memory/DRAM/n80 ), .B1(n169), .B2(
        \unit_memory/DRAM/n336 ), .ZN(\unit_memory/DRAM/n2190 ) );
  AOI21_X1 U5731 ( .B1(\unit_memory/DRAM/n568 ), .B2(\unit_memory/DRAM/n569 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n567 ) );
  AOI221_X1 U5732 ( .B1(n202), .B2(\unit_memory/DRAM/n242 ), .C1(n215), .C2(
        \unit_memory/DRAM/n498 ), .A(\unit_memory/DRAM/n578 ), .ZN(
        \unit_memory/DRAM/n568 ) );
  AOI221_X1 U5733 ( .B1(n150), .B2(\unit_memory/DRAM/n114 ), .C1(n163), .C2(
        \unit_memory/DRAM/n370 ), .A(\unit_memory/DRAM/n573 ), .ZN(
        \unit_memory/DRAM/n569 ) );
  AOI21_X1 U5734 ( .B1(\unit_memory/DRAM/n599 ), .B2(\unit_memory/DRAM/n600 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n598 ) );
  AOI221_X1 U5735 ( .B1(n199), .B2(\unit_memory/DRAM/n243 ), .C1(n212), .C2(
        \unit_memory/DRAM/n499 ), .A(\unit_memory/DRAM/n602 ), .ZN(
        \unit_memory/DRAM/n599 ) );
  AOI221_X1 U5736 ( .B1(n147), .B2(\unit_memory/DRAM/n115 ), .C1(n160), .C2(
        \unit_memory/DRAM/n371 ), .A(\unit_memory/DRAM/n601 ), .ZN(
        \unit_memory/DRAM/n600 ) );
  AOI21_X1 U5737 ( .B1(\unit_memory/DRAM/n620 ), .B2(\unit_memory/DRAM/n621 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n619 ) );
  AOI221_X1 U5738 ( .B1(n199), .B2(\unit_memory/DRAM/n244 ), .C1(n212), .C2(
        \unit_memory/DRAM/n500 ), .A(\unit_memory/DRAM/n623 ), .ZN(
        \unit_memory/DRAM/n620 ) );
  AOI221_X1 U5739 ( .B1(n147), .B2(\unit_memory/DRAM/n116 ), .C1(n160), .C2(
        \unit_memory/DRAM/n372 ), .A(\unit_memory/DRAM/n622 ), .ZN(
        \unit_memory/DRAM/n621 ) );
  AOI21_X1 U5740 ( .B1(\unit_memory/DRAM/n641 ), .B2(\unit_memory/DRAM/n642 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n640 ) );
  AOI221_X1 U5741 ( .B1(n200), .B2(\unit_memory/DRAM/n245 ), .C1(n213), .C2(
        \unit_memory/DRAM/n501 ), .A(\unit_memory/DRAM/n644 ), .ZN(
        \unit_memory/DRAM/n641 ) );
  AOI221_X1 U5742 ( .B1(n148), .B2(\unit_memory/DRAM/n117 ), .C1(n161), .C2(
        \unit_memory/DRAM/n373 ), .A(\unit_memory/DRAM/n643 ), .ZN(
        \unit_memory/DRAM/n642 ) );
  AOI21_X1 U5743 ( .B1(\unit_memory/DRAM/n662 ), .B2(\unit_memory/DRAM/n663 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n661 ) );
  AOI221_X1 U5744 ( .B1(n200), .B2(\unit_memory/DRAM/n246 ), .C1(n213), .C2(
        \unit_memory/DRAM/n502 ), .A(\unit_memory/DRAM/n665 ), .ZN(
        \unit_memory/DRAM/n662 ) );
  AOI221_X1 U5745 ( .B1(n148), .B2(\unit_memory/DRAM/n118 ), .C1(n161), .C2(
        \unit_memory/DRAM/n374 ), .A(\unit_memory/DRAM/n664 ), .ZN(
        \unit_memory/DRAM/n663 ) );
  AOI21_X1 U5746 ( .B1(\unit_memory/DRAM/n683 ), .B2(\unit_memory/DRAM/n684 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n682 ) );
  AOI221_X1 U5747 ( .B1(n200), .B2(\unit_memory/DRAM/n247 ), .C1(n213), .C2(
        \unit_memory/DRAM/n503 ), .A(\unit_memory/DRAM/n686 ), .ZN(
        \unit_memory/DRAM/n683 ) );
  AOI221_X1 U5748 ( .B1(n148), .B2(\unit_memory/DRAM/n119 ), .C1(n161), .C2(
        \unit_memory/DRAM/n375 ), .A(\unit_memory/DRAM/n685 ), .ZN(
        \unit_memory/DRAM/n684 ) );
  AOI21_X1 U5749 ( .B1(\unit_memory/DRAM/n704 ), .B2(\unit_memory/DRAM/n705 ), 
        .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n703 ) );
  AOI221_X1 U5750 ( .B1(n201), .B2(\unit_memory/DRAM/n248 ), .C1(n214), .C2(
        \unit_memory/DRAM/n504 ), .A(\unit_memory/DRAM/n707 ), .ZN(
        \unit_memory/DRAM/n704 ) );
  AOI221_X1 U5751 ( .B1(n149), .B2(\unit_memory/DRAM/n120 ), .C1(n162), .C2(
        \unit_memory/DRAM/n376 ), .A(\unit_memory/DRAM/n706 ), .ZN(
        \unit_memory/DRAM/n705 ) );
  AOI21_X1 U5752 ( .B1(\unit_memory/DRAM/n2225 ), .B2(\unit_memory/DRAM/n2226 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2224 ) );
  AOI221_X1 U5753 ( .B1(n203), .B2(\unit_memory/DRAM/n250 ), .C1(n216), .C2(
        \unit_memory/DRAM/n506 ), .A(\unit_memory/DRAM/n2228 ), .ZN(
        \unit_memory/DRAM/n2225 ) );
  AOI221_X1 U5754 ( .B1(n151), .B2(\unit_memory/DRAM/n122 ), .C1(n164), .C2(
        \unit_memory/DRAM/n378 ), .A(\unit_memory/DRAM/n2227 ), .ZN(
        \unit_memory/DRAM/n2226 ) );
  AOI21_X1 U5755 ( .B1(\unit_memory/DRAM/n2246 ), .B2(\unit_memory/DRAM/n2247 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2245 ) );
  AOI221_X1 U5756 ( .B1(n204), .B2(\unit_memory/DRAM/n251 ), .C1(n217), .C2(
        \unit_memory/DRAM/n507 ), .A(\unit_memory/DRAM/n2249 ), .ZN(
        \unit_memory/DRAM/n2246 ) );
  AOI221_X1 U5757 ( .B1(n152), .B2(\unit_memory/DRAM/n123 ), .C1(n165), .C2(
        \unit_memory/DRAM/n379 ), .A(\unit_memory/DRAM/n2248 ), .ZN(
        \unit_memory/DRAM/n2247 ) );
  AOI21_X1 U5758 ( .B1(\unit_memory/DRAM/n2267 ), .B2(\unit_memory/DRAM/n2268 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2266 ) );
  AOI221_X1 U5759 ( .B1(n203), .B2(\unit_memory/DRAM/n252 ), .C1(n216), .C2(
        \unit_memory/DRAM/n508 ), .A(\unit_memory/DRAM/n2270 ), .ZN(
        \unit_memory/DRAM/n2267 ) );
  AOI221_X1 U5760 ( .B1(n151), .B2(\unit_memory/DRAM/n124 ), .C1(n164), .C2(
        \unit_memory/DRAM/n380 ), .A(\unit_memory/DRAM/n2269 ), .ZN(
        \unit_memory/DRAM/n2268 ) );
  AOI21_X1 U5761 ( .B1(\unit_memory/DRAM/n2288 ), .B2(\unit_memory/DRAM/n2289 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2287 ) );
  AOI221_X1 U5762 ( .B1(n203), .B2(\unit_memory/DRAM/n253 ), .C1(n216), .C2(
        \unit_memory/DRAM/n509 ), .A(\unit_memory/DRAM/n2291 ), .ZN(
        \unit_memory/DRAM/n2288 ) );
  AOI221_X1 U5763 ( .B1(n151), .B2(\unit_memory/DRAM/n125 ), .C1(n164), .C2(
        \unit_memory/DRAM/n381 ), .A(\unit_memory/DRAM/n2290 ), .ZN(
        \unit_memory/DRAM/n2289 ) );
  AOI21_X1 U5764 ( .B1(\unit_memory/DRAM/n2309 ), .B2(\unit_memory/DRAM/n2310 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2308 ) );
  AOI221_X1 U5765 ( .B1(n204), .B2(\unit_memory/DRAM/n254 ), .C1(n217), .C2(
        \unit_memory/DRAM/n510 ), .A(\unit_memory/DRAM/n2312 ), .ZN(
        \unit_memory/DRAM/n2309 ) );
  AOI221_X1 U5766 ( .B1(n152), .B2(\unit_memory/DRAM/n126 ), .C1(n165), .C2(
        \unit_memory/DRAM/n382 ), .A(\unit_memory/DRAM/n2311 ), .ZN(
        \unit_memory/DRAM/n2310 ) );
  AOI21_X1 U5767 ( .B1(\unit_memory/DRAM/n2330 ), .B2(\unit_memory/DRAM/n2331 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2329 ) );
  AOI221_X1 U5768 ( .B1(n203), .B2(\unit_memory/DRAM/n255 ), .C1(n216), .C2(
        \unit_memory/DRAM/n511 ), .A(\unit_memory/DRAM/n2333 ), .ZN(
        \unit_memory/DRAM/n2330 ) );
  AOI221_X1 U5769 ( .B1(n151), .B2(\unit_memory/DRAM/n127 ), .C1(n164), .C2(
        \unit_memory/DRAM/n383 ), .A(\unit_memory/DRAM/n2332 ), .ZN(
        \unit_memory/DRAM/n2331 ) );
  AOI21_X1 U5770 ( .B1(\unit_memory/DRAM/n2351 ), .B2(\unit_memory/DRAM/n2352 ), .A(\unit_memory/DRAM/n570 ), .ZN(\unit_memory/DRAM/n2350 ) );
  AOI221_X1 U5771 ( .B1(n204), .B2(\unit_memory/DRAM/n256 ), .C1(n217), .C2(
        \unit_memory/DRAM/n512 ), .A(\unit_memory/DRAM/n2354 ), .ZN(
        \unit_memory/DRAM/n2351 ) );
  AOI221_X1 U5772 ( .B1(n152), .B2(\unit_memory/DRAM/n128 ), .C1(n165), .C2(
        \unit_memory/DRAM/n384 ), .A(\unit_memory/DRAM/n2353 ), .ZN(
        \unit_memory/DRAM/n2352 ) );
  AOI21_X1 U5773 ( .B1(\unit_memory/DRAM/n581 ), .B2(\unit_memory/DRAM/n582 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n566 ) );
  AOI221_X1 U5774 ( .B1(n199), .B2(\unit_memory/DRAM/n210 ), .C1(n212), .C2(
        \unit_memory/DRAM/n466 ), .A(\unit_memory/DRAM/n585 ), .ZN(
        \unit_memory/DRAM/n581 ) );
  AOI221_X1 U5775 ( .B1(n147), .B2(\unit_memory/DRAM/n82 ), .C1(n160), .C2(
        \unit_memory/DRAM/n338 ), .A(\unit_memory/DRAM/n584 ), .ZN(
        \unit_memory/DRAM/n582 ) );
  AOI21_X1 U5776 ( .B1(\unit_memory/DRAM/n603 ), .B2(\unit_memory/DRAM/n604 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n597 ) );
  AOI221_X1 U5777 ( .B1(n199), .B2(\unit_memory/DRAM/n211 ), .C1(n212), .C2(
        \unit_memory/DRAM/n467 ), .A(\unit_memory/DRAM/n606 ), .ZN(
        \unit_memory/DRAM/n603 ) );
  AOI221_X1 U5778 ( .B1(n147), .B2(\unit_memory/DRAM/n83 ), .C1(n160), .C2(
        \unit_memory/DRAM/n339 ), .A(\unit_memory/DRAM/n605 ), .ZN(
        \unit_memory/DRAM/n604 ) );
  AOI21_X1 U5779 ( .B1(\unit_memory/DRAM/n624 ), .B2(\unit_memory/DRAM/n625 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n618 ) );
  AOI221_X1 U5780 ( .B1(n199), .B2(\unit_memory/DRAM/n212 ), .C1(n212), .C2(
        \unit_memory/DRAM/n468 ), .A(\unit_memory/DRAM/n627 ), .ZN(
        \unit_memory/DRAM/n624 ) );
  AOI221_X1 U5781 ( .B1(n147), .B2(\unit_memory/DRAM/n84 ), .C1(n160), .C2(
        \unit_memory/DRAM/n340 ), .A(\unit_memory/DRAM/n626 ), .ZN(
        \unit_memory/DRAM/n625 ) );
  AOI21_X1 U5782 ( .B1(\unit_memory/DRAM/n645 ), .B2(\unit_memory/DRAM/n646 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n639 ) );
  AOI221_X1 U5783 ( .B1(n200), .B2(\unit_memory/DRAM/n213 ), .C1(n213), .C2(
        \unit_memory/DRAM/n469 ), .A(\unit_memory/DRAM/n648 ), .ZN(
        \unit_memory/DRAM/n645 ) );
  AOI221_X1 U5784 ( .B1(n148), .B2(\unit_memory/DRAM/n85 ), .C1(n161), .C2(
        \unit_memory/DRAM/n341 ), .A(\unit_memory/DRAM/n647 ), .ZN(
        \unit_memory/DRAM/n646 ) );
  AOI21_X1 U5785 ( .B1(\unit_memory/DRAM/n666 ), .B2(\unit_memory/DRAM/n667 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n660 ) );
  AOI221_X1 U5786 ( .B1(n200), .B2(\unit_memory/DRAM/n214 ), .C1(n213), .C2(
        \unit_memory/DRAM/n470 ), .A(\unit_memory/DRAM/n669 ), .ZN(
        \unit_memory/DRAM/n666 ) );
  AOI221_X1 U5787 ( .B1(n148), .B2(\unit_memory/DRAM/n86 ), .C1(n161), .C2(
        \unit_memory/DRAM/n342 ), .A(\unit_memory/DRAM/n668 ), .ZN(
        \unit_memory/DRAM/n667 ) );
  AOI21_X1 U5788 ( .B1(\unit_memory/DRAM/n687 ), .B2(\unit_memory/DRAM/n688 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n681 ) );
  AOI221_X1 U5789 ( .B1(n200), .B2(\unit_memory/DRAM/n215 ), .C1(n213), .C2(
        \unit_memory/DRAM/n471 ), .A(\unit_memory/DRAM/n690 ), .ZN(
        \unit_memory/DRAM/n687 ) );
  AOI221_X1 U5790 ( .B1(n148), .B2(\unit_memory/DRAM/n87 ), .C1(n161), .C2(
        \unit_memory/DRAM/n343 ), .A(\unit_memory/DRAM/n689 ), .ZN(
        \unit_memory/DRAM/n688 ) );
  AOI21_X1 U5791 ( .B1(\unit_memory/DRAM/n708 ), .B2(\unit_memory/DRAM/n709 ), 
        .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n702 ) );
  AOI221_X1 U5792 ( .B1(n201), .B2(\unit_memory/DRAM/n216 ), .C1(n214), .C2(
        \unit_memory/DRAM/n472 ), .A(\unit_memory/DRAM/n711 ), .ZN(
        \unit_memory/DRAM/n708 ) );
  AOI221_X1 U5793 ( .B1(n149), .B2(\unit_memory/DRAM/n88 ), .C1(n162), .C2(
        \unit_memory/DRAM/n344 ), .A(\unit_memory/DRAM/n710 ), .ZN(
        \unit_memory/DRAM/n709 ) );
  AOI21_X1 U5794 ( .B1(\unit_memory/DRAM/n2229 ), .B2(\unit_memory/DRAM/n2230 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2223 ) );
  AOI221_X1 U5795 ( .B1(n203), .B2(\unit_memory/DRAM/n218 ), .C1(n216), .C2(
        \unit_memory/DRAM/n474 ), .A(\unit_memory/DRAM/n2232 ), .ZN(
        \unit_memory/DRAM/n2229 ) );
  AOI221_X1 U5796 ( .B1(n151), .B2(\unit_memory/DRAM/n90 ), .C1(n164), .C2(
        \unit_memory/DRAM/n346 ), .A(\unit_memory/DRAM/n2231 ), .ZN(
        \unit_memory/DRAM/n2230 ) );
  AOI21_X1 U5797 ( .B1(\unit_memory/DRAM/n2250 ), .B2(\unit_memory/DRAM/n2251 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2244 ) );
  AOI221_X1 U5798 ( .B1(n202), .B2(\unit_memory/DRAM/n219 ), .C1(n215), .C2(
        \unit_memory/DRAM/n475 ), .A(\unit_memory/DRAM/n2253 ), .ZN(
        \unit_memory/DRAM/n2250 ) );
  AOI221_X1 U5799 ( .B1(n150), .B2(\unit_memory/DRAM/n91 ), .C1(n163), .C2(
        \unit_memory/DRAM/n347 ), .A(\unit_memory/DRAM/n2252 ), .ZN(
        \unit_memory/DRAM/n2251 ) );
  AOI21_X1 U5800 ( .B1(\unit_memory/DRAM/n2271 ), .B2(\unit_memory/DRAM/n2272 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2265 ) );
  AOI221_X1 U5801 ( .B1(n203), .B2(\unit_memory/DRAM/n220 ), .C1(n216), .C2(
        \unit_memory/DRAM/n476 ), .A(\unit_memory/DRAM/n2274 ), .ZN(
        \unit_memory/DRAM/n2271 ) );
  AOI221_X1 U5802 ( .B1(n151), .B2(\unit_memory/DRAM/n92 ), .C1(n164), .C2(
        \unit_memory/DRAM/n348 ), .A(\unit_memory/DRAM/n2273 ), .ZN(
        \unit_memory/DRAM/n2272 ) );
  AOI21_X1 U5803 ( .B1(\unit_memory/DRAM/n2292 ), .B2(\unit_memory/DRAM/n2293 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2286 ) );
  AOI221_X1 U5804 ( .B1(n204), .B2(\unit_memory/DRAM/n221 ), .C1(n217), .C2(
        \unit_memory/DRAM/n477 ), .A(\unit_memory/DRAM/n2295 ), .ZN(
        \unit_memory/DRAM/n2292 ) );
  AOI221_X1 U5805 ( .B1(n152), .B2(\unit_memory/DRAM/n93 ), .C1(n165), .C2(
        \unit_memory/DRAM/n349 ), .A(\unit_memory/DRAM/n2294 ), .ZN(
        \unit_memory/DRAM/n2293 ) );
  AOI21_X1 U5806 ( .B1(\unit_memory/DRAM/n2313 ), .B2(\unit_memory/DRAM/n2314 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2307 ) );
  AOI221_X1 U5807 ( .B1(n203), .B2(\unit_memory/DRAM/n222 ), .C1(n216), .C2(
        \unit_memory/DRAM/n478 ), .A(\unit_memory/DRAM/n2316 ), .ZN(
        \unit_memory/DRAM/n2313 ) );
  AOI221_X1 U5808 ( .B1(n151), .B2(\unit_memory/DRAM/n94 ), .C1(n164), .C2(
        \unit_memory/DRAM/n350 ), .A(\unit_memory/DRAM/n2315 ), .ZN(
        \unit_memory/DRAM/n2314 ) );
  AOI21_X1 U5809 ( .B1(\unit_memory/DRAM/n2334 ), .B2(\unit_memory/DRAM/n2335 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2328 ) );
  AOI221_X1 U5810 ( .B1(n204), .B2(\unit_memory/DRAM/n223 ), .C1(n217), .C2(
        \unit_memory/DRAM/n479 ), .A(\unit_memory/DRAM/n2337 ), .ZN(
        \unit_memory/DRAM/n2334 ) );
  AOI221_X1 U5811 ( .B1(n152), .B2(\unit_memory/DRAM/n95 ), .C1(n165), .C2(
        \unit_memory/DRAM/n351 ), .A(\unit_memory/DRAM/n2336 ), .ZN(
        \unit_memory/DRAM/n2335 ) );
  AOI21_X1 U5812 ( .B1(\unit_memory/DRAM/n2355 ), .B2(\unit_memory/DRAM/n2356 ), .A(\unit_memory/DRAM/n583 ), .ZN(\unit_memory/DRAM/n2349 ) );
  AOI221_X1 U5813 ( .B1(n204), .B2(\unit_memory/DRAM/n224 ), .C1(n217), .C2(
        \unit_memory/DRAM/n480 ), .A(\unit_memory/DRAM/n2358 ), .ZN(
        \unit_memory/DRAM/n2355 ) );
  AOI221_X1 U5814 ( .B1(n152), .B2(\unit_memory/DRAM/n96 ), .C1(n165), .C2(
        \unit_memory/DRAM/n352 ), .A(\unit_memory/DRAM/n2357 ), .ZN(
        \unit_memory/DRAM/n2356 ) );
  OAI21_X1 U5815 ( .B1(\unit_memory/DRAM/n2204 ), .B2(\unit_memory/DRAM/n2205 ), .A(\unit_memory/DRAM/n1143 ), .ZN(\unit_memory/DRAM/n2203 ) );
  OAI221_X1 U5816 ( .B1(\unit_memory/DRAM/n2391 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2647 ), .C2(n183), .A(\unit_memory/DRAM/n2207 ), 
        .ZN(\unit_memory/DRAM/n2204 ) );
  OAI221_X1 U5817 ( .B1(\unit_memory/DRAM/n2519 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2775 ), .C2(n235), .A(\unit_memory/DRAM/n2206 ), 
        .ZN(\unit_memory/DRAM/n2205 ) );
  AOI22_X1 U5818 ( .A1(n157), .A2(\unit_memory/DRAM/n25 ), .B1(n170), .B2(
        \unit_memory/DRAM/n281 ), .ZN(\unit_memory/DRAM/n2207 ) );
  OAI21_X1 U5819 ( .B1(\unit_memory/DRAM/n2212 ), .B2(\unit_memory/DRAM/n2213 ), .A(\unit_memory/DRAM/n549 ), .ZN(\unit_memory/DRAM/n2201 ) );
  OAI221_X1 U5820 ( .B1(\unit_memory/DRAM/n2455 ), .B2(n196), .C1(
        \unit_memory/DRAM/n2711 ), .C2(n183), .A(\unit_memory/DRAM/n2215 ), 
        .ZN(\unit_memory/DRAM/n2212 ) );
  OAI221_X1 U5821 ( .B1(\unit_memory/DRAM/n2583 ), .B2(n248), .C1(
        \unit_memory/DRAM/n2839 ), .C2(n235), .A(\unit_memory/DRAM/n2214 ), 
        .ZN(\unit_memory/DRAM/n2213 ) );
  AOI22_X1 U5822 ( .A1(n157), .A2(\unit_memory/DRAM/n89 ), .B1(n170), .B2(
        \unit_memory/DRAM/n345 ), .ZN(\unit_memory/DRAM/n2215 ) );
  NAND2_X1 U5823 ( .A1(aluout_regn[2]), .A2(\unit_memory/DRAM/n782 ), .ZN(
        \unit_memory/DRAM/n579 ) );
  NAND2_X1 U5824 ( .A1(aluout_regn[2]), .A2(\unit_memory/DRAM/n772 ), .ZN(
        \unit_memory/DRAM/n580 ) );
  OAI21_X1 U5825 ( .B1(\unit_memory/DRAM/n1141 ), .B2(\unit_memory/DRAM/n1142 ), .A(\unit_memory/DRAM/n1143 ), .ZN(\unit_memory/DRAM/n1140 ) );
  OAI221_X1 U5826 ( .B1(\unit_memory/DRAM/n2383 ), .B2(n195), .C1(
        \unit_memory/DRAM/n2639 ), .C2(n182), .A(\unit_memory/DRAM/n1145 ), 
        .ZN(\unit_memory/DRAM/n1141 ) );
  OAI221_X1 U5827 ( .B1(\unit_memory/DRAM/n2511 ), .B2(n247), .C1(
        \unit_memory/DRAM/n2767 ), .C2(n234), .A(\unit_memory/DRAM/n1144 ), 
        .ZN(\unit_memory/DRAM/n1142 ) );
  AOI22_X1 U5828 ( .A1(n156), .A2(\unit_memory/DRAM/n17 ), .B1(n169), .B2(
        \unit_memory/DRAM/n273 ), .ZN(\unit_memory/DRAM/n1145 ) );
  NOR4_X1 U5829 ( .A1(\unit_memory/DRAM/n564 ), .A2(\unit_memory/DRAM/n565 ), 
        .A3(\unit_memory/DRAM/n566 ), .A4(\unit_memory/DRAM/n567 ), .ZN(
        \unit_memory/DRAM/n563 ) );
  AOI21_X1 U5830 ( .B1(\unit_memory/DRAM/n590 ), .B2(\unit_memory/DRAM/n591 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n564 ) );
  AOI21_X1 U5831 ( .B1(\unit_memory/DRAM/n586 ), .B2(\unit_memory/DRAM/n587 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n565 ) );
  NOR4_X1 U5832 ( .A1(\unit_memory/DRAM/n595 ), .A2(\unit_memory/DRAM/n596 ), 
        .A3(\unit_memory/DRAM/n597 ), .A4(\unit_memory/DRAM/n598 ), .ZN(
        \unit_memory/DRAM/n594 ) );
  AOI21_X1 U5833 ( .B1(\unit_memory/DRAM/n611 ), .B2(\unit_memory/DRAM/n612 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n595 ) );
  AOI21_X1 U5834 ( .B1(\unit_memory/DRAM/n607 ), .B2(\unit_memory/DRAM/n608 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n596 ) );
  NOR4_X1 U5835 ( .A1(\unit_memory/DRAM/n616 ), .A2(\unit_memory/DRAM/n617 ), 
        .A3(\unit_memory/DRAM/n618 ), .A4(\unit_memory/DRAM/n619 ), .ZN(
        \unit_memory/DRAM/n615 ) );
  AOI21_X1 U5836 ( .B1(\unit_memory/DRAM/n632 ), .B2(\unit_memory/DRAM/n633 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n616 ) );
  AOI21_X1 U5837 ( .B1(\unit_memory/DRAM/n628 ), .B2(\unit_memory/DRAM/n629 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n617 ) );
  NOR4_X1 U5838 ( .A1(\unit_memory/DRAM/n637 ), .A2(\unit_memory/DRAM/n638 ), 
        .A3(\unit_memory/DRAM/n639 ), .A4(\unit_memory/DRAM/n640 ), .ZN(
        \unit_memory/DRAM/n636 ) );
  AOI21_X1 U5839 ( .B1(\unit_memory/DRAM/n653 ), .B2(\unit_memory/DRAM/n654 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n637 ) );
  AOI21_X1 U5840 ( .B1(\unit_memory/DRAM/n649 ), .B2(\unit_memory/DRAM/n650 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n638 ) );
  NOR4_X1 U5841 ( .A1(\unit_memory/DRAM/n658 ), .A2(\unit_memory/DRAM/n659 ), 
        .A3(\unit_memory/DRAM/n660 ), .A4(\unit_memory/DRAM/n661 ), .ZN(
        \unit_memory/DRAM/n657 ) );
  AOI21_X1 U5842 ( .B1(\unit_memory/DRAM/n674 ), .B2(\unit_memory/DRAM/n675 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n658 ) );
  AOI21_X1 U5843 ( .B1(\unit_memory/DRAM/n670 ), .B2(\unit_memory/DRAM/n671 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n659 ) );
  NOR4_X1 U5844 ( .A1(\unit_memory/DRAM/n679 ), .A2(\unit_memory/DRAM/n680 ), 
        .A3(\unit_memory/DRAM/n681 ), .A4(\unit_memory/DRAM/n682 ), .ZN(
        \unit_memory/DRAM/n678 ) );
  AOI21_X1 U5845 ( .B1(\unit_memory/DRAM/n695 ), .B2(\unit_memory/DRAM/n696 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n679 ) );
  AOI21_X1 U5846 ( .B1(\unit_memory/DRAM/n691 ), .B2(\unit_memory/DRAM/n692 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n680 ) );
  NOR4_X1 U5847 ( .A1(\unit_memory/DRAM/n700 ), .A2(\unit_memory/DRAM/n701 ), 
        .A3(\unit_memory/DRAM/n702 ), .A4(\unit_memory/DRAM/n703 ), .ZN(
        \unit_memory/DRAM/n699 ) );
  AOI21_X1 U5848 ( .B1(\unit_memory/DRAM/n716 ), .B2(\unit_memory/DRAM/n717 ), 
        .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n700 ) );
  AOI21_X1 U5849 ( .B1(\unit_memory/DRAM/n712 ), .B2(\unit_memory/DRAM/n713 ), 
        .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n701 ) );
  NAND2_X1 U5850 ( .A1(\unit_decode/n2430 ), .A2(\unit_decode/n2431 ), .ZN(
        \unit_decode/RegisterFile/N436 ) );
  NOR4_X1 U5851 ( .A1(\unit_decode/n2440 ), .A2(\unit_decode/n2441 ), .A3(
        \unit_decode/n2442 ), .A4(\unit_decode/n2443 ), .ZN(
        \unit_decode/n2430 ) );
  NOR4_X1 U5852 ( .A1(\unit_decode/n2432 ), .A2(\unit_decode/n2433 ), .A3(
        \unit_decode/n2434 ), .A4(\unit_decode/n2435 ), .ZN(
        \unit_decode/n2431 ) );
  OAI221_X1 U5853 ( .B1(\unit_decode/RegisterFile/n3811 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3843 ), .C2(n1182), .A(\unit_decode/n2447 ), 
        .ZN(\unit_decode/n2440 ) );
  NAND2_X1 U5854 ( .A1(\unit_decode/n2412 ), .A2(\unit_decode/n2413 ), .ZN(
        \unit_decode/RegisterFile/N437 ) );
  NOR4_X1 U5855 ( .A1(\unit_decode/n2422 ), .A2(\unit_decode/n2423 ), .A3(
        \unit_decode/n2424 ), .A4(\unit_decode/n2425 ), .ZN(
        \unit_decode/n2412 ) );
  NOR4_X1 U5856 ( .A1(\unit_decode/n2414 ), .A2(\unit_decode/n2415 ), .A3(
        \unit_decode/n2416 ), .A4(\unit_decode/n2417 ), .ZN(
        \unit_decode/n2413 ) );
  OAI221_X1 U5857 ( .B1(\unit_decode/RegisterFile/n3810 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3842 ), .C2(n1182), .A(\unit_decode/n2429 ), 
        .ZN(\unit_decode/n2422 ) );
  NAND2_X1 U5858 ( .A1(\unit_decode/n2394 ), .A2(\unit_decode/n2395 ), .ZN(
        \unit_decode/RegisterFile/N438 ) );
  NOR4_X1 U5859 ( .A1(\unit_decode/n2404 ), .A2(\unit_decode/n2405 ), .A3(
        \unit_decode/n2406 ), .A4(\unit_decode/n2407 ), .ZN(
        \unit_decode/n2394 ) );
  NOR4_X1 U5860 ( .A1(\unit_decode/n2396 ), .A2(\unit_decode/n2397 ), .A3(
        \unit_decode/n2398 ), .A4(\unit_decode/n2399 ), .ZN(
        \unit_decode/n2395 ) );
  OAI221_X1 U5861 ( .B1(\unit_decode/RegisterFile/n3809 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3841 ), .C2(n1182), .A(\unit_decode/n2411 ), 
        .ZN(\unit_decode/n2404 ) );
  NAND2_X1 U5862 ( .A1(\unit_decode/n2376 ), .A2(\unit_decode/n2377 ), .ZN(
        \unit_decode/RegisterFile/N439 ) );
  NOR4_X1 U5863 ( .A1(\unit_decode/n2386 ), .A2(\unit_decode/n2387 ), .A3(
        \unit_decode/n2388 ), .A4(\unit_decode/n2389 ), .ZN(
        \unit_decode/n2376 ) );
  NOR4_X1 U5864 ( .A1(\unit_decode/n2378 ), .A2(\unit_decode/n2379 ), .A3(
        \unit_decode/n2380 ), .A4(\unit_decode/n2381 ), .ZN(
        \unit_decode/n2377 ) );
  OAI221_X1 U5865 ( .B1(\unit_decode/RegisterFile/n3808 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3840 ), .C2(n1182), .A(\unit_decode/n2393 ), 
        .ZN(\unit_decode/n2386 ) );
  NAND2_X1 U5866 ( .A1(\unit_decode/n2358 ), .A2(\unit_decode/n2359 ), .ZN(
        \unit_decode/RegisterFile/N440 ) );
  NOR4_X1 U5867 ( .A1(\unit_decode/n2368 ), .A2(\unit_decode/n2369 ), .A3(
        \unit_decode/n2370 ), .A4(\unit_decode/n2371 ), .ZN(
        \unit_decode/n2358 ) );
  NOR4_X1 U5868 ( .A1(\unit_decode/n2360 ), .A2(\unit_decode/n2361 ), .A3(
        \unit_decode/n2362 ), .A4(\unit_decode/n2363 ), .ZN(
        \unit_decode/n2359 ) );
  OAI221_X1 U5869 ( .B1(\unit_decode/RegisterFile/n3807 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3839 ), .C2(n1182), .A(\unit_decode/n2375 ), 
        .ZN(\unit_decode/n2368 ) );
  NAND2_X1 U5870 ( .A1(\unit_decode/n2340 ), .A2(\unit_decode/n2341 ), .ZN(
        \unit_decode/RegisterFile/N441 ) );
  NOR4_X1 U5871 ( .A1(\unit_decode/n2350 ), .A2(\unit_decode/n2351 ), .A3(
        \unit_decode/n2352 ), .A4(\unit_decode/n2353 ), .ZN(
        \unit_decode/n2340 ) );
  NOR4_X1 U5872 ( .A1(\unit_decode/n2342 ), .A2(\unit_decode/n2343 ), .A3(
        \unit_decode/n2344 ), .A4(\unit_decode/n2345 ), .ZN(
        \unit_decode/n2341 ) );
  OAI221_X1 U5873 ( .B1(\unit_decode/RegisterFile/n3806 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3838 ), .C2(n1182), .A(\unit_decode/n2357 ), 
        .ZN(\unit_decode/n2350 ) );
  NAND2_X1 U5874 ( .A1(\unit_decode/n2322 ), .A2(\unit_decode/n2323 ), .ZN(
        \unit_decode/RegisterFile/N442 ) );
  NOR4_X1 U5875 ( .A1(\unit_decode/n2332 ), .A2(\unit_decode/n2333 ), .A3(
        \unit_decode/n2334 ), .A4(\unit_decode/n2335 ), .ZN(
        \unit_decode/n2322 ) );
  NOR4_X1 U5876 ( .A1(\unit_decode/n2324 ), .A2(\unit_decode/n2325 ), .A3(
        \unit_decode/n2326 ), .A4(\unit_decode/n2327 ), .ZN(
        \unit_decode/n2323 ) );
  OAI221_X1 U5877 ( .B1(\unit_decode/RegisterFile/n3805 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3837 ), .C2(n1182), .A(\unit_decode/n2339 ), 
        .ZN(\unit_decode/n2332 ) );
  NAND2_X1 U5878 ( .A1(\unit_decode/n2272 ), .A2(\unit_decode/n2273 ), .ZN(
        \unit_decode/RegisterFile/N443 ) );
  NOR4_X1 U5879 ( .A1(\unit_decode/n2298 ), .A2(\unit_decode/n2299 ), .A3(
        \unit_decode/n2300 ), .A4(\unit_decode/n2301 ), .ZN(
        \unit_decode/n2272 ) );
  NOR4_X1 U5880 ( .A1(\unit_decode/n2274 ), .A2(\unit_decode/n2275 ), .A3(
        \unit_decode/n2276 ), .A4(\unit_decode/n2277 ), .ZN(
        \unit_decode/n2273 ) );
  OAI221_X1 U5881 ( .B1(\unit_decode/RegisterFile/n3804 ), .B2(n1179), .C1(
        \unit_decode/RegisterFile/n3836 ), .C2(n1182), .A(\unit_decode/n2319 ), 
        .ZN(\unit_decode/n2298 ) );
  NAND2_X1 U5882 ( .A1(\unit_decode/n3050 ), .A2(\unit_decode/n3051 ), .ZN(
        \unit_decode/RegisterFile/N403 ) );
  NOR4_X1 U5883 ( .A1(\unit_decode/n3060 ), .A2(\unit_decode/n3061 ), .A3(
        \unit_decode/n3062 ), .A4(\unit_decode/n3063 ), .ZN(
        \unit_decode/n3050 ) );
  NOR4_X1 U5884 ( .A1(\unit_decode/n3052 ), .A2(\unit_decode/n3053 ), .A3(
        \unit_decode/n3054 ), .A4(\unit_decode/n3055 ), .ZN(
        \unit_decode/n3051 ) );
  OAI221_X1 U5885 ( .B1(\unit_decode/RegisterFile/n3811 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3843 ), .C2(n1278), .A(\unit_decode/n3067 ), 
        .ZN(\unit_decode/n3060 ) );
  NAND2_X1 U5886 ( .A1(\unit_decode/n3032 ), .A2(\unit_decode/n3033 ), .ZN(
        \unit_decode/RegisterFile/N404 ) );
  NOR4_X1 U5887 ( .A1(\unit_decode/n3042 ), .A2(\unit_decode/n3043 ), .A3(
        \unit_decode/n3044 ), .A4(\unit_decode/n3045 ), .ZN(
        \unit_decode/n3032 ) );
  NOR4_X1 U5888 ( .A1(\unit_decode/n3034 ), .A2(\unit_decode/n3035 ), .A3(
        \unit_decode/n3036 ), .A4(\unit_decode/n3037 ), .ZN(
        \unit_decode/n3033 ) );
  OAI221_X1 U5889 ( .B1(\unit_decode/RegisterFile/n3810 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3842 ), .C2(n1278), .A(\unit_decode/n3049 ), 
        .ZN(\unit_decode/n3042 ) );
  NAND2_X1 U5890 ( .A1(\unit_decode/n3014 ), .A2(\unit_decode/n3015 ), .ZN(
        \unit_decode/RegisterFile/N405 ) );
  NOR4_X1 U5891 ( .A1(\unit_decode/n3024 ), .A2(\unit_decode/n3025 ), .A3(
        \unit_decode/n3026 ), .A4(\unit_decode/n3027 ), .ZN(
        \unit_decode/n3014 ) );
  NOR4_X1 U5892 ( .A1(\unit_decode/n3016 ), .A2(\unit_decode/n3017 ), .A3(
        \unit_decode/n3018 ), .A4(\unit_decode/n3019 ), .ZN(
        \unit_decode/n3015 ) );
  OAI221_X1 U5893 ( .B1(\unit_decode/RegisterFile/n3809 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3841 ), .C2(n1278), .A(\unit_decode/n3031 ), 
        .ZN(\unit_decode/n3024 ) );
  NAND2_X1 U5894 ( .A1(\unit_decode/n2996 ), .A2(\unit_decode/n2997 ), .ZN(
        \unit_decode/RegisterFile/N406 ) );
  NOR4_X1 U5895 ( .A1(\unit_decode/n3006 ), .A2(\unit_decode/n3007 ), .A3(
        \unit_decode/n3008 ), .A4(\unit_decode/n3009 ), .ZN(
        \unit_decode/n2996 ) );
  NOR4_X1 U5896 ( .A1(\unit_decode/n2998 ), .A2(\unit_decode/n2999 ), .A3(
        \unit_decode/n3000 ), .A4(\unit_decode/n3001 ), .ZN(
        \unit_decode/n2997 ) );
  OAI221_X1 U5897 ( .B1(\unit_decode/RegisterFile/n3808 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3840 ), .C2(n1278), .A(\unit_decode/n3013 ), 
        .ZN(\unit_decode/n3006 ) );
  NAND2_X1 U5898 ( .A1(\unit_decode/n2978 ), .A2(\unit_decode/n2979 ), .ZN(
        \unit_decode/RegisterFile/N407 ) );
  NOR4_X1 U5899 ( .A1(\unit_decode/n2988 ), .A2(\unit_decode/n2989 ), .A3(
        \unit_decode/n2990 ), .A4(\unit_decode/n2991 ), .ZN(
        \unit_decode/n2978 ) );
  NOR4_X1 U5900 ( .A1(\unit_decode/n2980 ), .A2(\unit_decode/n2981 ), .A3(
        \unit_decode/n2982 ), .A4(\unit_decode/n2983 ), .ZN(
        \unit_decode/n2979 ) );
  OAI221_X1 U5901 ( .B1(\unit_decode/RegisterFile/n3807 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3839 ), .C2(n1278), .A(\unit_decode/n2995 ), 
        .ZN(\unit_decode/n2988 ) );
  NAND2_X1 U5902 ( .A1(\unit_decode/n2960 ), .A2(\unit_decode/n2961 ), .ZN(
        \unit_decode/RegisterFile/N408 ) );
  NOR4_X1 U5903 ( .A1(\unit_decode/n2970 ), .A2(\unit_decode/n2971 ), .A3(
        \unit_decode/n2972 ), .A4(\unit_decode/n2973 ), .ZN(
        \unit_decode/n2960 ) );
  NOR4_X1 U5904 ( .A1(\unit_decode/n2962 ), .A2(\unit_decode/n2963 ), .A3(
        \unit_decode/n2964 ), .A4(\unit_decode/n2965 ), .ZN(
        \unit_decode/n2961 ) );
  OAI221_X1 U5905 ( .B1(\unit_decode/RegisterFile/n3806 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3838 ), .C2(n1278), .A(\unit_decode/n2977 ), 
        .ZN(\unit_decode/n2970 ) );
  NAND2_X1 U5906 ( .A1(\unit_decode/n2942 ), .A2(\unit_decode/n2943 ), .ZN(
        \unit_decode/RegisterFile/N409 ) );
  NOR4_X1 U5907 ( .A1(\unit_decode/n2952 ), .A2(\unit_decode/n2953 ), .A3(
        \unit_decode/n2954 ), .A4(\unit_decode/n2955 ), .ZN(
        \unit_decode/n2942 ) );
  NOR4_X1 U5908 ( .A1(\unit_decode/n2944 ), .A2(\unit_decode/n2945 ), .A3(
        \unit_decode/n2946 ), .A4(\unit_decode/n2947 ), .ZN(
        \unit_decode/n2943 ) );
  OAI221_X1 U5909 ( .B1(\unit_decode/RegisterFile/n3805 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3837 ), .C2(n1278), .A(\unit_decode/n2959 ), 
        .ZN(\unit_decode/n2952 ) );
  NAND2_X1 U5910 ( .A1(\unit_decode/n2892 ), .A2(\unit_decode/n2893 ), .ZN(
        \unit_decode/RegisterFile/N410 ) );
  NOR4_X1 U5911 ( .A1(\unit_decode/n2918 ), .A2(\unit_decode/n2919 ), .A3(
        \unit_decode/n2920 ), .A4(\unit_decode/n2921 ), .ZN(
        \unit_decode/n2892 ) );
  NOR4_X1 U5912 ( .A1(\unit_decode/n2894 ), .A2(\unit_decode/n2895 ), .A3(
        \unit_decode/n2896 ), .A4(\unit_decode/n2897 ), .ZN(
        \unit_decode/n2893 ) );
  OAI221_X1 U5913 ( .B1(\unit_decode/RegisterFile/n3804 ), .B2(n1275), .C1(
        \unit_decode/RegisterFile/n3836 ), .C2(n1278), .A(\unit_decode/n2939 ), 
        .ZN(\unit_decode/n2918 ) );
  AND2_X1 U5914 ( .A1(aluout_regn[2]), .A2(\unit_memory/DRAM/n792 ), .ZN(
        \unit_memory/DRAM/n576 ) );
  AND2_X1 U5915 ( .A1(aluout_regn[2]), .A2(\unit_memory/DRAM/n809 ), .ZN(
        \unit_memory/DRAM/n577 ) );
  NOR4_X1 U5916 ( .A1(\unit_memory/DRAM/n2221 ), .A2(\unit_memory/DRAM/n2222 ), 
        .A3(\unit_memory/DRAM/n2223 ), .A4(\unit_memory/DRAM/n2224 ), .ZN(
        \unit_memory/DRAM/n2220 ) );
  AOI21_X1 U5917 ( .B1(\unit_memory/DRAM/n2237 ), .B2(\unit_memory/DRAM/n2238 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2221 ) );
  AOI21_X1 U5918 ( .B1(\unit_memory/DRAM/n2233 ), .B2(\unit_memory/DRAM/n2234 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2222 ) );
  NOR4_X1 U5919 ( .A1(\unit_memory/DRAM/n2242 ), .A2(\unit_memory/DRAM/n2243 ), 
        .A3(\unit_memory/DRAM/n2244 ), .A4(\unit_memory/DRAM/n2245 ), .ZN(
        \unit_memory/DRAM/n2241 ) );
  AOI21_X1 U5920 ( .B1(\unit_memory/DRAM/n2258 ), .B2(\unit_memory/DRAM/n2259 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2242 ) );
  AOI21_X1 U5921 ( .B1(\unit_memory/DRAM/n2254 ), .B2(\unit_memory/DRAM/n2255 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2243 ) );
  NOR4_X1 U5922 ( .A1(\unit_memory/DRAM/n2263 ), .A2(\unit_memory/DRAM/n2264 ), 
        .A3(\unit_memory/DRAM/n2265 ), .A4(\unit_memory/DRAM/n2266 ), .ZN(
        \unit_memory/DRAM/n2262 ) );
  AOI21_X1 U5923 ( .B1(\unit_memory/DRAM/n2279 ), .B2(\unit_memory/DRAM/n2280 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2263 ) );
  AOI21_X1 U5924 ( .B1(\unit_memory/DRAM/n2275 ), .B2(\unit_memory/DRAM/n2276 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2264 ) );
  NOR4_X1 U5925 ( .A1(\unit_memory/DRAM/n2284 ), .A2(\unit_memory/DRAM/n2285 ), 
        .A3(\unit_memory/DRAM/n2286 ), .A4(\unit_memory/DRAM/n2287 ), .ZN(
        \unit_memory/DRAM/n2283 ) );
  AOI21_X1 U5926 ( .B1(\unit_memory/DRAM/n2300 ), .B2(\unit_memory/DRAM/n2301 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2284 ) );
  AOI21_X1 U5927 ( .B1(\unit_memory/DRAM/n2296 ), .B2(\unit_memory/DRAM/n2297 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2285 ) );
  NOR4_X1 U5928 ( .A1(\unit_memory/DRAM/n2305 ), .A2(\unit_memory/DRAM/n2306 ), 
        .A3(\unit_memory/DRAM/n2307 ), .A4(\unit_memory/DRAM/n2308 ), .ZN(
        \unit_memory/DRAM/n2304 ) );
  AOI21_X1 U5929 ( .B1(\unit_memory/DRAM/n2321 ), .B2(\unit_memory/DRAM/n2322 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2305 ) );
  AOI21_X1 U5930 ( .B1(\unit_memory/DRAM/n2317 ), .B2(\unit_memory/DRAM/n2318 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2306 ) );
  NOR4_X1 U5931 ( .A1(\unit_memory/DRAM/n2326 ), .A2(\unit_memory/DRAM/n2327 ), 
        .A3(\unit_memory/DRAM/n2328 ), .A4(\unit_memory/DRAM/n2329 ), .ZN(
        \unit_memory/DRAM/n2325 ) );
  AOI21_X1 U5932 ( .B1(\unit_memory/DRAM/n2342 ), .B2(\unit_memory/DRAM/n2343 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2326 ) );
  AOI21_X1 U5933 ( .B1(\unit_memory/DRAM/n2338 ), .B2(\unit_memory/DRAM/n2339 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2327 ) );
  NOR4_X1 U5934 ( .A1(\unit_memory/DRAM/n2347 ), .A2(\unit_memory/DRAM/n2348 ), 
        .A3(\unit_memory/DRAM/n2349 ), .A4(\unit_memory/DRAM/n2350 ), .ZN(
        \unit_memory/DRAM/n2346 ) );
  AOI21_X1 U5935 ( .B1(\unit_memory/DRAM/n2363 ), .B2(\unit_memory/DRAM/n2364 ), .A(\unit_memory/DRAM/n551 ), .ZN(\unit_memory/DRAM/n2347 ) );
  AOI21_X1 U5936 ( .B1(\unit_memory/DRAM/n2359 ), .B2(\unit_memory/DRAM/n2360 ), .A(\unit_memory/DRAM/n550 ), .ZN(\unit_memory/DRAM/n2348 ) );
  AND2_X1 U5937 ( .A1(cw_dec[3]), .A2(n136), .ZN(
        \unit_decode/RegisterFile/N445 ) );
  AND2_X1 U5938 ( .A1(cw_dec[4]), .A2(n134), .ZN(
        \unit_decode/RegisterFile/N444 ) );
  BUF_X1 U5939 ( .A(RST), .Z(n1343) );
  BUF_X1 U5940 ( .A(RST), .Z(n1342) );
  BUF_X1 U5941 ( .A(RST), .Z(n1344) );
  NAND4_X1 U5942 ( .A1(\unit_memory/DRAM/n2200 ), .A2(\unit_memory/DRAM/n2201 ), .A3(\unit_memory/DRAM/n2202 ), .A4(\unit_memory/DRAM/n2203 ), .ZN(
        \unit_memory/DRAM/N573 ) );
  OAI21_X1 U5943 ( .B1(\unit_memory/DRAM/n2208 ), .B2(\unit_memory/DRAM/n2209 ), .A(\unit_memory/DRAM/n1148 ), .ZN(\unit_memory/DRAM/n2202 ) );
  OAI21_X1 U5944 ( .B1(\unit_memory/DRAM/n2216 ), .B2(\unit_memory/DRAM/n2217 ), .A(\unit_memory/DRAM/n548 ), .ZN(\unit_memory/DRAM/n2200 ) );
  NOR2_X1 U5950 ( .A1(IR_OUT[31]), .A2(IR_OUT[29]), .ZN(\unit_decode/n3517 )
         );
  BUF_X1 U5951 ( .A(\unit_fetch/n329 ), .Z(n114) );
  XNOR2_X1 U5952 ( .A(n35), .B(n114), .ZN(\unit_fetch/n674 ) );
  OAI22_X1 U5953 ( .A1(n1285), .A2(\unit_decode/n2194 ), .B1(n1374), .B2(n1296), .ZN(\unit_decode/RD1reg/ffi_0/n5 ) );
  OAI22_X1 U5954 ( .A1(IR_OUT[11]), .A2(n40), .B1(IR_OUT[16]), .B2(
        \unit_decode/n3515 ), .ZN(\unit_decode/n2194 ) );
  INV_X1 U5955 ( .A(n77), .ZN(n1401) );
  INV_X1 U5956 ( .A(n141), .ZN(n139) );
  INV_X1 U5957 ( .A(n141), .ZN(n138) );
  INV_X1 U5958 ( .A(n46), .ZN(net130914) );
  BUF_X1 U5959 ( .A(\unit_decode/n2193 ), .Z(n116) );
  OAI22_X1 U5960 ( .A1(IR_OUT[12]), .A2(n40), .B1(IR_OUT[17]), .B2(
        \unit_decode/n3515 ), .ZN(\unit_decode/n2193 ) );
  BUF_X1 U5961 ( .A(n1423), .Z(n117) );
  INV_X1 U5962 ( .A(n1463), .ZN(n119) );
  AND2_X1 U5963 ( .A1(n1383), .A2(n1471), .ZN(n120) );
  CLKBUF_X1 U5964 ( .A(n119), .Z(n122) );
  CLKBUF_X1 U5965 ( .A(n118), .Z(n123) );
  NAND3_X1 U5966 ( .A1(n78), .A2(n1426), .A3(n1427), .ZN(n1428) );
  CLKBUF_X1 U5967 ( .A(n1471), .Z(n125) );
  OR2_X1 U5968 ( .A1(n1430), .A2(n1429), .ZN(n126) );
  NAND2_X1 U5969 ( .A1(n1428), .A2(n126), .ZN(n1432) );
  INV_X2 U5970 ( .A(n89), .ZN(n141) );
  INV_X1 U5971 ( .A(n1322), .ZN(n1352) );
  INV_X1 U5972 ( .A(cw_dec[2]), .ZN(n128) );
  INV_X1 U5973 ( .A(cw_dec[2]), .ZN(n129) );
  INV_X1 U5974 ( .A(n128), .ZN(n130) );
  INV_X1 U5975 ( .A(n128), .ZN(n131) );
  INV_X1 U5976 ( .A(n128), .ZN(n132) );
  INV_X1 U5977 ( .A(n128), .ZN(n133) );
  INV_X1 U5978 ( .A(n129), .ZN(n134) );
  INV_X1 U5979 ( .A(n129), .ZN(n135) );
  INV_X1 U5980 ( .A(n129), .ZN(n136) );
  INV_X1 U5981 ( .A(n2), .ZN(n137) );
  CLKBUF_X1 U5982 ( .A(net130302), .Z(net130312) );
  INV_X1 U5983 ( .A(n141), .ZN(n140) );
  CLKBUF_X1 U5984 ( .A(n146), .Z(n157) );
  CLKBUF_X1 U5985 ( .A(n159), .Z(n170) );
  CLKBUF_X1 U5986 ( .A(n172), .Z(n183) );
  CLKBUF_X1 U5987 ( .A(n185), .Z(n196) );
  CLKBUF_X1 U5988 ( .A(n198), .Z(n209) );
  CLKBUF_X1 U5989 ( .A(n211), .Z(n222) );
  CLKBUF_X1 U5990 ( .A(n224), .Z(n235) );
  CLKBUF_X1 U5991 ( .A(n237), .Z(n248) );
  INV_X1 U5992 ( .A(\unit_decode/n3512 ), .ZN(n1293) );
  CLKBUF_X1 U5993 ( .A(n1295), .Z(n1305) );
  OAI22_X1 U5994 ( .A1(IR_OUT[15]), .A2(n40), .B1(IR_OUT[20]), .B2(
        \unit_decode/n3515 ), .ZN(\unit_decode/n2190 ) );
  OAI22_X1 U5995 ( .A1(IR_OUT[14]), .A2(n40), .B1(IR_OUT[19]), .B2(n41), .ZN(
        \unit_decode/n2191 ) );
  OAI22_X1 U5996 ( .A1(IR_OUT[13]), .A2(n40), .B1(IR_OUT[18]), .B2(n41), .ZN(
        \unit_decode/n2192 ) );
  NAND2_X1 U5997 ( .A1(\unit_fetch/pc_regout[3] ), .A2(n1539), .ZN(n1492) );
  INV_X1 U5998 ( .A(n1492), .ZN(n1353) );
  NAND4_X1 U5999 ( .A1(n92), .A2(n121), .A3(n124), .A4(n112), .ZN(n1354) );
  NOR4_X1 U6000 ( .A1(n1354), .A2(\unit_fetch/pc_regout[29] ), .A3(
        \unit_fetch/pc_regout[30] ), .A4(\unit_fetch/pc_regout[15] ), .ZN(
        n1360) );
  NAND3_X1 U6001 ( .A1(n1581), .A2(n87), .A3(n76), .ZN(n1355) );
  NOR4_X1 U6002 ( .A1(n1355), .A2(\unit_fetch/pc_regout[26] ), .A3(
        \unit_fetch/pc_regout[27] ), .A4(\unit_fetch/pc_regout[28] ), .ZN(
        n1359) );
  INV_X1 U6003 ( .A(\unit_fetch/pc_regout[11] ), .ZN(n1549) );
  NAND3_X1 U6004 ( .A1(n38), .A2(n1545), .A3(n1543), .ZN(n1356) );
  NOR4_X1 U6005 ( .A1(n1356), .A2(\unit_fetch/pc_regout[12] ), .A3(
        \unit_fetch/pc_regout[14] ), .A4(\unit_fetch/pc_regout[16] ), .ZN(
        n1357) );
  OAI21_X1 U6006 ( .B1(n104), .B2(n105), .A(n72), .ZN(n1478) );
  INV_X1 U6007 ( .A(n1478), .ZN(n1452) );
  INV_X1 U6008 ( .A(n1446), .ZN(n1388) );
  NAND2_X1 U6009 ( .A1(n1452), .A2(n103), .ZN(n1460) );
  INV_X1 U6010 ( .A(n1460), .ZN(n1368) );
  NAND2_X1 U6011 ( .A1(\unit_fetch/pc_regout[2] ), .A2(n114), .ZN(n1421) );
  INV_X1 U6012 ( .A(n1421), .ZN(n1369) );
  NAND2_X1 U6013 ( .A1(n1369), .A2(net130925), .ZN(n1361) );
  NAND2_X1 U6014 ( .A1(n105), .A2(n42), .ZN(n1377) );
  NAND2_X1 U6015 ( .A1(n110), .A2(n104), .ZN(n1380) );
  INV_X1 U6016 ( .A(n1380), .ZN(n1362) );
  INV_X1 U6017 ( .A(n1361), .ZN(n1451) );
  NAND2_X1 U6018 ( .A1(n1362), .A2(n1451), .ZN(n1610) );
  OAI21_X1 U6019 ( .B1(n1361), .B2(n1377), .A(n1610), .ZN(n1621) );
  NAND2_X1 U6020 ( .A1(\unit_fetch/pc_regout[4] ), .A2(n1655), .ZN(n1493) );
  INV_X1 U6021 ( .A(n1493), .ZN(n1392) );
  NAND3_X1 U6022 ( .A1(n114), .A2(n35), .A3(n81), .ZN(n1455) );
  NAND2_X1 U6023 ( .A1(n107), .A2(n81), .ZN(n1400) );
  INV_X1 U6024 ( .A(n1400), .ZN(n1376) );
  NAND2_X1 U6025 ( .A1(n1376), .A2(n77), .ZN(n1384) );
  NAND2_X1 U6026 ( .A1(n1388), .A2(\unit_fetch/pc_regout[2] ), .ZN(n1402) );
  INV_X1 U6027 ( .A(n1402), .ZN(n1378) );
  NAND2_X1 U6028 ( .A1(n1362), .A2(n1378), .ZN(n1476) );
  NAND2_X1 U6029 ( .A1(n1384), .A2(n1476), .ZN(n1464) );
  INV_X1 U6030 ( .A(n1464), .ZN(n1472) );
  NAND3_X1 U6031 ( .A1(net130925), .A2(n110), .A3(n111), .ZN(n1399) );
  INV_X1 U6032 ( .A(n1399), .ZN(n1465) );
  NAND2_X1 U6033 ( .A1(n104), .A2(n1465), .ZN(n1454) );
  OAI211_X1 U6034 ( .C1(n1401), .C2(n1455), .A(n1472), .B(n1454), .ZN(n1363)
         );
  INV_X1 U6035 ( .A(n1363), .ZN(n1436) );
  NAND2_X1 U6036 ( .A1(n106), .A2(n81), .ZN(n1367) );
  INV_X1 U6037 ( .A(n1367), .ZN(n1449) );
  NAND2_X1 U6038 ( .A1(n127), .A2(n1449), .ZN(n1471) );
  NAND2_X1 U6039 ( .A1(n1436), .A2(n125), .ZN(n1620) );
  MUX2_X1 U6040 ( .A(\unit_fetch/pc_regout[3] ), .B(n1539), .S(
        \unit_fetch/pc_regout[5] ), .Z(n1364) );
  NAND3_X1 U6041 ( .A1(n42), .A2(n1492), .A3(n1364), .ZN(n1456) );
  INV_X1 U6042 ( .A(\unit_fetch/n682 ), .ZN(n1365) );
  NAND3_X1 U6043 ( .A1(n1451), .A2(n72), .A3(n1365), .ZN(n1366) );
  OAI21_X1 U6044 ( .B1(n1367), .B2(n1456), .A(n1366), .ZN(n1600) );
  NOR4_X1 U6045 ( .A1(n1368), .A2(n1621), .A3(n1620), .A4(n1600), .ZN(n1435)
         );
  INV_X1 U6046 ( .A(n1455), .ZN(n1382) );
  NAND2_X1 U6047 ( .A1(n1382), .A2(n1452), .ZN(n1608) );
  INV_X1 U6048 ( .A(n1608), .ZN(n1371) );
  NAND2_X1 U6049 ( .A1(n1369), .A2(n35), .ZN(n1479) );
  INV_X1 U6050 ( .A(n1479), .ZN(n1370) );
  NAND2_X1 U6051 ( .A1(n1370), .A2(n72), .ZN(n1457) );
  INV_X1 U6052 ( .A(n1457), .ZN(n1437) );
  NAND2_X1 U6053 ( .A1(n1437), .A2(n104), .ZN(n1473) );
  INV_X1 U6054 ( .A(n1473), .ZN(n1466) );
  NAND2_X1 U6055 ( .A1(n1452), .A2(n1376), .ZN(n1623) );
  INV_X1 U6056 ( .A(n1623), .ZN(n1607) );
  NOR3_X1 U6057 ( .A1(n1371), .A2(n1466), .A3(n1607), .ZN(n1434) );
  NOR3_X1 U6058 ( .A1(rd1_out[2]), .A2(rd1_out[1]), .A3(rd1_out[0]), .ZN(n1373) );
  NAND3_X1 U6059 ( .A1(n1397), .A2(n1386), .A3(n1373), .ZN(n1692) );
  OAI21_X1 U6060 ( .B1(n98), .B2(n1374), .A(\unit_decode/n2194 ), .ZN(n1423)
         );
  OAI21_X1 U6061 ( .B1(n98), .B2(n1375), .A(\unit_decode/n2192 ), .ZN(n1414)
         );
  NOR4_X1 U6062 ( .A1(n103), .A2(n1376), .A3(n1449), .A4(n1382), .ZN(n1381) );
  INV_X1 U6063 ( .A(n1377), .ZN(n1379) );
  NAND2_X1 U6064 ( .A1(n1379), .A2(n1378), .ZN(n1445) );
  OAI211_X1 U6065 ( .C1(n1381), .C2(n1380), .A(n1445), .B(n1610), .ZN(n1613)
         );
  INV_X1 U6066 ( .A(n1613), .ZN(n1385) );
  OAI21_X1 U6067 ( .B1(n1382), .B2(n103), .A(n127), .ZN(n1383) );
  NAND2_X1 U6068 ( .A1(n1383), .A2(n1471), .ZN(n1463) );
  NAND2_X1 U6069 ( .A1(n1451), .A2(n77), .ZN(n1470) );
  NAND4_X1 U6070 ( .A1(n119), .A2(n1454), .A3(n1470), .A4(n1384), .ZN(n1658)
         );
  INV_X1 U6071 ( .A(n1658), .ZN(n1477) );
  NAND3_X1 U6072 ( .A1(n1385), .A2(n1477), .A3(n1473), .ZN(n1484) );
  OAI21_X1 U6073 ( .B1(n98), .B2(n1386), .A(\unit_decode/n2191 ), .ZN(n1417)
         );
  NAND4_X1 U6074 ( .A1(n117), .A2(n1414), .A3(n1484), .A4(n74), .ZN(n1430) );
  OAI21_X1 U6075 ( .B1(n106), .B2(n1388), .A(n1421), .ZN(n1387) );
  NAND2_X1 U6076 ( .A1(n1392), .A2(n1387), .ZN(n1628) );
  INV_X1 U6077 ( .A(n1628), .ZN(n1406) );
  OAI21_X1 U6078 ( .B1(\unit_fetch/n674 ), .B2(\unit_fetch/pc_regout[2] ), .A(
        n88), .ZN(n1390) );
  NAND3_X1 U6079 ( .A1(\unit_fetch/pc_regout[4] ), .A2(
        \unit_fetch/pc_regout[3] ), .A3(n1388), .ZN(n1389) );
  NAND2_X1 U6080 ( .A1(n103), .A2(\unit_fetch/pc_regout[5] ), .ZN(n1395) );
  NAND3_X1 U6081 ( .A1(n1390), .A2(n1389), .A3(n1395), .ZN(n1403) );
  INV_X1 U6082 ( .A(n1403), .ZN(n1598) );
  NAND3_X1 U6083 ( .A1(n1392), .A2(n36), .A3(n81), .ZN(n1419) );
  OAI21_X1 U6084 ( .B1(\unit_fetch/pc_regout[2] ), .B2(net130925), .A(n1421), 
        .ZN(n1391) );
  NAND2_X1 U6085 ( .A1(n88), .A2(n1391), .ZN(n1411) );
  NAND3_X1 U6086 ( .A1(n1419), .A2(n1492), .A3(n1411), .ZN(n1679) );
  NAND2_X1 U6087 ( .A1(\unit_fetch/pc_regout[2] ), .A2(n1697), .ZN(n1393) );
  MUX2_X1 U6088 ( .A(n1393), .B(n1446), .S(\unit_fetch/pc_regout[4] ), .Z(
        n1394) );
  OAI211_X1 U6089 ( .C1(n1493), .C2(n111), .A(n1395), .B(n1394), .ZN(n1669) );
  NAND3_X1 U6090 ( .A1(n1406), .A2(n101), .A3(n1669), .ZN(n1408) );
  INV_X1 U6091 ( .A(n1408), .ZN(n1688) );
  OAI21_X1 U6092 ( .B1(n118), .B2(n1396), .A(n116), .ZN(n1424) );
  OAI21_X1 U6093 ( .B1(n1694), .B2(n1397), .A(\unit_decode/n2190 ), .ZN(n1398)
         );
  INV_X1 U6094 ( .A(n1398), .ZN(n1413) );
  OAI22_X1 U6095 ( .A1(n1456), .A2(n1400), .B1(\unit_fetch/n682 ), .B2(n1399), 
        .ZN(n1480) );
  OAI21_X1 U6096 ( .B1(n1401), .B2(n1421), .A(n120), .ZN(n1416) );
  INV_X1 U6097 ( .A(n1416), .ZN(n1486) );
  INV_X1 U6098 ( .A(n1599), .ZN(n1425) );
  NAND4_X1 U6099 ( .A1(n1688), .A2(n1424), .A3(n1413), .A4(n1425), .ZN(n1429)
         );
  OAI21_X1 U6100 ( .B1(n1492), .B2(n1402), .A(n1628), .ZN(n1404) );
  INV_X1 U6101 ( .A(n1404), .ZN(n1681) );
  NAND2_X1 U6102 ( .A1(n1681), .A2(n1403), .ZN(n1405) );
  INV_X1 U6103 ( .A(n1405), .ZN(n1676) );
  NAND2_X1 U6104 ( .A1(n1676), .A2(n1679), .ZN(n1674) );
  NAND2_X1 U6105 ( .A1(n59), .A2(n58), .ZN(n1673) );
  OAI211_X1 U6106 ( .C1(n1405), .C2(n1669), .A(n1674), .B(n1673), .ZN(n1670)
         );
  INV_X1 U6107 ( .A(n1670), .ZN(n1409) );
  NAND2_X1 U6108 ( .A1(n57), .A2(n101), .ZN(n1667) );
  INV_X1 U6109 ( .A(n1679), .ZN(n1490) );
  NAND2_X1 U6110 ( .A1(n1490), .A2(n1406), .ZN(n1686) );
  NAND2_X1 U6111 ( .A1(n1667), .A2(n1686), .ZN(n1687) );
  INV_X1 U6112 ( .A(n1687), .ZN(n1407) );
  NAND3_X1 U6113 ( .A1(n1409), .A2(n1408), .A3(n1407), .ZN(n1410) );
  NAND2_X1 U6114 ( .A1(n1410), .A2(n1667), .ZN(n1666) );
  OAI21_X1 U6115 ( .B1(n80), .B2(\unit_fetch/pc_regout[3] ), .A(
        \unit_fetch/pc_regout[4] ), .ZN(n1418) );
  NAND3_X1 U6116 ( .A1(n1697), .A2(n36), .A3(n1418), .ZN(n1412) );
  NAND2_X1 U6117 ( .A1(n1412), .A2(n1411), .ZN(n1488) );
  INV_X1 U6118 ( .A(n1414), .ZN(n1415) );
  NAND3_X1 U6119 ( .A1(n1697), .A2(n35), .A3(n1418), .ZN(n1420) );
  OAI211_X1 U6120 ( .C1(n1493), .C2(n1421), .A(n1420), .B(n1419), .ZN(n1422)
         );
  INV_X1 U6121 ( .A(n1422), .ZN(n1487) );
  AOI21_X1 U6122 ( .B1(n1435), .B2(n1434), .A(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n96 ) );
  NAND2_X1 U6123 ( .A1(n77), .A2(n103), .ZN(n1469) );
  NAND2_X1 U6124 ( .A1(n1436), .A2(n1469), .ZN(n1601) );
  INV_X1 U6125 ( .A(n1601), .ZN(n1611) );
  NOR2_X1 U6126 ( .A1(n1611), .A2(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n91 ) );
  NAND2_X1 U6127 ( .A1(n105), .A2(n1437), .ZN(n1612) );
  NAND4_X1 U6128 ( .A1(n1472), .A2(n122), .A3(n1612), .A4(n1473), .ZN(n1458)
         );
  INV_X1 U6129 ( .A(n1458), .ZN(n1438) );
  NAND2_X1 U6130 ( .A1(n1438), .A2(n1608), .ZN(n1450) );
  INV_X1 U6131 ( .A(n1450), .ZN(n1448) );
  NOR4_X1 U6132 ( .A1(n1593), .A2(n1589), .A3(n1583), .A4(n1587), .ZN(n1444)
         );
  NOR4_X1 U6133 ( .A1(n1581), .A2(n87), .A3(n76), .A4(n1573), .ZN(n1443) );
  NOR4_X1 U6134 ( .A1(n1559), .A2(n1555), .A3(n1553), .A4(n1651), .ZN(n1441)
         );
  NAND3_X1 U6135 ( .A1(\unit_fetch/pc_regout[2] ), .A2(
        \unit_fetch/pc_regout[3] ), .A3(\unit_fetch/pc_regout[4] ), .ZN(n1647)
         );
  INV_X1 U6136 ( .A(n1498), .ZN(n1646) );
  NOR4_X1 U6137 ( .A1(n92), .A2(n1543), .A3(n121), .A4(n124), .ZN(n1439) );
  NAND2_X1 U6138 ( .A1(n1646), .A2(n1439), .ZN(n1504) );
  INV_X1 U6139 ( .A(n1504), .ZN(n1540) );
  NOR4_X1 U6140 ( .A1(n112), .A2(n1551), .A3(n1549), .A4(n1545), .ZN(n1440) );
  NAND2_X1 U6141 ( .A1(n1540), .A2(n1440), .ZN(n1510) );
  INV_X1 U6142 ( .A(n1510), .ZN(n1636) );
  NAND2_X1 U6143 ( .A1(n1441), .A2(n1636), .ZN(n1516) );
  NOR3_X1 U6144 ( .A1(n1561), .A2(n1516), .A3(n1565), .ZN(n1442) );
  NAND3_X1 U6145 ( .A1(\unit_fetch/pc_regout[20] ), .A2(
        \unit_fetch/pc_regout[21] ), .A3(n1442), .ZN(n1522) );
  INV_X1 U6146 ( .A(n1522), .ZN(n1568) );
  NAND2_X1 U6147 ( .A1(n1443), .A2(n1568), .ZN(n1528) );
  INV_X1 U6148 ( .A(n1528), .ZN(n1578) );
  NAND2_X1 U6149 ( .A1(n1444), .A2(n1578), .ZN(n1535) );
  INV_X1 U6150 ( .A(n1535), .ZN(n1590) );
  NAND2_X1 U6151 ( .A1(\unit_fetch/pc_regout[30] ), .A2(n1590), .ZN(n1534) );
  OAI211_X1 U6152 ( .C1(n1446), .C2(n1534), .A(n1445), .B(n1460), .ZN(n1617)
         );
  INV_X1 U6153 ( .A(n1617), .ZN(n1447) );
  AOI21_X1 U6154 ( .B1(n1448), .B2(n1447), .A(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n90 ) );
  NAND2_X1 U6155 ( .A1(n1452), .A2(n1449), .ZN(n1624) );
  INV_X1 U6156 ( .A(n1624), .ZN(n1618) );
  NOR2_X1 U6157 ( .A1(n1618), .A2(n1450), .ZN(n1453) );
  NAND2_X1 U6158 ( .A1(n1452), .A2(n1451), .ZN(n1659) );
  AOI21_X1 U6159 ( .B1(n1453), .B2(n1659), .A(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n89 ) );
  INV_X1 U6160 ( .A(n1454), .ZN(n1459) );
  OAI22_X1 U6161 ( .A1(\unit_fetch/n682 ), .A2(n1457), .B1(n1456), .B2(n1455), 
        .ZN(n1603) );
  NOR3_X1 U6162 ( .A1(n1459), .A2(n1603), .A3(n1458), .ZN(n1462) );
  NAND2_X1 U6163 ( .A1(n1659), .A2(n1460), .ZN(n1475) );
  NOR2_X1 U6164 ( .A1(n1607), .A2(n1475), .ZN(n1461) );
  AOI21_X1 U6165 ( .B1(n1462), .B2(n1461), .A(n140), .ZN(
        \unit_fetch/unit_instructionRegister/n88 ) );
  NOR3_X1 U6166 ( .A1(n1464), .A2(n1463), .A3(n1613), .ZN(n1468) );
  NAND2_X1 U6167 ( .A1(n105), .A2(n1465), .ZN(n1622) );
  INV_X1 U6168 ( .A(n1622), .ZN(n1614) );
  NOR2_X1 U6169 ( .A1(n1466), .A2(n1614), .ZN(n1467) );
  AOI21_X1 U6170 ( .B1(n1468), .B2(n1467), .A(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n87 ) );
  NAND4_X1 U6171 ( .A1(n1472), .A2(n125), .A3(n1470), .A4(n1469), .ZN(n1604)
         );
  INV_X1 U6172 ( .A(n1604), .ZN(n1474) );
  AOI21_X1 U6173 ( .B1(n1474), .B2(n1473), .A(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n85 ) );
  NOR2_X1 U6174 ( .A1(n1474), .A2(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n83 ) );
  INV_X1 U6175 ( .A(n1475), .ZN(n1483) );
  INV_X1 U6176 ( .A(n1476), .ZN(n1481) );
  OAI211_X1 U6177 ( .C1(n1479), .C2(n1478), .A(n1477), .B(n1622), .ZN(n1606)
         );
  NOR3_X1 U6178 ( .A1(n1481), .A2(n1480), .A3(n1606), .ZN(n1482) );
  AOI21_X1 U6179 ( .B1(n1483), .B2(n1482), .A(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n80 ) );
  INV_X1 U6180 ( .A(n1484), .ZN(n1485) );
  NOR2_X1 U6181 ( .A1(n1485), .A2(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n79 ) );
  NOR2_X1 U6182 ( .A1(n1486), .A2(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n67 ) );
  NOR2_X1 U6183 ( .A1(n1487), .A2(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n75 ) );
  INV_X1 U6184 ( .A(n1488), .ZN(n1489) );
  NOR2_X1 U6185 ( .A1(n1489), .A2(n140), .ZN(
        \unit_fetch/unit_instructionRegister/n74 ) );
  NOR2_X1 U6186 ( .A1(n1490), .A2(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n73 ) );
  NOR2_X1 U6187 ( .A1(n57), .A2(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n72 ) );
  NAND2_X1 U6188 ( .A1(n115), .A2(n1352), .ZN(net126982) );
  MUX2_X1 U6189 ( .A(n1539), .B(n1492), .S(n80), .Z(n1494) );
  NAND2_X1 U6190 ( .A1(n1494), .A2(n1493), .ZN(n1495) );
  MUX2_X1 U6191 ( .A(n1495), .B(alu_out[4]), .S(jump), .Z(n1496) );
  NAND2_X1 U6192 ( .A1(n1496), .A2(n141), .ZN(n1538) );
  OAI21_X1 U6193 ( .B1(\unit_decode/n2144 ), .B2(net130306), .A(n1538), .ZN(
        \unit_fetch/unit_npcregister/ffi_4/n5 ) );
  NAND2_X1 U6194 ( .A1(n1646), .A2(\unit_fetch/pc_regout[6] ), .ZN(n1644) );
  INV_X1 U6195 ( .A(n1644), .ZN(n1500) );
  INV_X1 U6196 ( .A(jump), .ZN(n1497) );
  AOI211_X1 U6197 ( .C1(n1498), .C2(n124), .A(n1500), .B(n45), .ZN(n1499) );
  AOI21_X1 U6198 ( .B1(alu_out[6]), .B2(net130324), .A(n1499), .ZN(n1661) );
  OAI21_X1 U6199 ( .B1(\unit_decode/n2142 ), .B2(net130312), .A(n1661), .ZN(
        \unit_fetch/unit_npcregister/ffi_6/n5 ) );
  NAND2_X1 U6200 ( .A1(n1500), .A2(\unit_fetch/pc_regout[7] ), .ZN(n1502) );
  INV_X1 U6201 ( .A(n1502), .ZN(n1643) );
  NAND2_X1 U6202 ( .A1(n1643), .A2(\unit_fetch/pc_regout[8] ), .ZN(n1541) );
  INV_X1 U6203 ( .A(n1541), .ZN(n1501) );
  AOI211_X1 U6204 ( .C1(n1502), .C2(n92), .A(n1501), .B(n45), .ZN(n1503) );
  AOI21_X1 U6205 ( .B1(alu_out[8]), .B2(net130326), .A(n1503), .ZN(n1656) );
  OAI21_X1 U6206 ( .B1(\unit_decode/n2140 ), .B2(net130312), .A(n1656), .ZN(
        \unit_fetch/unit_npcregister/ffi_8/n5 ) );
  NAND2_X1 U6207 ( .A1(n1540), .A2(\unit_fetch/pc_regout[10] ), .ZN(n1547) );
  INV_X1 U6208 ( .A(n1547), .ZN(n1506) );
  AOI211_X1 U6209 ( .C1(n1504), .C2(n1545), .A(n1506), .B(n45), .ZN(n1505) );
  AOI21_X1 U6210 ( .B1(alu_out[10]), .B2(n50), .A(n1505), .ZN(n1544) );
  OAI21_X1 U6211 ( .B1(\unit_decode/n2138 ), .B2(net130312), .A(n1544), .ZN(
        \unit_fetch/unit_npcregister/ffi_10/n5 ) );
  NAND2_X1 U6212 ( .A1(n1506), .A2(\unit_fetch/pc_regout[11] ), .ZN(n1508) );
  INV_X1 U6213 ( .A(n1508), .ZN(n1546) );
  NAND2_X1 U6214 ( .A1(n1546), .A2(\unit_fetch/pc_regout[12] ), .ZN(n1637) );
  INV_X1 U6215 ( .A(n1637), .ZN(n1507) );
  AOI211_X1 U6216 ( .C1(n1508), .C2(n1551), .A(n1507), .B(n47), .ZN(n1509) );
  AOI21_X1 U6217 ( .B1(alu_out[12]), .B2(n50), .A(n1509), .ZN(n1550) );
  OAI21_X1 U6218 ( .B1(\unit_decode/n2136 ), .B2(net130310), .A(n1550), .ZN(
        \unit_fetch/unit_npcregister/ffi_12/n5 ) );
  NAND2_X1 U6219 ( .A1(\unit_fetch/pc_regout[14] ), .A2(n1636), .ZN(n1634) );
  INV_X1 U6220 ( .A(n1634), .ZN(n1512) );
  AOI211_X1 U6221 ( .C1(n1510), .C2(n1553), .A(n1512), .B(n46), .ZN(n1511) );
  AOI21_X1 U6222 ( .B1(alu_out[14]), .B2(net130324), .A(n1511), .ZN(n1552) );
  OAI21_X1 U6223 ( .B1(\unit_decode/n2134 ), .B2(net130310), .A(n1552), .ZN(
        \unit_fetch/unit_npcregister/ffi_14/n5 ) );
  NAND2_X1 U6224 ( .A1(\unit_fetch/pc_regout[15] ), .A2(n1512), .ZN(n1514) );
  INV_X1 U6225 ( .A(n1514), .ZN(n1633) );
  NAND2_X1 U6226 ( .A1(n1633), .A2(\unit_fetch/pc_regout[16] ), .ZN(n1557) );
  INV_X1 U6227 ( .A(n1557), .ZN(n1513) );
  AOI211_X1 U6228 ( .C1(n1514), .C2(n1555), .A(n1513), .B(n45), .ZN(n1515) );
  AOI21_X1 U6229 ( .B1(alu_out[16]), .B2(net130324), .A(n1515), .ZN(n1554) );
  OAI21_X1 U6230 ( .B1(\unit_decode/n2132 ), .B2(net130310), .A(n1554), .ZN(
        \unit_fetch/unit_npcregister/ffi_16/n5 ) );
  INV_X1 U6231 ( .A(n1516), .ZN(n1556) );
  NAND2_X1 U6232 ( .A1(\unit_fetch/pc_regout[18] ), .A2(n1556), .ZN(n1563) );
  INV_X1 U6233 ( .A(n1563), .ZN(n1518) );
  AOI211_X1 U6234 ( .C1(n1516), .C2(n1561), .A(n1518), .B(n46), .ZN(n1517) );
  AOI21_X1 U6235 ( .B1(alu_out[18]), .B2(net130326), .A(n1517), .ZN(n1560) );
  OAI21_X1 U6236 ( .B1(\unit_decode/n2130 ), .B2(net130310), .A(n1560), .ZN(
        \unit_fetch/unit_npcregister/ffi_18/n5 ) );
  NAND2_X1 U6237 ( .A1(n1518), .A2(\unit_fetch/pc_regout[19] ), .ZN(n1520) );
  INV_X1 U6238 ( .A(n1520), .ZN(n1562) );
  NAND2_X1 U6239 ( .A1(n1562), .A2(\unit_fetch/pc_regout[20] ), .ZN(n1569) );
  INV_X1 U6240 ( .A(n1569), .ZN(n1519) );
  AOI211_X1 U6241 ( .C1(n1520), .C2(n1567), .A(n1519), .B(n46), .ZN(n1521) );
  AOI21_X1 U6242 ( .B1(alu_out[20]), .B2(n50), .A(n1521), .ZN(n1566) );
  OAI21_X1 U6243 ( .B1(\unit_decode/n2128 ), .B2(net130310), .A(n1566), .ZN(
        \unit_fetch/unit_npcregister/ffi_20/n5 ) );
  NAND2_X1 U6244 ( .A1(n1568), .A2(\unit_fetch/pc_regout[22] ), .ZN(n1575) );
  INV_X1 U6245 ( .A(n1575), .ZN(n1524) );
  AOI211_X1 U6246 ( .C1(n1522), .C2(n1573), .A(n1524), .B(n46), .ZN(n1523) );
  AOI21_X1 U6247 ( .B1(alu_out[22]), .B2(net130324), .A(n1523), .ZN(n1572) );
  OAI21_X1 U6248 ( .B1(\unit_decode/n2126 ), .B2(net130310), .A(n1572), .ZN(
        \unit_fetch/unit_npcregister/ffi_22/n5 ) );
  NAND2_X1 U6249 ( .A1(n1524), .A2(\unit_fetch/pc_regout[23] ), .ZN(n1526) );
  INV_X1 U6250 ( .A(n1526), .ZN(n1574) );
  NAND2_X1 U6251 ( .A1(n1574), .A2(\unit_fetch/pc_regout[24] ), .ZN(n1579) );
  INV_X1 U6252 ( .A(n1579), .ZN(n1525) );
  AOI211_X1 U6253 ( .C1(n1526), .C2(n87), .A(n1525), .B(n45), .ZN(n1527) );
  AOI21_X1 U6254 ( .B1(alu_out[24]), .B2(net130326), .A(n1527), .ZN(n1577) );
  OAI21_X1 U6255 ( .B1(\unit_decode/n2124 ), .B2(net130310), .A(n1577), .ZN(
        \unit_fetch/unit_npcregister/ffi_24/n5 ) );
  NAND2_X1 U6256 ( .A1(\unit_fetch/pc_regout[26] ), .A2(n1578), .ZN(n1585) );
  INV_X1 U6257 ( .A(n1585), .ZN(n1530) );
  AOI211_X1 U6258 ( .C1(n1528), .C2(n1583), .A(n1530), .B(n46), .ZN(n1529) );
  AOI21_X1 U6259 ( .B1(alu_out[26]), .B2(net130324), .A(n1529), .ZN(n1582) );
  OAI21_X1 U6260 ( .B1(\unit_decode/n2122 ), .B2(net130310), .A(n1582), .ZN(
        \unit_fetch/unit_npcregister/ffi_26/n5 ) );
  NAND2_X1 U6261 ( .A1(\unit_fetch/pc_regout[27] ), .A2(n1530), .ZN(n1532) );
  INV_X1 U6262 ( .A(n1532), .ZN(n1584) );
  NAND2_X1 U6263 ( .A1(n1584), .A2(\unit_fetch/pc_regout[28] ), .ZN(n1591) );
  INV_X1 U6264 ( .A(n1591), .ZN(n1531) );
  AOI211_X1 U6265 ( .C1(n1532), .C2(n1589), .A(n1531), .B(n47), .ZN(n1533) );
  AOI21_X1 U6266 ( .B1(alu_out[28]), .B2(net130326), .A(n1533), .ZN(n1588) );
  OAI21_X1 U6267 ( .B1(\unit_decode/n2120 ), .B2(net130310), .A(n1588), .ZN(
        \unit_fetch/unit_npcregister/ffi_28/n5 ) );
  INV_X1 U6268 ( .A(n1534), .ZN(n1625) );
  AOI211_X1 U6269 ( .C1(n1535), .C2(n1595), .A(n1625), .B(n45), .ZN(n1536) );
  AOI21_X1 U6270 ( .B1(alu_out[30]), .B2(net130326), .A(n1536), .ZN(n1594) );
  OAI21_X1 U6271 ( .B1(\unit_decode/n2118 ), .B2(net130310), .A(n1594), .ZN(
        \unit_fetch/unit_npcregister/ffi_30/n5 ) );
  XOR2_X1 U6272 ( .A(\unit_fetch/pc_regout[31] ), .B(n1625), .Z(n1537) );
  AOI22_X1 U6273 ( .A1(n1537), .A2(net130914), .B1(alu_out[31]), .B2(net130328), .ZN(n1596) );
  OAI21_X1 U6274 ( .B1(\unit_decode/n2117 ), .B2(net130310), .A(n1596), .ZN(
        \unit_fetch/unit_npcregister/ffi_31/n5 ) );
  OAI21_X1 U6275 ( .B1(n1539), .B2(net130310), .A(n1538), .ZN(
        \unit_fetch/unit_programCounter/ffi_4/n5 ) );
  AOI211_X1 U6276 ( .C1(n1541), .C2(n1543), .A(n1540), .B(n47), .ZN(n1542) );
  AOI21_X1 U6277 ( .B1(alu_out[9]), .B2(n50), .A(n1542), .ZN(n1640) );
  OAI21_X1 U6278 ( .B1(net141182), .B2(n1543), .A(n1640), .ZN(
        \unit_fetch/unit_programCounter/ffi_9/n5 ) );
  OAI21_X1 U6279 ( .B1(net141182), .B2(n1545), .A(n1544), .ZN(
        \unit_fetch/unit_programCounter/ffi_10/n5 ) );
  AOI211_X1 U6280 ( .C1(n1547), .C2(n1549), .A(n1546), .B(n46), .ZN(n1548) );
  AOI21_X1 U6281 ( .B1(alu_out[11]), .B2(net130326), .A(n1548), .ZN(n1639) );
  OAI21_X1 U6282 ( .B1(net130304), .B2(n1549), .A(n1639), .ZN(
        \unit_fetch/unit_programCounter/ffi_11/n5 ) );
  OAI21_X1 U6283 ( .B1(net130304), .B2(n1551), .A(n1550), .ZN(
        \unit_fetch/unit_programCounter/ffi_12/n5 ) );
  OAI21_X1 U6284 ( .B1(net141182), .B2(n1553), .A(n1552), .ZN(
        \unit_fetch/unit_programCounter/ffi_14/n5 ) );
  OAI21_X1 U6285 ( .B1(net130304), .B2(n1555), .A(n1554), .ZN(
        \unit_fetch/unit_programCounter/ffi_16/n5 ) );
  AOI211_X1 U6286 ( .C1(n1557), .C2(n1559), .A(n1556), .B(n45), .ZN(n1558) );
  OAI21_X1 U6287 ( .B1(net130304), .B2(n1559), .A(n60), .ZN(
        \unit_fetch/unit_programCounter/ffi_17/n5 ) );
  OAI21_X1 U6288 ( .B1(net141182), .B2(n1561), .A(n1560), .ZN(
        \unit_fetch/unit_programCounter/ffi_18/n5 ) );
  AOI211_X1 U6289 ( .C1(n1563), .C2(n1565), .A(n1562), .B(n45), .ZN(n1564) );
  AOI21_X1 U6290 ( .B1(alu_out[19]), .B2(net130328), .A(n1564), .ZN(n1632) );
  OAI21_X1 U6291 ( .B1(net130304), .B2(n1565), .A(n1632), .ZN(
        \unit_fetch/unit_programCounter/ffi_19/n5 ) );
  OAI21_X1 U6292 ( .B1(net141182), .B2(n1567), .A(n1566), .ZN(
        \unit_fetch/unit_programCounter/ffi_20/n5 ) );
  AOI211_X1 U6293 ( .C1(n1569), .C2(n1571), .A(n1568), .B(n46), .ZN(n1570) );
  AOI21_X1 U6294 ( .B1(alu_out[21]), .B2(net130328), .A(n1570), .ZN(n1631) );
  OAI21_X1 U6295 ( .B1(net141182), .B2(n1571), .A(n1631), .ZN(
        \unit_fetch/unit_programCounter/ffi_21/n5 ) );
  OAI21_X1 U6296 ( .B1(net130304), .B2(n1573), .A(n1572), .ZN(
        \unit_fetch/unit_programCounter/ffi_22/n5 ) );
  AOI211_X1 U6297 ( .C1(n1575), .C2(n76), .A(n1574), .B(n47), .ZN(n1576) );
  AOI21_X1 U6298 ( .B1(alu_out[23]), .B2(n50), .A(n1576), .ZN(n1630) );
  OAI21_X1 U6299 ( .B1(net130304), .B2(n76), .A(n1630), .ZN(
        \unit_fetch/unit_programCounter/ffi_23/n5 ) );
  OAI21_X1 U6300 ( .B1(net130304), .B2(n87), .A(n1577), .ZN(
        \unit_fetch/unit_programCounter/ffi_24/n5 ) );
  AOI211_X1 U6301 ( .C1(n1579), .C2(n1581), .A(n1578), .B(n46), .ZN(n1580) );
  AOI21_X1 U6302 ( .B1(alu_out[25]), .B2(n50), .A(n1580), .ZN(n1629) );
  OAI21_X1 U6303 ( .B1(net130306), .B2(n1583), .A(n1582), .ZN(
        \unit_fetch/unit_programCounter/ffi_26/n5 ) );
  AOI211_X1 U6304 ( .C1(n1585), .C2(n1587), .A(n1584), .B(n47), .ZN(n1586) );
  AOI21_X1 U6305 ( .B1(alu_out[27]), .B2(net130326), .A(n1586), .ZN(n1642) );
  OAI21_X1 U6306 ( .B1(net130304), .B2(n1587), .A(n52), .ZN(
        \unit_fetch/unit_programCounter/ffi_27/n5 ) );
  OAI21_X1 U6307 ( .B1(net130304), .B2(n1589), .A(n1588), .ZN(
        \unit_fetch/unit_programCounter/ffi_28/n5 ) );
  AOI211_X1 U6308 ( .C1(n1591), .C2(n1593), .A(n1590), .B(n45), .ZN(n1592) );
  AOI21_X1 U6309 ( .B1(alu_out[29]), .B2(net130326), .A(n1592), .ZN(n1641) );
  OAI21_X1 U6310 ( .B1(net130306), .B2(n1593), .A(n1641), .ZN(
        \unit_fetch/unit_programCounter/ffi_29/n5 ) );
  OAI21_X1 U6311 ( .B1(net130304), .B2(n1595), .A(n1594), .ZN(
        \unit_fetch/unit_programCounter/ffi_30/n5 ) );
  OAI21_X1 U6312 ( .B1(net130306), .B2(n1597), .A(n1596), .ZN(
        \unit_fetch/unit_programCounter/ffi_31/n5 ) );
  INV_X1 U6313 ( .A(n1669), .ZN(n1680) );
  NAND2_X1 U6314 ( .A1(n1680), .A2(n48), .ZN(
        \unit_fetch/unit_instructionRegister/n68 ) );
  NAND2_X1 U6315 ( .A1(n48), .A2(n1598), .ZN(
        \unit_fetch/unit_instructionRegister/n69 ) );
  OAI21_X1 U6316 ( .B1(n1601), .B2(n1600), .A(n141), .ZN(n1602) );
  INV_X1 U6317 ( .A(n1602), .ZN(\unit_fetch/unit_instructionRegister/n92 ) );
  OAI21_X1 U6318 ( .B1(n1604), .B2(n1603), .A(n141), .ZN(n1605) );
  INV_X1 U6319 ( .A(n1605), .ZN(\unit_fetch/unit_instructionRegister/n84 ) );
  NOR2_X1 U6320 ( .A1(n1607), .A2(n1606), .ZN(n1609) );
  AOI21_X1 U6321 ( .B1(n1609), .B2(n1608), .A(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n81 ) );
  AOI21_X1 U6322 ( .B1(n1611), .B2(n1610), .A(n140), .ZN(
        \unit_fetch/unit_instructionRegister/n93 ) );
  INV_X1 U6323 ( .A(n1612), .ZN(n1615) );
  NOR4_X1 U6324 ( .A1(n1615), .A2(n1614), .A3(n1613), .A4(n1620), .ZN(n1616)
         );
  NOR2_X1 U6325 ( .A1(n1616), .A2(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n95 ) );
  NOR4_X1 U6326 ( .A1(n1618), .A2(n1621), .A3(n1620), .A4(n1617), .ZN(n1619)
         );
  NOR2_X1 U6327 ( .A1(n1619), .A2(n138), .ZN(
        \unit_fetch/unit_instructionRegister/n97 ) );
  NOR2_X1 U6328 ( .A1(n1621), .A2(n1620), .ZN(n1627) );
  NAND3_X1 U6329 ( .A1(n1624), .A2(n1623), .A3(n1622), .ZN(n1657) );
  AOI21_X1 U6330 ( .B1(n1625), .B2(n107), .A(n1657), .ZN(n1626) );
  AOI21_X1 U6331 ( .B1(n1627), .B2(n1626), .A(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n98 ) );
  NOR2_X1 U6332 ( .A1(n58), .A2(n139), .ZN(
        \unit_fetch/unit_instructionRegister/n71 ) );
  OAI21_X1 U6333 ( .B1(\unit_decode/n2123 ), .B2(net130308), .A(n1629), .ZN(
        \unit_fetch/unit_npcregister/ffi_25/n5 ) );
  OAI21_X1 U6334 ( .B1(\unit_decode/n2125 ), .B2(net130308), .A(n1630), .ZN(
        \unit_fetch/unit_npcregister/ffi_23/n5 ) );
  OAI21_X1 U6335 ( .B1(\unit_decode/n2127 ), .B2(net130308), .A(n1631), .ZN(
        \unit_fetch/unit_npcregister/ffi_21/n5 ) );
  OAI21_X1 U6336 ( .B1(\unit_decode/n2129 ), .B2(net130308), .A(n1632), .ZN(
        \unit_fetch/unit_npcregister/ffi_19/n5 ) );
  OAI21_X1 U6337 ( .B1(\unit_decode/n2131 ), .B2(net130308), .A(n60), .ZN(
        \unit_fetch/unit_npcregister/ffi_17/n5 ) );
  AOI211_X1 U6338 ( .C1(n1634), .C2(n1651), .A(n1633), .B(n45), .ZN(n1635) );
  AOI21_X1 U6339 ( .B1(alu_out[15]), .B2(n50), .A(n1635), .ZN(n1650) );
  OAI21_X1 U6340 ( .B1(\unit_decode/n2133 ), .B2(net130308), .A(n1650), .ZN(
        \unit_fetch/unit_npcregister/ffi_15/n5 ) );
  AOI211_X1 U6341 ( .C1(n1637), .C2(n112), .A(n1636), .B(n46), .ZN(n1638) );
  AOI21_X1 U6342 ( .B1(alu_out[13]), .B2(net130326), .A(n1638), .ZN(n1663) );
  OAI21_X1 U6343 ( .B1(\unit_decode/n2135 ), .B2(net130308), .A(n1663), .ZN(
        \unit_fetch/unit_npcregister/ffi_13/n5 ) );
  OAI21_X1 U6344 ( .B1(\unit_decode/n2137 ), .B2(net130308), .A(n1639), .ZN(
        \unit_fetch/unit_npcregister/ffi_11/n5 ) );
  OAI21_X1 U6345 ( .B1(\unit_decode/n2139 ), .B2(net130308), .A(n1640), .ZN(
        \unit_fetch/unit_npcregister/ffi_9/n5 ) );
  OAI21_X1 U6346 ( .B1(\unit_decode/n2119 ), .B2(net130306), .A(n1641), .ZN(
        \unit_fetch/unit_npcregister/ffi_29/n5 ) );
  OAI21_X1 U6347 ( .B1(\unit_decode/n2121 ), .B2(net130308), .A(n1642), .ZN(
        \unit_fetch/unit_npcregister/ffi_27/n5 ) );
  AOI211_X1 U6348 ( .C1(n1644), .C2(n121), .A(n1643), .B(n47), .ZN(n1645) );
  OAI21_X1 U6349 ( .B1(\unit_decode/n2141 ), .B2(net130306), .A(n1662), .ZN(
        \unit_fetch/unit_npcregister/ffi_7/n5 ) );
  AOI211_X1 U6350 ( .C1(n1647), .C2(n1697), .A(n1646), .B(n47), .ZN(n1648) );
  AOI21_X1 U6351 ( .B1(alu_out[5]), .B2(net130324), .A(n1648), .ZN(n1653) );
  OAI21_X1 U6352 ( .B1(\unit_decode/n2143 ), .B2(net130306), .A(n1653), .ZN(
        \unit_fetch/unit_npcregister/ffi_5/n5 ) );
  XOR2_X1 U6353 ( .A(n80), .B(\unit_fetch/pc_regout[3] ), .Z(n1649) );
  AOI22_X1 U6354 ( .A1(net130914), .A2(n1649), .B1(alu_out[3]), .B2(net130328), 
        .ZN(n1654) );
  OAI21_X1 U6355 ( .B1(\unit_decode/n2145 ), .B2(net130306), .A(n1654), .ZN(
        \unit_fetch/unit_npcregister/ffi_3/n5 ) );
  AOI22_X1 U6356 ( .A1(net130914), .A2(n81), .B1(alu_out[2]), .B2(net130328), 
        .ZN(n1664) );
  OAI21_X1 U6357 ( .B1(\unit_decode/n2146 ), .B2(net130306), .A(n1664), .ZN(
        \unit_fetch/unit_npcregister/ffi_2/n5 ) );
  NAND2_X1 U6358 ( .A1(alu_out[1]), .A2(n50), .ZN(n1652) );
  OAI221_X1 U6359 ( .B1(n114), .B2(n46), .C1(\unit_decode/n2147 ), .C2(
        net130306), .A(n1652), .ZN(\unit_fetch/unit_npcregister/ffi_1/n5 ) );
  OAI21_X1 U6360 ( .B1(net141182), .B2(n1651), .A(n1650), .ZN(
        \unit_fetch/unit_programCounter/ffi_15/n5 ) );
  OAI21_X1 U6361 ( .B1(jump), .B2(n1336), .A(net141181), .ZN(net127003) );
  INV_X1 U6362 ( .A(net127003), .ZN(net126984) );
  OAI21_X1 U6363 ( .B1(n114), .B2(net126984), .A(n1652), .ZN(
        \unit_fetch/unit_programCounter/ffi_1/n5 ) );
  OAI21_X1 U6364 ( .B1(n1697), .B2(net130306), .A(n1653), .ZN(
        \unit_fetch/unit_programCounter/ffi_5/n5 ) );
  OAI21_X1 U6365 ( .B1(n1655), .B2(net130308), .A(n1654), .ZN(
        \unit_fetch/unit_programCounter/ffi_3/n5 ) );
  OAI21_X1 U6366 ( .B1(net141182), .B2(n92), .A(n1656), .ZN(
        \unit_fetch/unit_programCounter/ffi_8/n5 ) );
  NOR2_X1 U6367 ( .A1(n102), .A2(n140), .ZN(\unit_fetch/n462 ) );
  NOR2_X1 U6368 ( .A1(n1658), .A2(n1657), .ZN(n1660) );
  AOI21_X1 U6369 ( .B1(n1660), .B2(n1659), .A(n138), .ZN(\unit_fetch/n447 ) );
  OAI21_X1 U6370 ( .B1(net141182), .B2(n124), .A(n1661), .ZN(
        \unit_fetch/unit_programCounter/ffi_6/n5 ) );
  OAI21_X1 U6371 ( .B1(net141182), .B2(n121), .A(n51), .ZN(
        \unit_fetch/unit_programCounter/ffi_7/n5 ) );
  OAI21_X1 U6372 ( .B1(net141182), .B2(n112), .A(n1663), .ZN(
        \unit_fetch/unit_programCounter/ffi_13/n5 ) );
  OAI21_X1 U6373 ( .B1(n81), .B2(net130308), .A(n1664), .ZN(
        \unit_fetch/unit_programCounter/ffi_2/n5 ) );
  INV_X1 U6374 ( .A(n123), .ZN(n1665) );
  NOR3_X1 U6375 ( .A1(n1665), .A2(n1693), .A3(n1695), .ZN(
        \unit_control/next_state[1] ) );
  NOR2_X1 U6376 ( .A1(n1666), .A2(n139), .ZN(
        \unit_control/uut_second_stage/ffi_24/n5 ) );
  INV_X1 U6377 ( .A(n1667), .ZN(n1668) );
  NAND2_X1 U6378 ( .A1(n1668), .A2(n141), .ZN(n1685) );
  INV_X1 U6379 ( .A(n1685), .ZN(\unit_control/uut_second_stage/ffi_15/n5 ) );
  NAND2_X1 U6380 ( .A1(\unit_control/uut_second_stage/ffi_15/n5 ), .A2(n1669), 
        .ZN(n1672) );
  NAND2_X1 U6381 ( .A1(n141), .A2(n1670), .ZN(n1690) );
  OAI21_X1 U6382 ( .B1(n1680), .B2(n1673), .A(n1686), .ZN(n1671) );
  NAND2_X1 U6383 ( .A1(n141), .A2(n1671), .ZN(n1691) );
  INV_X1 U6384 ( .A(n1686), .ZN(n1677) );
  INV_X1 U6385 ( .A(n1673), .ZN(n1683) );
  NOR2_X1 U6386 ( .A1(n1677), .A2(n1683), .ZN(n1675) );
  AOI21_X1 U6387 ( .B1(n1675), .B2(n1678), .A(n138), .ZN(
        \unit_control/uut_second_stage/ffi_9/n5 ) );
  NAND2_X1 U6388 ( .A1(n1676), .A2(n1679), .ZN(n1678) );
  NAND2_X1 U6389 ( .A1(n1677), .A2(n1680), .ZN(n1682) );
  AOI21_X1 U6390 ( .B1(n1678), .B2(n1682), .A(n140), .ZN(
        \unit_control/uut_second_stage/ffi_10/n5 ) );
  NOR4_X1 U6391 ( .A1(n140), .A2(n57), .A3(n1680), .A4(n1679), .ZN(
        \unit_control/uut_second_stage/ffi_11/n5 ) );
  NOR2_X1 U6392 ( .A1(n140), .A2(n1682), .ZN(
        \unit_control/uut_second_stage/ffi_12/n5 ) );
  OAI21_X1 U6393 ( .B1(n1688), .B2(n1683), .A(n141), .ZN(n1684) );
  NAND2_X1 U6394 ( .A1(n1685), .A2(n1684), .ZN(
        \unit_control/uut_second_stage/ffi_13/n5 ) );
  NOR2_X1 U6395 ( .A1(n138), .A2(n1686), .ZN(
        \unit_control/uut_second_stage/ffi_14/n5 ) );
  OAI21_X1 U6396 ( .B1(n1688), .B2(n1687), .A(n141), .ZN(n1689) );
  NAND2_X1 U6397 ( .A1(n1690), .A2(n1689), .ZN(
        \unit_control/uut_second_stage/ffi_17/n5 ) );
  INV_X1 U6398 ( .A(n1691), .ZN(\unit_control/n418 ) );
  INV_X1 U6399 ( .A(n1692), .ZN(n1696) );
  NOR4_X1 U6400 ( .A1(n1696), .A2(n1695), .A3(n123), .A4(n1693), .ZN(
        \unit_control/next_state[0] ) );
endmodule

