
module register_file_WORD_SIZE32_ADDR_SIZE5 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n2163), .CK(CLK), .Q(\REGISTERS[0][31] )
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n2162), .CK(CLK), .Q(\REGISTERS[0][30] )
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n2161), .CK(CLK), .Q(\REGISTERS[0][29] )
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n2160), .CK(CLK), .Q(\REGISTERS[0][28] )
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n2159), .CK(CLK), .Q(\REGISTERS[0][27] )
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n2158), .CK(CLK), .Q(\REGISTERS[0][26] )
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n2157), .CK(CLK), .Q(\REGISTERS[0][25] )
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n2156), .CK(CLK), .Q(\REGISTERS[0][24] )
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n2155), .CK(CLK), .Q(\REGISTERS[0][23] )
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n2154), .CK(CLK), .Q(\REGISTERS[0][22] )
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n2153), .CK(CLK), .Q(\REGISTERS[0][21] )
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n2152), .CK(CLK), .Q(\REGISTERS[0][20] )
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n2151), .CK(CLK), .Q(\REGISTERS[0][19] )
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n2150), .CK(CLK), .Q(\REGISTERS[0][18] )
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n2149), .CK(CLK), .Q(\REGISTERS[0][17] )
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n2148), .CK(CLK), .Q(\REGISTERS[0][16] )
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n2147), .CK(CLK), .Q(\REGISTERS[0][15] )
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n2146), .CK(CLK), .Q(\REGISTERS[0][14] )
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n2145), .CK(CLK), .Q(\REGISTERS[0][13] )
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n2144), .CK(CLK), .Q(\REGISTERS[0][12] )
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n2143), .CK(CLK), .Q(\REGISTERS[0][11] )
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n2142), .CK(CLK), .Q(\REGISTERS[0][10] )
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n2141), .CK(CLK), .Q(\REGISTERS[0][9] ) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n2140), .CK(CLK), .Q(\REGISTERS[0][8] ) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n2139), .CK(CLK), .Q(\REGISTERS[0][7] ) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n2138), .CK(CLK), .Q(\REGISTERS[0][6] ) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n2137), .CK(CLK), .Q(\REGISTERS[0][5] ) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n2136), .CK(CLK), .Q(\REGISTERS[0][4] ) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n2135), .CK(CLK), .Q(\REGISTERS[0][3] ) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n2134), .CK(CLK), .Q(\REGISTERS[0][2] ) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n2133), .CK(CLK), .Q(\REGISTERS[0][1] ) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n2132), .CK(CLK), .Q(\REGISTERS[0][0] ) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n2131), .CK(CLK), .Q(\REGISTERS[1][31] )
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n2130), .CK(CLK), .Q(\REGISTERS[1][30] )
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n2129), .CK(CLK), .Q(\REGISTERS[1][29] )
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n2128), .CK(CLK), .Q(\REGISTERS[1][28] )
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n2127), .CK(CLK), .Q(\REGISTERS[1][27] )
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n2126), .CK(CLK), .Q(\REGISTERS[1][26] )
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n2125), .CK(CLK), .Q(\REGISTERS[1][25] )
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n2124), .CK(CLK), .Q(\REGISTERS[1][24] )
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n2123), .CK(CLK), .Q(\REGISTERS[1][23] )
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n2122), .CK(CLK), .Q(\REGISTERS[1][22] )
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n2121), .CK(CLK), .Q(\REGISTERS[1][21] )
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n2120), .CK(CLK), .Q(\REGISTERS[1][20] )
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n2119), .CK(CLK), .Q(\REGISTERS[1][19] )
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n2118), .CK(CLK), .Q(\REGISTERS[1][18] )
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n2117), .CK(CLK), .Q(\REGISTERS[1][17] )
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n2116), .CK(CLK), .Q(\REGISTERS[1][16] )
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n2115), .CK(CLK), .Q(\REGISTERS[1][15] )
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n2114), .CK(CLK), .Q(\REGISTERS[1][14] )
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n2113), .CK(CLK), .Q(\REGISTERS[1][13] )
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n2112), .CK(CLK), .Q(\REGISTERS[1][12] )
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n2111), .CK(CLK), .Q(\REGISTERS[1][11] )
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n2110), .CK(CLK), .Q(\REGISTERS[1][10] )
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n2109), .CK(CLK), .Q(\REGISTERS[1][9] ) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n2108), .CK(CLK), .Q(\REGISTERS[1][8] ) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n2107), .CK(CLK), .Q(\REGISTERS[1][7] ) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n2106), .CK(CLK), .Q(\REGISTERS[1][6] ) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n2105), .CK(CLK), .Q(\REGISTERS[1][5] ) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n2104), .CK(CLK), .Q(\REGISTERS[1][4] ) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n2103), .CK(CLK), .Q(\REGISTERS[1][3] ) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n2102), .CK(CLK), .Q(\REGISTERS[1][2] ) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n2101), .CK(CLK), .Q(\REGISTERS[1][1] ) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n2100), .CK(CLK), .Q(\REGISTERS[1][0] ) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n2099), .CK(CLK), .Q(\REGISTERS[2][31] )
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n2098), .CK(CLK), .Q(\REGISTERS[2][30] )
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n2097), .CK(CLK), .Q(\REGISTERS[2][29] )
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n2096), .CK(CLK), .Q(\REGISTERS[2][28] )
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n2095), .CK(CLK), .Q(\REGISTERS[2][27] )
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n2094), .CK(CLK), .Q(\REGISTERS[2][26] )
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n2093), .CK(CLK), .Q(\REGISTERS[2][25] )
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n2092), .CK(CLK), .Q(\REGISTERS[2][24] )
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n2091), .CK(CLK), .Q(\REGISTERS[2][23] )
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n2090), .CK(CLK), .Q(\REGISTERS[2][22] )
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n2089), .CK(CLK), .Q(\REGISTERS[2][21] )
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n2088), .CK(CLK), .Q(\REGISTERS[2][20] )
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n2087), .CK(CLK), .Q(\REGISTERS[2][19] )
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n2086), .CK(CLK), .Q(\REGISTERS[2][18] )
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n2085), .CK(CLK), .Q(\REGISTERS[2][17] )
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n2084), .CK(CLK), .Q(\REGISTERS[2][16] )
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n2083), .CK(CLK), .Q(\REGISTERS[2][15] )
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n2082), .CK(CLK), .Q(\REGISTERS[2][14] )
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n2081), .CK(CLK), .Q(\REGISTERS[2][13] )
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n2080), .CK(CLK), .Q(\REGISTERS[2][12] )
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n2079), .CK(CLK), .Q(\REGISTERS[2][11] )
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n2078), .CK(CLK), .Q(\REGISTERS[2][10] )
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n2077), .CK(CLK), .Q(\REGISTERS[2][9] ) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n2076), .CK(CLK), .Q(\REGISTERS[2][8] ) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n2075), .CK(CLK), .Q(\REGISTERS[2][7] ) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n2074), .CK(CLK), .Q(\REGISTERS[2][6] ) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n2073), .CK(CLK), .Q(\REGISTERS[2][5] ) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n2072), .CK(CLK), .Q(\REGISTERS[2][4] ) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n2071), .CK(CLK), .Q(\REGISTERS[2][3] ) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n2070), .CK(CLK), .Q(\REGISTERS[2][2] ) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n2069), .CK(CLK), .Q(\REGISTERS[2][1] ) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n2068), .CK(CLK), .Q(\REGISTERS[2][0] ) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n2067), .CK(CLK), .Q(\REGISTERS[3][31] )
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n2066), .CK(CLK), .Q(\REGISTERS[3][30] )
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n2065), .CK(CLK), .Q(\REGISTERS[3][29] )
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n2064), .CK(CLK), .Q(\REGISTERS[3][28] )
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n2063), .CK(CLK), .Q(\REGISTERS[3][27] )
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n2062), .CK(CLK), .Q(\REGISTERS[3][26] )
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n2061), .CK(CLK), .Q(\REGISTERS[3][25] )
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n2060), .CK(CLK), .Q(\REGISTERS[3][24] )
         );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n2059), .CK(CLK), .Q(\REGISTERS[3][23] )
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n2058), .CK(CLK), .Q(\REGISTERS[3][22] )
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n2057), .CK(CLK), .Q(\REGISTERS[3][21] )
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n2056), .CK(CLK), .Q(\REGISTERS[3][20] )
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n2055), .CK(CLK), .Q(\REGISTERS[3][19] )
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n2054), .CK(CLK), .Q(\REGISTERS[3][18] )
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n2053), .CK(CLK), .Q(\REGISTERS[3][17] )
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n2052), .CK(CLK), .Q(\REGISTERS[3][16] )
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n2051), .CK(CLK), .Q(\REGISTERS[3][15] )
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n2050), .CK(CLK), .Q(\REGISTERS[3][14] )
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n2049), .CK(CLK), .Q(\REGISTERS[3][13] )
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n2048), .CK(CLK), .Q(\REGISTERS[3][12] )
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n2047), .CK(CLK), .Q(\REGISTERS[3][11] )
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n2046), .CK(CLK), .Q(\REGISTERS[3][10] )
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n2045), .CK(CLK), .Q(\REGISTERS[3][9] ) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n2044), .CK(CLK), .Q(\REGISTERS[3][8] ) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n2043), .CK(CLK), .Q(\REGISTERS[3][7] ) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n2042), .CK(CLK), .Q(\REGISTERS[3][6] ) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n2041), .CK(CLK), .Q(\REGISTERS[3][5] ) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n2040), .CK(CLK), .Q(\REGISTERS[3][4] ) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n2039), .CK(CLK), .Q(\REGISTERS[3][3] ) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n2038), .CK(CLK), .Q(\REGISTERS[3][2] ) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n2037), .CK(CLK), .Q(\REGISTERS[3][1] ) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n2036), .CK(CLK), .Q(\REGISTERS[3][0] ) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n2035), .CK(CLK), .Q(\REGISTERS[4][31] )
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n2034), .CK(CLK), .Q(\REGISTERS[4][30] )
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n2033), .CK(CLK), .Q(\REGISTERS[4][29] )
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n2032), .CK(CLK), .Q(\REGISTERS[4][28] )
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n2031), .CK(CLK), .Q(\REGISTERS[4][27] )
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n2030), .CK(CLK), .Q(\REGISTERS[4][26] )
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n2029), .CK(CLK), .Q(\REGISTERS[4][25] )
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n2028), .CK(CLK), .Q(\REGISTERS[4][24] )
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n2027), .CK(CLK), .Q(\REGISTERS[4][23] )
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n2026), .CK(CLK), .Q(\REGISTERS[4][22] )
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n2025), .CK(CLK), .Q(\REGISTERS[4][21] )
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n2024), .CK(CLK), .Q(\REGISTERS[4][20] )
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n2023), .CK(CLK), .Q(\REGISTERS[4][19] )
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n2022), .CK(CLK), .Q(\REGISTERS[4][18] )
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n2021), .CK(CLK), .Q(\REGISTERS[4][17] )
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n2020), .CK(CLK), .Q(\REGISTERS[4][16] )
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n2019), .CK(CLK), .Q(\REGISTERS[4][15] )
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n2018), .CK(CLK), .Q(\REGISTERS[4][14] )
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n2017), .CK(CLK), .Q(\REGISTERS[4][13] )
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n2016), .CK(CLK), .Q(\REGISTERS[4][12] )
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n2015), .CK(CLK), .Q(\REGISTERS[4][11] )
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n2014), .CK(CLK), .Q(\REGISTERS[4][10] )
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n2013), .CK(CLK), .Q(\REGISTERS[4][9] ) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n2012), .CK(CLK), .Q(\REGISTERS[4][8] ) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n2011), .CK(CLK), .Q(\REGISTERS[4][7] ) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n2010), .CK(CLK), .Q(\REGISTERS[4][6] ) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n2009), .CK(CLK), .Q(\REGISTERS[4][5] ) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n2008), .CK(CLK), .Q(\REGISTERS[4][4] ) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n2007), .CK(CLK), .Q(\REGISTERS[4][3] ) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n2006), .CK(CLK), .Q(\REGISTERS[4][2] ) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n2005), .CK(CLK), .Q(\REGISTERS[4][1] ) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n2004), .CK(CLK), .Q(\REGISTERS[4][0] ) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n2003), .CK(CLK), .Q(\REGISTERS[5][31] )
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n2002), .CK(CLK), .Q(\REGISTERS[5][30] )
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n2001), .CK(CLK), .Q(\REGISTERS[5][29] )
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n2000), .CK(CLK), .Q(\REGISTERS[5][28] )
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n1999), .CK(CLK), .Q(\REGISTERS[5][27] )
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n1998), .CK(CLK), .Q(\REGISTERS[5][26] )
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n1997), .CK(CLK), .Q(\REGISTERS[5][25] )
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n1996), .CK(CLK), .Q(\REGISTERS[5][24] )
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n1995), .CK(CLK), .Q(\REGISTERS[5][23] )
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n1994), .CK(CLK), .Q(\REGISTERS[5][22] )
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n1993), .CK(CLK), .Q(\REGISTERS[5][21] )
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n1992), .CK(CLK), .Q(\REGISTERS[5][20] )
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n1991), .CK(CLK), .Q(\REGISTERS[5][19] )
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n1990), .CK(CLK), .Q(\REGISTERS[5][18] )
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n1989), .CK(CLK), .Q(\REGISTERS[5][17] )
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n1988), .CK(CLK), .Q(\REGISTERS[5][16] )
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n1987), .CK(CLK), .Q(\REGISTERS[5][15] )
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n1986), .CK(CLK), .Q(\REGISTERS[5][14] )
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n1985), .CK(CLK), .Q(\REGISTERS[5][13] )
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n1984), .CK(CLK), .Q(\REGISTERS[5][12] )
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n1983), .CK(CLK), .Q(\REGISTERS[5][11] )
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n1982), .CK(CLK), .Q(\REGISTERS[5][10] )
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n1981), .CK(CLK), .Q(\REGISTERS[5][9] ) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n1980), .CK(CLK), .Q(\REGISTERS[5][8] ) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n1979), .CK(CLK), .Q(\REGISTERS[5][7] ) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n1978), .CK(CLK), .Q(\REGISTERS[5][6] ) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n1977), .CK(CLK), .Q(\REGISTERS[5][5] ) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n1976), .CK(CLK), .Q(\REGISTERS[5][4] ) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n1975), .CK(CLK), .Q(\REGISTERS[5][3] ) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n1974), .CK(CLK), .Q(\REGISTERS[5][2] ) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n1973), .CK(CLK), .Q(\REGISTERS[5][1] ) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n1972), .CK(CLK), .Q(\REGISTERS[5][0] ) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n1971), .CK(CLK), .Q(\REGISTERS[6][31] )
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n1970), .CK(CLK), .Q(\REGISTERS[6][30] )
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n1969), .CK(CLK), .Q(\REGISTERS[6][29] )
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n1968), .CK(CLK), .Q(\REGISTERS[6][28] )
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n1967), .CK(CLK), .Q(\REGISTERS[6][27] )
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n1966), .CK(CLK), .Q(\REGISTERS[6][26] )
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n1965), .CK(CLK), .Q(\REGISTERS[6][25] )
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n1964), .CK(CLK), .Q(\REGISTERS[6][24] )
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n1963), .CK(CLK), .Q(\REGISTERS[6][23] )
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n1962), .CK(CLK), .Q(\REGISTERS[6][22] )
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n1961), .CK(CLK), .Q(\REGISTERS[6][21] )
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n1960), .CK(CLK), .Q(\REGISTERS[6][20] )
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n1959), .CK(CLK), .Q(\REGISTERS[6][19] )
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n1958), .CK(CLK), .Q(\REGISTERS[6][18] )
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n1957), .CK(CLK), .Q(\REGISTERS[6][17] )
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n1956), .CK(CLK), .Q(\REGISTERS[6][16] )
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n1955), .CK(CLK), .Q(\REGISTERS[6][15] )
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n1954), .CK(CLK), .Q(\REGISTERS[6][14] )
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n1953), .CK(CLK), .Q(\REGISTERS[6][13] )
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n1952), .CK(CLK), .Q(\REGISTERS[6][12] )
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n1951), .CK(CLK), .Q(\REGISTERS[6][11] )
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n1950), .CK(CLK), .Q(\REGISTERS[6][10] )
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n1949), .CK(CLK), .Q(\REGISTERS[6][9] ) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n1948), .CK(CLK), .Q(\REGISTERS[6][8] ) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n1947), .CK(CLK), .Q(\REGISTERS[6][7] ) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n1946), .CK(CLK), .Q(\REGISTERS[6][6] ) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n1945), .CK(CLK), .Q(\REGISTERS[6][5] ) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n1944), .CK(CLK), .Q(\REGISTERS[6][4] ) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n1943), .CK(CLK), .Q(\REGISTERS[6][3] ) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n1942), .CK(CLK), .Q(\REGISTERS[6][2] ) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n1941), .CK(CLK), .Q(\REGISTERS[6][1] ) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n1940), .CK(CLK), .Q(\REGISTERS[6][0] ) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n1939), .CK(CLK), .Q(\REGISTERS[7][31] )
         );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n1938), .CK(CLK), .Q(\REGISTERS[7][30] )
         );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n1937), .CK(CLK), .Q(\REGISTERS[7][29] )
         );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n1936), .CK(CLK), .Q(\REGISTERS[7][28] )
         );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n1935), .CK(CLK), .Q(\REGISTERS[7][27] )
         );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n1934), .CK(CLK), .Q(\REGISTERS[7][26] )
         );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n1933), .CK(CLK), .Q(\REGISTERS[7][25] )
         );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n1932), .CK(CLK), .Q(\REGISTERS[7][24] )
         );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n1931), .CK(CLK), .Q(\REGISTERS[7][23] )
         );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n1930), .CK(CLK), .Q(\REGISTERS[7][22] )
         );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n1929), .CK(CLK), .Q(\REGISTERS[7][21] )
         );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n1928), .CK(CLK), .Q(\REGISTERS[7][20] )
         );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n1927), .CK(CLK), .Q(\REGISTERS[7][19] )
         );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n1926), .CK(CLK), .Q(\REGISTERS[7][18] )
         );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n1925), .CK(CLK), .Q(\REGISTERS[7][17] )
         );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n1924), .CK(CLK), .Q(\REGISTERS[7][16] )
         );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n1923), .CK(CLK), .Q(\REGISTERS[7][15] )
         );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n1922), .CK(CLK), .Q(\REGISTERS[7][14] )
         );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n1921), .CK(CLK), .Q(\REGISTERS[7][13] )
         );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n1920), .CK(CLK), .Q(\REGISTERS[7][12] )
         );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n1919), .CK(CLK), .Q(\REGISTERS[7][11] )
         );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n1918), .CK(CLK), .Q(\REGISTERS[7][10] )
         );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n1917), .CK(CLK), .Q(\REGISTERS[7][9] ) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n1916), .CK(CLK), .Q(\REGISTERS[7][8] ) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n1915), .CK(CLK), .Q(\REGISTERS[7][7] ) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n1914), .CK(CLK), .Q(\REGISTERS[7][6] ) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n1913), .CK(CLK), .Q(\REGISTERS[7][5] ) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n1912), .CK(CLK), .Q(\REGISTERS[7][4] ) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n1911), .CK(CLK), .Q(\REGISTERS[7][3] ) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n1910), .CK(CLK), .Q(\REGISTERS[7][2] ) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n1909), .CK(CLK), .Q(\REGISTERS[7][1] ) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n1908), .CK(CLK), .Q(\REGISTERS[7][0] ) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n1907), .CK(CLK), .Q(\REGISTERS[8][31] )
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n1906), .CK(CLK), .Q(\REGISTERS[8][30] )
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n1905), .CK(CLK), .Q(\REGISTERS[8][29] )
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n1904), .CK(CLK), .Q(\REGISTERS[8][28] )
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n1903), .CK(CLK), .Q(\REGISTERS[8][27] )
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n1902), .CK(CLK), .Q(\REGISTERS[8][26] )
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n1901), .CK(CLK), .Q(\REGISTERS[8][25] )
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n1900), .CK(CLK), .Q(\REGISTERS[8][24] )
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n1899), .CK(CLK), .Q(\REGISTERS[8][23] )
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n1898), .CK(CLK), .Q(\REGISTERS[8][22] )
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n1897), .CK(CLK), .Q(\REGISTERS[8][21] )
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n1896), .CK(CLK), .Q(\REGISTERS[8][20] )
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n1895), .CK(CLK), .Q(\REGISTERS[8][19] )
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n1894), .CK(CLK), .Q(\REGISTERS[8][18] )
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n1893), .CK(CLK), .Q(\REGISTERS[8][17] )
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n1892), .CK(CLK), .Q(\REGISTERS[8][16] )
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n1891), .CK(CLK), .Q(\REGISTERS[8][15] )
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n1890), .CK(CLK), .Q(\REGISTERS[8][14] )
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n1889), .CK(CLK), .Q(\REGISTERS[8][13] )
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n1888), .CK(CLK), .Q(\REGISTERS[8][12] )
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n1887), .CK(CLK), .Q(\REGISTERS[8][11] )
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n1886), .CK(CLK), .Q(\REGISTERS[8][10] )
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n1885), .CK(CLK), .Q(\REGISTERS[8][9] ) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n1884), .CK(CLK), .Q(\REGISTERS[8][8] ) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n1883), .CK(CLK), .Q(\REGISTERS[8][7] ) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n1882), .CK(CLK), .Q(\REGISTERS[8][6] ) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n1881), .CK(CLK), .Q(\REGISTERS[8][5] ) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n1880), .CK(CLK), .Q(\REGISTERS[8][4] ) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n1879), .CK(CLK), .Q(\REGISTERS[8][3] ) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n1878), .CK(CLK), .Q(\REGISTERS[8][2] ) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n1877), .CK(CLK), .Q(\REGISTERS[8][1] ) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n1876), .CK(CLK), .Q(\REGISTERS[8][0] ) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n1875), .CK(CLK), .Q(\REGISTERS[9][31] )
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n1874), .CK(CLK), .Q(\REGISTERS[9][30] )
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n1873), .CK(CLK), .Q(\REGISTERS[9][29] )
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n1872), .CK(CLK), .Q(\REGISTERS[9][28] )
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n1871), .CK(CLK), .Q(\REGISTERS[9][27] )
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n1870), .CK(CLK), .Q(\REGISTERS[9][26] )
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n1869), .CK(CLK), .Q(\REGISTERS[9][25] )
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n1868), .CK(CLK), .Q(\REGISTERS[9][24] )
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n1867), .CK(CLK), .Q(\REGISTERS[9][23] )
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n1866), .CK(CLK), .Q(\REGISTERS[9][22] )
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n1865), .CK(CLK), .Q(\REGISTERS[9][21] )
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n1864), .CK(CLK), .Q(\REGISTERS[9][20] )
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n1863), .CK(CLK), .Q(\REGISTERS[9][19] )
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n1862), .CK(CLK), .Q(\REGISTERS[9][18] )
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n1861), .CK(CLK), .Q(\REGISTERS[9][17] )
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n1860), .CK(CLK), .Q(\REGISTERS[9][16] )
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n1859), .CK(CLK), .Q(\REGISTERS[9][15] )
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n1858), .CK(CLK), .Q(\REGISTERS[9][14] )
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n1857), .CK(CLK), .Q(\REGISTERS[9][13] )
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n1856), .CK(CLK), .Q(\REGISTERS[9][12] )
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n1855), .CK(CLK), .Q(\REGISTERS[9][11] )
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n1854), .CK(CLK), .Q(\REGISTERS[9][10] )
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n1853), .CK(CLK), .Q(\REGISTERS[9][9] ) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n1852), .CK(CLK), .Q(\REGISTERS[9][8] ) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n1851), .CK(CLK), .Q(\REGISTERS[9][7] ) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n1850), .CK(CLK), .Q(\REGISTERS[9][6] ) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n1849), .CK(CLK), .Q(\REGISTERS[9][5] ) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n1848), .CK(CLK), .Q(\REGISTERS[9][4] ) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n1847), .CK(CLK), .Q(\REGISTERS[9][3] ) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n1846), .CK(CLK), .Q(\REGISTERS[9][2] ) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n1845), .CK(CLK), .Q(\REGISTERS[9][1] ) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n1844), .CK(CLK), .Q(\REGISTERS[9][0] ) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n1843), .CK(CLK), .Q(\REGISTERS[10][31] ) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n1842), .CK(CLK), .Q(\REGISTERS[10][30] ) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n1841), .CK(CLK), .Q(\REGISTERS[10][29] ) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n1840), .CK(CLK), .Q(\REGISTERS[10][28] ) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n1839), .CK(CLK), .Q(\REGISTERS[10][27] ) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n1838), .CK(CLK), .Q(\REGISTERS[10][26] ) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n1837), .CK(CLK), .Q(\REGISTERS[10][25] ) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n1836), .CK(CLK), .Q(\REGISTERS[10][24] ) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n1835), .CK(CLK), .Q(\REGISTERS[10][23] ) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n1834), .CK(CLK), .Q(\REGISTERS[10][22] ) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n1833), .CK(CLK), .Q(\REGISTERS[10][21] ) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n1832), .CK(CLK), .Q(\REGISTERS[10][20] ) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n1831), .CK(CLK), .Q(\REGISTERS[10][19] ) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n1830), .CK(CLK), .Q(\REGISTERS[10][18] ) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n1829), .CK(CLK), .Q(\REGISTERS[10][17] ) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n1828), .CK(CLK), .Q(\REGISTERS[10][16] ) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n1827), .CK(CLK), .Q(\REGISTERS[10][15] ) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n1826), .CK(CLK), .Q(\REGISTERS[10][14] ) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n1825), .CK(CLK), .Q(\REGISTERS[10][13] ) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n1824), .CK(CLK), .Q(\REGISTERS[10][12] ) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n1823), .CK(CLK), .Q(\REGISTERS[10][11] ) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n1822), .CK(CLK), .Q(\REGISTERS[10][10] ) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n1821), .CK(CLK), .Q(\REGISTERS[10][9] )
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n1820), .CK(CLK), .Q(\REGISTERS[10][8] )
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n1819), .CK(CLK), .Q(\REGISTERS[10][7] )
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n1818), .CK(CLK), .Q(\REGISTERS[10][6] )
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n1817), .CK(CLK), .Q(\REGISTERS[10][5] )
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n1816), .CK(CLK), .Q(\REGISTERS[10][4] )
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n1815), .CK(CLK), .Q(\REGISTERS[10][3] )
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n1814), .CK(CLK), .Q(\REGISTERS[10][2] )
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n1813), .CK(CLK), .Q(\REGISTERS[10][1] )
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n1812), .CK(CLK), .Q(\REGISTERS[10][0] )
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n1811), .CK(CLK), .Q(\REGISTERS[11][31] ) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n1810), .CK(CLK), .Q(\REGISTERS[11][30] ) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n1809), .CK(CLK), .Q(\REGISTERS[11][29] ) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n1808), .CK(CLK), .Q(\REGISTERS[11][28] ) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n1807), .CK(CLK), .Q(\REGISTERS[11][27] ) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n1806), .CK(CLK), .Q(\REGISTERS[11][26] ) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n1805), .CK(CLK), .Q(\REGISTERS[11][25] ) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n1804), .CK(CLK), .Q(\REGISTERS[11][24] ) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n1803), .CK(CLK), .Q(\REGISTERS[11][23] ) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n1802), .CK(CLK), .Q(\REGISTERS[11][22] ) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n1801), .CK(CLK), .Q(\REGISTERS[11][21] ) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n1800), .CK(CLK), .Q(\REGISTERS[11][20] ) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n1799), .CK(CLK), .Q(\REGISTERS[11][19] ) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n1798), .CK(CLK), .Q(\REGISTERS[11][18] ) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n1797), .CK(CLK), .Q(\REGISTERS[11][17] ) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n1796), .CK(CLK), .Q(\REGISTERS[11][16] ) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n1795), .CK(CLK), .Q(\REGISTERS[11][15] ) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n1794), .CK(CLK), .Q(\REGISTERS[11][14] ) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n1793), .CK(CLK), .Q(\REGISTERS[11][13] ) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n1792), .CK(CLK), .Q(\REGISTERS[11][12] ) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n1791), .CK(CLK), .Q(\REGISTERS[11][11] ) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n1790), .CK(CLK), .Q(\REGISTERS[11][10] ) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n1789), .CK(CLK), .Q(\REGISTERS[11][9] )
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n1788), .CK(CLK), .Q(\REGISTERS[11][8] )
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n1787), .CK(CLK), .Q(\REGISTERS[11][7] )
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n1786), .CK(CLK), .Q(\REGISTERS[11][6] )
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n1785), .CK(CLK), .Q(\REGISTERS[11][5] )
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n1784), .CK(CLK), .Q(\REGISTERS[11][4] )
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n1783), .CK(CLK), .Q(\REGISTERS[11][3] )
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n1782), .CK(CLK), .Q(\REGISTERS[11][2] )
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n1781), .CK(CLK), .Q(\REGISTERS[11][1] )
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n1780), .CK(CLK), .Q(\REGISTERS[11][0] )
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n1779), .CK(CLK), .Q(\REGISTERS[12][31] ) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n1778), .CK(CLK), .Q(\REGISTERS[12][30] ) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n1777), .CK(CLK), .Q(\REGISTERS[12][29] ) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n1776), .CK(CLK), .Q(\REGISTERS[12][28] ) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n1775), .CK(CLK), .Q(\REGISTERS[12][27] ) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n1774), .CK(CLK), .Q(\REGISTERS[12][26] ) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n1773), .CK(CLK), .Q(\REGISTERS[12][25] ) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n1772), .CK(CLK), .Q(\REGISTERS[12][24] ) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n1771), .CK(CLK), .Q(\REGISTERS[12][23] ) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n1770), .CK(CLK), .Q(\REGISTERS[12][22] ) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n1769), .CK(CLK), .Q(\REGISTERS[12][21] ) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n1768), .CK(CLK), .Q(\REGISTERS[12][20] ) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n1767), .CK(CLK), .Q(\REGISTERS[12][19] ) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n1766), .CK(CLK), .Q(\REGISTERS[12][18] ) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n1765), .CK(CLK), .Q(\REGISTERS[12][17] ) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n1764), .CK(CLK), .Q(\REGISTERS[12][16] ) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n1763), .CK(CLK), .Q(\REGISTERS[12][15] ) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n1762), .CK(CLK), .Q(\REGISTERS[12][14] ) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n1761), .CK(CLK), .Q(\REGISTERS[12][13] ) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n1760), .CK(CLK), .Q(\REGISTERS[12][12] ) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n1759), .CK(CLK), .Q(\REGISTERS[12][11] ) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n1758), .CK(CLK), .Q(\REGISTERS[12][10] ) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n1757), .CK(CLK), .Q(\REGISTERS[12][9] )
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n1756), .CK(CLK), .Q(\REGISTERS[12][8] )
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n1755), .CK(CLK), .Q(\REGISTERS[12][7] )
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n1754), .CK(CLK), .Q(\REGISTERS[12][6] )
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n1753), .CK(CLK), .Q(\REGISTERS[12][5] )
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n1752), .CK(CLK), .Q(\REGISTERS[12][4] )
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n1751), .CK(CLK), .Q(\REGISTERS[12][3] )
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n1750), .CK(CLK), .Q(\REGISTERS[12][2] )
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n1749), .CK(CLK), .Q(\REGISTERS[12][1] )
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n1748), .CK(CLK), .Q(\REGISTERS[12][0] )
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n1747), .CK(CLK), .Q(\REGISTERS[13][31] ) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n1746), .CK(CLK), .Q(\REGISTERS[13][30] ) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n1745), .CK(CLK), .Q(\REGISTERS[13][29] ) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n1744), .CK(CLK), .Q(\REGISTERS[13][28] ) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n1743), .CK(CLK), .Q(\REGISTERS[13][27] ) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n1742), .CK(CLK), .Q(\REGISTERS[13][26] ) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n1741), .CK(CLK), .Q(\REGISTERS[13][25] ) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n1740), .CK(CLK), .Q(\REGISTERS[13][24] ) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n1739), .CK(CLK), .Q(\REGISTERS[13][23] ) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n1738), .CK(CLK), .Q(\REGISTERS[13][22] ) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n1737), .CK(CLK), .Q(\REGISTERS[13][21] ) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n1736), .CK(CLK), .Q(\REGISTERS[13][20] ) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n1735), .CK(CLK), .Q(\REGISTERS[13][19] ) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n1734), .CK(CLK), .Q(\REGISTERS[13][18] ) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n1733), .CK(CLK), .Q(\REGISTERS[13][17] ) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n1732), .CK(CLK), .Q(\REGISTERS[13][16] ) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n1731), .CK(CLK), .Q(\REGISTERS[13][15] ) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n1730), .CK(CLK), .Q(\REGISTERS[13][14] ) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n1729), .CK(CLK), .Q(\REGISTERS[13][13] ) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n1728), .CK(CLK), .Q(\REGISTERS[13][12] ) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n1727), .CK(CLK), .Q(\REGISTERS[13][11] ) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n1726), .CK(CLK), .Q(\REGISTERS[13][10] ) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n1725), .CK(CLK), .Q(\REGISTERS[13][9] )
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n1724), .CK(CLK), .Q(\REGISTERS[13][8] )
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n1723), .CK(CLK), .Q(\REGISTERS[13][7] )
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n1722), .CK(CLK), .Q(\REGISTERS[13][6] )
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n1721), .CK(CLK), .Q(\REGISTERS[13][5] )
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n1720), .CK(CLK), .Q(\REGISTERS[13][4] )
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n1719), .CK(CLK), .Q(\REGISTERS[13][3] )
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n1718), .CK(CLK), .Q(\REGISTERS[13][2] )
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n1717), .CK(CLK), .Q(\REGISTERS[13][1] )
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n1716), .CK(CLK), .Q(\REGISTERS[13][0] )
         );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n1715), .CK(CLK), .Q(\REGISTERS[14][31] ) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n1714), .CK(CLK), .Q(\REGISTERS[14][30] ) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n1713), .CK(CLK), .Q(\REGISTERS[14][29] ) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n1712), .CK(CLK), .Q(\REGISTERS[14][28] ) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n1711), .CK(CLK), .Q(\REGISTERS[14][27] ) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n1710), .CK(CLK), .Q(\REGISTERS[14][26] ) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n1709), .CK(CLK), .Q(\REGISTERS[14][25] ) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n1708), .CK(CLK), .Q(\REGISTERS[14][24] ) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n1707), .CK(CLK), .Q(\REGISTERS[14][23] ) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n1706), .CK(CLK), .Q(\REGISTERS[14][22] ) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n1705), .CK(CLK), .Q(\REGISTERS[14][21] ) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n1704), .CK(CLK), .Q(\REGISTERS[14][20] ) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n1703), .CK(CLK), .Q(\REGISTERS[14][19] ) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n1702), .CK(CLK), .Q(\REGISTERS[14][18] ) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n1701), .CK(CLK), .Q(\REGISTERS[14][17] ) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n1700), .CK(CLK), .Q(\REGISTERS[14][16] ) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n1699), .CK(CLK), .Q(\REGISTERS[14][15] ) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n1698), .CK(CLK), .Q(\REGISTERS[14][14] ) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n1697), .CK(CLK), .Q(\REGISTERS[14][13] ) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n1696), .CK(CLK), .Q(\REGISTERS[14][12] ) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n1695), .CK(CLK), .Q(\REGISTERS[14][11] ) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n1694), .CK(CLK), .Q(\REGISTERS[14][10] ) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n1693), .CK(CLK), .Q(\REGISTERS[14][9] )
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n1692), .CK(CLK), .Q(\REGISTERS[14][8] )
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n1691), .CK(CLK), .Q(\REGISTERS[14][7] )
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n1690), .CK(CLK), .Q(\REGISTERS[14][6] )
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n1689), .CK(CLK), .Q(\REGISTERS[14][5] )
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n1688), .CK(CLK), .Q(\REGISTERS[14][4] )
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n1687), .CK(CLK), .Q(\REGISTERS[14][3] )
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n1686), .CK(CLK), .Q(\REGISTERS[14][2] )
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n1685), .CK(CLK), .Q(\REGISTERS[14][1] )
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n1684), .CK(CLK), .Q(\REGISTERS[14][0] )
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n1683), .CK(CLK), .Q(\REGISTERS[15][31] ) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n1682), .CK(CLK), .Q(\REGISTERS[15][30] ) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n1681), .CK(CLK), .Q(\REGISTERS[15][29] ) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n1680), .CK(CLK), .Q(\REGISTERS[15][28] ) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n1679), .CK(CLK), .Q(\REGISTERS[15][27] ) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n1678), .CK(CLK), .Q(\REGISTERS[15][26] ) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n1677), .CK(CLK), .Q(\REGISTERS[15][25] ) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n1676), .CK(CLK), .Q(\REGISTERS[15][24] ) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n1675), .CK(CLK), .Q(\REGISTERS[15][23] ) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n1674), .CK(CLK), .Q(\REGISTERS[15][22] ) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n1673), .CK(CLK), .Q(\REGISTERS[15][21] ) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n1672), .CK(CLK), .Q(\REGISTERS[15][20] ) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n1671), .CK(CLK), .Q(\REGISTERS[15][19] ) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n1670), .CK(CLK), .Q(\REGISTERS[15][18] ) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n1669), .CK(CLK), .Q(\REGISTERS[15][17] ) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n1668), .CK(CLK), .Q(\REGISTERS[15][16] ) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n1667), .CK(CLK), .Q(\REGISTERS[15][15] ) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n1666), .CK(CLK), .Q(\REGISTERS[15][14] ) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n1665), .CK(CLK), .Q(\REGISTERS[15][13] ) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n1664), .CK(CLK), .Q(\REGISTERS[15][12] ) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n1663), .CK(CLK), .Q(\REGISTERS[15][11] ) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n1662), .CK(CLK), .Q(\REGISTERS[15][10] ) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n1661), .CK(CLK), .Q(\REGISTERS[15][9] )
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n1660), .CK(CLK), .Q(\REGISTERS[15][8] )
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n1659), .CK(CLK), .Q(\REGISTERS[15][7] )
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n1658), .CK(CLK), .Q(\REGISTERS[15][6] )
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n1657), .CK(CLK), .Q(\REGISTERS[15][5] )
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n1656), .CK(CLK), .Q(\REGISTERS[15][4] )
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n1655), .CK(CLK), .Q(\REGISTERS[15][3] )
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n1654), .CK(CLK), .Q(\REGISTERS[15][2] )
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n1653), .CK(CLK), .Q(\REGISTERS[15][1] )
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n1652), .CK(CLK), .Q(\REGISTERS[15][0] )
         );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n1651), .CK(CLK), .Q(\REGISTERS[16][31] ) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n1650), .CK(CLK), .Q(\REGISTERS[16][30] ) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n1649), .CK(CLK), .Q(\REGISTERS[16][29] ) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n1648), .CK(CLK), .Q(\REGISTERS[16][28] ) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n1647), .CK(CLK), .Q(\REGISTERS[16][27] ) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n1646), .CK(CLK), .Q(\REGISTERS[16][26] ) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n1645), .CK(CLK), .Q(\REGISTERS[16][25] ) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n1644), .CK(CLK), .Q(\REGISTERS[16][24] ) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n1643), .CK(CLK), .Q(\REGISTERS[16][23] ) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n1642), .CK(CLK), .Q(\REGISTERS[16][22] ) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n1641), .CK(CLK), .Q(\REGISTERS[16][21] ) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n1640), .CK(CLK), .Q(\REGISTERS[16][20] ) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n1639), .CK(CLK), .Q(\REGISTERS[16][19] ) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n1638), .CK(CLK), .Q(\REGISTERS[16][18] ) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n1637), .CK(CLK), .Q(\REGISTERS[16][17] ) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n1636), .CK(CLK), .Q(\REGISTERS[16][16] ) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n1635), .CK(CLK), .Q(\REGISTERS[16][15] ) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n1634), .CK(CLK), .Q(\REGISTERS[16][14] ) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n1633), .CK(CLK), .Q(\REGISTERS[16][13] ) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n1632), .CK(CLK), .Q(\REGISTERS[16][12] ) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n1631), .CK(CLK), .Q(\REGISTERS[16][11] ) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n1630), .CK(CLK), .Q(\REGISTERS[16][10] ) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n1629), .CK(CLK), .Q(\REGISTERS[16][9] )
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n1628), .CK(CLK), .Q(\REGISTERS[16][8] )
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n1627), .CK(CLK), .Q(\REGISTERS[16][7] )
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n1626), .CK(CLK), .Q(\REGISTERS[16][6] )
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n1625), .CK(CLK), .Q(\REGISTERS[16][5] )
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n1624), .CK(CLK), .Q(\REGISTERS[16][4] )
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n1623), .CK(CLK), .Q(\REGISTERS[16][3] )
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n1622), .CK(CLK), .Q(\REGISTERS[16][2] )
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n1621), .CK(CLK), .Q(\REGISTERS[16][1] )
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n1620), .CK(CLK), .Q(\REGISTERS[16][0] )
         );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n1619), .CK(CLK), .Q(\REGISTERS[17][31] ) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n1618), .CK(CLK), .Q(\REGISTERS[17][30] ) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n1617), .CK(CLK), .Q(\REGISTERS[17][29] ) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n1616), .CK(CLK), .Q(\REGISTERS[17][28] ) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n1615), .CK(CLK), .Q(\REGISTERS[17][27] ) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n1614), .CK(CLK), .Q(\REGISTERS[17][26] ) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n1613), .CK(CLK), .Q(\REGISTERS[17][25] ) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n1612), .CK(CLK), .Q(\REGISTERS[17][24] ) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n1611), .CK(CLK), .Q(\REGISTERS[17][23] ) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n1610), .CK(CLK), .Q(\REGISTERS[17][22] ) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n1609), .CK(CLK), .Q(\REGISTERS[17][21] ) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n1608), .CK(CLK), .Q(\REGISTERS[17][20] ) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n1607), .CK(CLK), .Q(\REGISTERS[17][19] ) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n1606), .CK(CLK), .Q(\REGISTERS[17][18] ) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n1605), .CK(CLK), .Q(\REGISTERS[17][17] ) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n1604), .CK(CLK), .Q(\REGISTERS[17][16] ) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n1603), .CK(CLK), .Q(\REGISTERS[17][15] ) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n1602), .CK(CLK), .Q(\REGISTERS[17][14] ) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n1601), .CK(CLK), .Q(\REGISTERS[17][13] ) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n1600), .CK(CLK), .Q(\REGISTERS[17][12] ) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n1599), .CK(CLK), .Q(\REGISTERS[17][11] ) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n1598), .CK(CLK), .Q(\REGISTERS[17][10] ) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n1597), .CK(CLK), .Q(\REGISTERS[17][9] )
         );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n1596), .CK(CLK), .Q(\REGISTERS[17][8] )
         );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n1595), .CK(CLK), .Q(\REGISTERS[17][7] )
         );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n1594), .CK(CLK), .Q(\REGISTERS[17][6] )
         );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n1593), .CK(CLK), .Q(\REGISTERS[17][5] )
         );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n1592), .CK(CLK), .Q(\REGISTERS[17][4] )
         );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n1591), .CK(CLK), .Q(\REGISTERS[17][3] )
         );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n1590), .CK(CLK), .Q(\REGISTERS[17][2] )
         );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n1589), .CK(CLK), .Q(\REGISTERS[17][1] )
         );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n1588), .CK(CLK), .Q(\REGISTERS[17][0] )
         );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n1587), .CK(CLK), .Q(\REGISTERS[18][31] ) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n1586), .CK(CLK), .Q(\REGISTERS[18][30] ) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n1585), .CK(CLK), .Q(\REGISTERS[18][29] ) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n1584), .CK(CLK), .Q(\REGISTERS[18][28] ) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n1583), .CK(CLK), .Q(\REGISTERS[18][27] ) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n1582), .CK(CLK), .Q(\REGISTERS[18][26] ) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n1581), .CK(CLK), .Q(\REGISTERS[18][25] ) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n1580), .CK(CLK), .Q(\REGISTERS[18][24] ) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n1579), .CK(CLK), .Q(\REGISTERS[18][23] ) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n1578), .CK(CLK), .Q(\REGISTERS[18][22] ) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n1577), .CK(CLK), .Q(\REGISTERS[18][21] ) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n1576), .CK(CLK), .Q(\REGISTERS[18][20] ) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n1575), .CK(CLK), .Q(\REGISTERS[18][19] ) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n1574), .CK(CLK), .Q(\REGISTERS[18][18] ) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n1573), .CK(CLK), .Q(\REGISTERS[18][17] ) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n1572), .CK(CLK), .Q(\REGISTERS[18][16] ) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n1571), .CK(CLK), .Q(\REGISTERS[18][15] ) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n1570), .CK(CLK), .Q(\REGISTERS[18][14] ) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n1569), .CK(CLK), .Q(\REGISTERS[18][13] ) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n1568), .CK(CLK), .Q(\REGISTERS[18][12] ) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n1567), .CK(CLK), .Q(\REGISTERS[18][11] ) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n1566), .CK(CLK), .Q(\REGISTERS[18][10] ) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n1565), .CK(CLK), .Q(\REGISTERS[18][9] )
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n1564), .CK(CLK), .Q(\REGISTERS[18][8] )
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n1563), .CK(CLK), .Q(\REGISTERS[18][7] )
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n1562), .CK(CLK), .Q(\REGISTERS[18][6] )
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n1561), .CK(CLK), .Q(\REGISTERS[18][5] )
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n1560), .CK(CLK), .Q(\REGISTERS[18][4] )
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n1559), .CK(CLK), .Q(\REGISTERS[18][3] )
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n1558), .CK(CLK), .Q(\REGISTERS[18][2] )
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n1557), .CK(CLK), .Q(\REGISTERS[18][1] )
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n1556), .CK(CLK), .Q(\REGISTERS[18][0] )
         );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n1555), .CK(CLK), .Q(\REGISTERS[19][31] ) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n1554), .CK(CLK), .Q(\REGISTERS[19][30] ) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n1553), .CK(CLK), .Q(\REGISTERS[19][29] ) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n1552), .CK(CLK), .Q(\REGISTERS[19][28] ) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n1551), .CK(CLK), .Q(\REGISTERS[19][27] ) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n1550), .CK(CLK), .Q(\REGISTERS[19][26] ) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n1549), .CK(CLK), .Q(\REGISTERS[19][25] ) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n1548), .CK(CLK), .Q(\REGISTERS[19][24] ) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n1547), .CK(CLK), .Q(\REGISTERS[19][23] ) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n1546), .CK(CLK), .Q(\REGISTERS[19][22] ) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n1545), .CK(CLK), .Q(\REGISTERS[19][21] ) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n1544), .CK(CLK), .Q(\REGISTERS[19][20] ) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n1543), .CK(CLK), .Q(\REGISTERS[19][19] ) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n1542), .CK(CLK), .Q(\REGISTERS[19][18] ) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n1541), .CK(CLK), .Q(\REGISTERS[19][17] ) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n1540), .CK(CLK), .Q(\REGISTERS[19][16] ) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n1539), .CK(CLK), .Q(\REGISTERS[19][15] ) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n1538), .CK(CLK), .Q(\REGISTERS[19][14] ) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n1537), .CK(CLK), .Q(\REGISTERS[19][13] ) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n1536), .CK(CLK), .Q(\REGISTERS[19][12] ) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n1535), .CK(CLK), .Q(\REGISTERS[19][11] ) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n1534), .CK(CLK), .Q(\REGISTERS[19][10] ) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n1533), .CK(CLK), .Q(\REGISTERS[19][9] )
         );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n1532), .CK(CLK), .Q(\REGISTERS[19][8] )
         );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n1531), .CK(CLK), .Q(\REGISTERS[19][7] )
         );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n1530), .CK(CLK), .Q(\REGISTERS[19][6] )
         );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n1529), .CK(CLK), .Q(\REGISTERS[19][5] )
         );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n1528), .CK(CLK), .Q(\REGISTERS[19][4] )
         );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n1527), .CK(CLK), .Q(\REGISTERS[19][3] )
         );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n1526), .CK(CLK), .Q(\REGISTERS[19][2] )
         );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n1525), .CK(CLK), .Q(\REGISTERS[19][1] )
         );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n1524), .CK(CLK), .Q(\REGISTERS[19][0] )
         );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n1523), .CK(CLK), .Q(\REGISTERS[20][31] ) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n1522), .CK(CLK), .Q(\REGISTERS[20][30] ) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n1521), .CK(CLK), .Q(\REGISTERS[20][29] ) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n1520), .CK(CLK), .Q(\REGISTERS[20][28] ) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n1519), .CK(CLK), .Q(\REGISTERS[20][27] ) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n1518), .CK(CLK), .Q(\REGISTERS[20][26] ) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n1517), .CK(CLK), .Q(\REGISTERS[20][25] ) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n1516), .CK(CLK), .Q(\REGISTERS[20][24] ) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n1515), .CK(CLK), .Q(\REGISTERS[20][23] ) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n1514), .CK(CLK), .Q(\REGISTERS[20][22] ) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n1513), .CK(CLK), .Q(\REGISTERS[20][21] ) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n1512), .CK(CLK), .Q(\REGISTERS[20][20] ) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n1511), .CK(CLK), .Q(\REGISTERS[20][19] ) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n1510), .CK(CLK), .Q(\REGISTERS[20][18] ) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n1509), .CK(CLK), .Q(\REGISTERS[20][17] ) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n1508), .CK(CLK), .Q(\REGISTERS[20][16] ) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n1507), .CK(CLK), .Q(\REGISTERS[20][15] ) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n1506), .CK(CLK), .Q(\REGISTERS[20][14] ) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n1505), .CK(CLK), .Q(\REGISTERS[20][13] ) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n1504), .CK(CLK), .Q(\REGISTERS[20][12] ) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n1503), .CK(CLK), .Q(\REGISTERS[20][11] ) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n1502), .CK(CLK), .Q(\REGISTERS[20][10] ) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n1501), .CK(CLK), .Q(\REGISTERS[20][9] )
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n1500), .CK(CLK), .Q(\REGISTERS[20][8] )
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n1499), .CK(CLK), .Q(\REGISTERS[20][7] )
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n1498), .CK(CLK), .Q(\REGISTERS[20][6] )
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n1497), .CK(CLK), .Q(\REGISTERS[20][5] )
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n1496), .CK(CLK), .Q(\REGISTERS[20][4] )
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n1495), .CK(CLK), .Q(\REGISTERS[20][3] )
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n1494), .CK(CLK), .Q(\REGISTERS[20][2] )
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n1493), .CK(CLK), .Q(\REGISTERS[20][1] )
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n1492), .CK(CLK), .Q(\REGISTERS[20][0] )
         );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n1491), .CK(CLK), .Q(\REGISTERS[21][31] ) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n1490), .CK(CLK), .Q(\REGISTERS[21][30] ) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n1489), .CK(CLK), .Q(\REGISTERS[21][29] ) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n1488), .CK(CLK), .Q(\REGISTERS[21][28] ) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n1487), .CK(CLK), .Q(\REGISTERS[21][27] ) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n1486), .CK(CLK), .Q(\REGISTERS[21][26] ) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n1485), .CK(CLK), .Q(\REGISTERS[21][25] ) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n1484), .CK(CLK), .Q(\REGISTERS[21][24] ) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n1483), .CK(CLK), .Q(\REGISTERS[21][23] ) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n1482), .CK(CLK), .Q(\REGISTERS[21][22] ) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n1481), .CK(CLK), .Q(\REGISTERS[21][21] ) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n1480), .CK(CLK), .Q(\REGISTERS[21][20] ) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n1479), .CK(CLK), .Q(\REGISTERS[21][19] ) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n1478), .CK(CLK), .Q(\REGISTERS[21][18] ) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n1477), .CK(CLK), .Q(\REGISTERS[21][17] ) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n1476), .CK(CLK), .Q(\REGISTERS[21][16] ) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n1475), .CK(CLK), .Q(\REGISTERS[21][15] ) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n1474), .CK(CLK), .Q(\REGISTERS[21][14] ) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n1473), .CK(CLK), .Q(\REGISTERS[21][13] ) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n1472), .CK(CLK), .Q(\REGISTERS[21][12] ) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n1471), .CK(CLK), .Q(\REGISTERS[21][11] ) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n1470), .CK(CLK), .Q(\REGISTERS[21][10] ) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n1469), .CK(CLK), .Q(\REGISTERS[21][9] )
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n1468), .CK(CLK), .Q(\REGISTERS[21][8] )
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n1467), .CK(CLK), .Q(\REGISTERS[21][7] )
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n1466), .CK(CLK), .Q(\REGISTERS[21][6] )
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n1465), .CK(CLK), .Q(\REGISTERS[21][5] )
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n1464), .CK(CLK), .Q(\REGISTERS[21][4] )
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n1463), .CK(CLK), .Q(\REGISTERS[21][3] )
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n1462), .CK(CLK), .Q(\REGISTERS[21][2] )
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n1461), .CK(CLK), .Q(\REGISTERS[21][1] )
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n1460), .CK(CLK), .Q(\REGISTERS[21][0] )
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n1459), .CK(CLK), .Q(\REGISTERS[22][31] ) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n1458), .CK(CLK), .Q(\REGISTERS[22][30] ) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n1457), .CK(CLK), .Q(\REGISTERS[22][29] ) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n1456), .CK(CLK), .Q(\REGISTERS[22][28] ) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n1455), .CK(CLK), .Q(\REGISTERS[22][27] ) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n1454), .CK(CLK), .Q(\REGISTERS[22][26] ) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n1453), .CK(CLK), .Q(\REGISTERS[22][25] ) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n1452), .CK(CLK), .Q(\REGISTERS[22][24] ) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n1451), .CK(CLK), .Q(\REGISTERS[22][23] ) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n1450), .CK(CLK), .Q(\REGISTERS[22][22] ) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n1449), .CK(CLK), .Q(\REGISTERS[22][21] ) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n1448), .CK(CLK), .Q(\REGISTERS[22][20] ) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n1447), .CK(CLK), .Q(\REGISTERS[22][19] ) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n1446), .CK(CLK), .Q(\REGISTERS[22][18] ) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n1445), .CK(CLK), .Q(\REGISTERS[22][17] ) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n1444), .CK(CLK), .Q(\REGISTERS[22][16] ) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n1443), .CK(CLK), .Q(\REGISTERS[22][15] ) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n1442), .CK(CLK), .Q(\REGISTERS[22][14] ) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n1441), .CK(CLK), .Q(\REGISTERS[22][13] ) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n1440), .CK(CLK), .Q(\REGISTERS[22][12] ) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n1439), .CK(CLK), .Q(\REGISTERS[22][11] ) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n1438), .CK(CLK), .Q(\REGISTERS[22][10] ) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n1437), .CK(CLK), .Q(\REGISTERS[22][9] )
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n1436), .CK(CLK), .Q(\REGISTERS[22][8] )
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n1435), .CK(CLK), .Q(\REGISTERS[22][7] )
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n1434), .CK(CLK), .Q(\REGISTERS[22][6] )
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n1433), .CK(CLK), .Q(\REGISTERS[22][5] )
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n1432), .CK(CLK), .Q(\REGISTERS[22][4] )
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n1431), .CK(CLK), .Q(\REGISTERS[22][3] )
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n1430), .CK(CLK), .Q(\REGISTERS[22][2] )
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n1429), .CK(CLK), .Q(\REGISTERS[22][1] )
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n1428), .CK(CLK), .Q(\REGISTERS[22][0] )
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n1427), .CK(CLK), .Q(\REGISTERS[23][31] ) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n1426), .CK(CLK), .Q(\REGISTERS[23][30] ) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n1425), .CK(CLK), .Q(\REGISTERS[23][29] ) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n1424), .CK(CLK), .Q(\REGISTERS[23][28] ) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n1423), .CK(CLK), .Q(\REGISTERS[23][27] ) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n1422), .CK(CLK), .Q(\REGISTERS[23][26] ) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n1421), .CK(CLK), .Q(\REGISTERS[23][25] ) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n1420), .CK(CLK), .Q(\REGISTERS[23][24] ) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n1419), .CK(CLK), .Q(\REGISTERS[23][23] ) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n1418), .CK(CLK), .Q(\REGISTERS[23][22] ) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n1417), .CK(CLK), .Q(\REGISTERS[23][21] ) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n1416), .CK(CLK), .Q(\REGISTERS[23][20] ) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n1415), .CK(CLK), .Q(\REGISTERS[23][19] ) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n1414), .CK(CLK), .Q(\REGISTERS[23][18] ) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n1413), .CK(CLK), .Q(\REGISTERS[23][17] ) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n1412), .CK(CLK), .Q(\REGISTERS[23][16] ) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n1411), .CK(CLK), .Q(\REGISTERS[23][15] ) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n1410), .CK(CLK), .Q(\REGISTERS[23][14] ) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n1409), .CK(CLK), .Q(\REGISTERS[23][13] ) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n1408), .CK(CLK), .Q(\REGISTERS[23][12] ) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n1407), .CK(CLK), .Q(\REGISTERS[23][11] ) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n1406), .CK(CLK), .Q(\REGISTERS[23][10] ) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n1405), .CK(CLK), .Q(\REGISTERS[23][9] )
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n1404), .CK(CLK), .Q(\REGISTERS[23][8] )
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n1403), .CK(CLK), .Q(\REGISTERS[23][7] )
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n1402), .CK(CLK), .Q(\REGISTERS[23][6] )
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n1401), .CK(CLK), .Q(\REGISTERS[23][5] )
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n1400), .CK(CLK), .Q(\REGISTERS[23][4] )
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n1399), .CK(CLK), .Q(\REGISTERS[23][3] )
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n1398), .CK(CLK), .Q(\REGISTERS[23][2] )
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n1397), .CK(CLK), .Q(\REGISTERS[23][1] )
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n1396), .CK(CLK), .Q(\REGISTERS[23][0] )
         );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n1395), .CK(CLK), .Q(\REGISTERS[24][31] ) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n1394), .CK(CLK), .Q(\REGISTERS[24][30] ) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n1393), .CK(CLK), .Q(\REGISTERS[24][29] ) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n1392), .CK(CLK), .Q(\REGISTERS[24][28] ) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n1391), .CK(CLK), .Q(\REGISTERS[24][27] ) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n1390), .CK(CLK), .Q(\REGISTERS[24][26] ) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n1389), .CK(CLK), .Q(\REGISTERS[24][25] ) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n1388), .CK(CLK), .Q(\REGISTERS[24][24] ) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n1387), .CK(CLK), .Q(\REGISTERS[24][23] ) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n1386), .CK(CLK), .Q(\REGISTERS[24][22] ) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n1385), .CK(CLK), .Q(\REGISTERS[24][21] ) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n1384), .CK(CLK), .Q(\REGISTERS[24][20] ) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n1383), .CK(CLK), .Q(\REGISTERS[24][19] ) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n1382), .CK(CLK), .Q(\REGISTERS[24][18] ) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n1381), .CK(CLK), .Q(\REGISTERS[24][17] ) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n1380), .CK(CLK), .Q(\REGISTERS[24][16] ) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n1379), .CK(CLK), .Q(\REGISTERS[24][15] ) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n1378), .CK(CLK), .Q(\REGISTERS[24][14] ) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n1377), .CK(CLK), .Q(\REGISTERS[24][13] ) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n1376), .CK(CLK), .Q(\REGISTERS[24][12] ) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n1375), .CK(CLK), .Q(\REGISTERS[24][11] ) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n1374), .CK(CLK), .Q(\REGISTERS[24][10] ) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n1373), .CK(CLK), .Q(\REGISTERS[24][9] )
         );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n1372), .CK(CLK), .Q(\REGISTERS[24][8] )
         );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n1371), .CK(CLK), .Q(\REGISTERS[24][7] )
         );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n1370), .CK(CLK), .Q(\REGISTERS[24][6] )
         );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n1369), .CK(CLK), .Q(\REGISTERS[24][5] )
         );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n1368), .CK(CLK), .Q(\REGISTERS[24][4] )
         );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n1367), .CK(CLK), .Q(\REGISTERS[24][3] )
         );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n1366), .CK(CLK), .Q(\REGISTERS[24][2] )
         );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n1365), .CK(CLK), .Q(\REGISTERS[24][1] )
         );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n1364), .CK(CLK), .Q(\REGISTERS[24][0] )
         );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n1363), .CK(CLK), .Q(\REGISTERS[25][31] ) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n1362), .CK(CLK), .Q(\REGISTERS[25][30] ) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n1361), .CK(CLK), .Q(\REGISTERS[25][29] ) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n1360), .CK(CLK), .Q(\REGISTERS[25][28] ) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n1359), .CK(CLK), .Q(\REGISTERS[25][27] ) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n1358), .CK(CLK), .Q(\REGISTERS[25][26] ) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n1357), .CK(CLK), .Q(\REGISTERS[25][25] ) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n1356), .CK(CLK), .Q(\REGISTERS[25][24] ) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n1355), .CK(CLK), .Q(\REGISTERS[25][23] ) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n1354), .CK(CLK), .Q(\REGISTERS[25][22] ) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n1353), .CK(CLK), .Q(\REGISTERS[25][21] ) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n1352), .CK(CLK), .Q(\REGISTERS[25][20] ) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n1351), .CK(CLK), .Q(\REGISTERS[25][19] ) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n1350), .CK(CLK), .Q(\REGISTERS[25][18] ) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n1349), .CK(CLK), .Q(\REGISTERS[25][17] ) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n1348), .CK(CLK), .Q(\REGISTERS[25][16] ) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n1347), .CK(CLK), .Q(\REGISTERS[25][15] ) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n1346), .CK(CLK), .Q(\REGISTERS[25][14] ) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n1345), .CK(CLK), .Q(\REGISTERS[25][13] ) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n1344), .CK(CLK), .Q(\REGISTERS[25][12] ) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n1343), .CK(CLK), .Q(\REGISTERS[25][11] ) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n1342), .CK(CLK), .Q(\REGISTERS[25][10] ) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n1341), .CK(CLK), .Q(\REGISTERS[25][9] )
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n1340), .CK(CLK), .Q(\REGISTERS[25][8] )
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n1339), .CK(CLK), .Q(\REGISTERS[25][7] )
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n1338), .CK(CLK), .Q(\REGISTERS[25][6] )
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n1337), .CK(CLK), .Q(\REGISTERS[25][5] )
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n1336), .CK(CLK), .Q(\REGISTERS[25][4] )
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n1335), .CK(CLK), .Q(\REGISTERS[25][3] )
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n1334), .CK(CLK), .Q(\REGISTERS[25][2] )
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n1333), .CK(CLK), .Q(\REGISTERS[25][1] )
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n1332), .CK(CLK), .Q(\REGISTERS[25][0] )
         );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n1331), .CK(CLK), .Q(\REGISTERS[26][31] ) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n1330), .CK(CLK), .Q(\REGISTERS[26][30] ) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n1329), .CK(CLK), .Q(\REGISTERS[26][29] ) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n1328), .CK(CLK), .Q(\REGISTERS[26][28] ) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n1327), .CK(CLK), .Q(\REGISTERS[26][27] ) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n1326), .CK(CLK), .Q(\REGISTERS[26][26] ) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n1325), .CK(CLK), .Q(\REGISTERS[26][25] ) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n1324), .CK(CLK), .Q(\REGISTERS[26][24] ) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n1323), .CK(CLK), .Q(\REGISTERS[26][23] ) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n1322), .CK(CLK), .Q(\REGISTERS[26][22] ) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n1321), .CK(CLK), .Q(\REGISTERS[26][21] ) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n1320), .CK(CLK), .Q(\REGISTERS[26][20] ) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n1319), .CK(CLK), .Q(\REGISTERS[26][19] ) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n1318), .CK(CLK), .Q(\REGISTERS[26][18] ) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n1317), .CK(CLK), .Q(\REGISTERS[26][17] ) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n1316), .CK(CLK), .Q(\REGISTERS[26][16] ) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n1315), .CK(CLK), .Q(\REGISTERS[26][15] ) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n1314), .CK(CLK), .Q(\REGISTERS[26][14] ) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n1313), .CK(CLK), .Q(\REGISTERS[26][13] ) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n1312), .CK(CLK), .Q(\REGISTERS[26][12] ) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n1311), .CK(CLK), .Q(\REGISTERS[26][11] ) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n1310), .CK(CLK), .Q(\REGISTERS[26][10] ) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n1309), .CK(CLK), .Q(\REGISTERS[26][9] )
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n1308), .CK(CLK), .Q(\REGISTERS[26][8] )
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n1307), .CK(CLK), .Q(\REGISTERS[26][7] )
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n1306), .CK(CLK), .Q(\REGISTERS[26][6] )
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n1305), .CK(CLK), .Q(\REGISTERS[26][5] )
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n1304), .CK(CLK), .Q(\REGISTERS[26][4] )
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n1303), .CK(CLK), .Q(\REGISTERS[26][3] )
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n1302), .CK(CLK), .Q(\REGISTERS[26][2] )
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n1301), .CK(CLK), .Q(\REGISTERS[26][1] )
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n1300), .CK(CLK), .Q(\REGISTERS[26][0] )
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n1299), .CK(CLK), .Q(\REGISTERS[27][31] ) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n1298), .CK(CLK), .Q(\REGISTERS[27][30] ) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n1297), .CK(CLK), .Q(\REGISTERS[27][29] ) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n1296), .CK(CLK), .Q(\REGISTERS[27][28] ) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n1295), .CK(CLK), .Q(\REGISTERS[27][27] ) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n1294), .CK(CLK), .Q(\REGISTERS[27][26] ) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n1293), .CK(CLK), .Q(\REGISTERS[27][25] ) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n1292), .CK(CLK), .Q(\REGISTERS[27][24] ) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n1291), .CK(CLK), .Q(\REGISTERS[27][23] ) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n1290), .CK(CLK), .Q(\REGISTERS[27][22] ) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n1289), .CK(CLK), .Q(\REGISTERS[27][21] ) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n1288), .CK(CLK), .Q(\REGISTERS[27][20] ) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n1287), .CK(CLK), .Q(\REGISTERS[27][19] ) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n1286), .CK(CLK), .Q(\REGISTERS[27][18] ) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n1285), .CK(CLK), .Q(\REGISTERS[27][17] ) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n1284), .CK(CLK), .Q(\REGISTERS[27][16] ) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n1283), .CK(CLK), .Q(\REGISTERS[27][15] ) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n1282), .CK(CLK), .Q(\REGISTERS[27][14] ) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n1281), .CK(CLK), .Q(\REGISTERS[27][13] ) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n1280), .CK(CLK), .Q(\REGISTERS[27][12] ) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n1279), .CK(CLK), .Q(\REGISTERS[27][11] ) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n1278), .CK(CLK), .Q(\REGISTERS[27][10] ) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n1277), .CK(CLK), .Q(\REGISTERS[27][9] )
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n1276), .CK(CLK), .Q(\REGISTERS[27][8] )
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n1275), .CK(CLK), .Q(\REGISTERS[27][7] )
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n1274), .CK(CLK), .Q(\REGISTERS[27][6] )
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n1273), .CK(CLK), .Q(\REGISTERS[27][5] )
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n1272), .CK(CLK), .Q(\REGISTERS[27][4] )
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n1271), .CK(CLK), .Q(\REGISTERS[27][3] )
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n1270), .CK(CLK), .Q(\REGISTERS[27][2] )
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n1269), .CK(CLK), .Q(\REGISTERS[27][1] )
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n1268), .CK(CLK), .Q(\REGISTERS[27][0] )
         );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n1267), .CK(CLK), .Q(\REGISTERS[28][31] ) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n1266), .CK(CLK), .Q(\REGISTERS[28][30] ) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n1265), .CK(CLK), .Q(\REGISTERS[28][29] ) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n1264), .CK(CLK), .Q(\REGISTERS[28][28] ) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n1263), .CK(CLK), .Q(\REGISTERS[28][27] ) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n1262), .CK(CLK), .Q(\REGISTERS[28][26] ) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n1261), .CK(CLK), .Q(\REGISTERS[28][25] ) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n1260), .CK(CLK), .Q(\REGISTERS[28][24] ) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n1259), .CK(CLK), .Q(\REGISTERS[28][23] ) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n1258), .CK(CLK), .Q(\REGISTERS[28][22] ) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n1257), .CK(CLK), .Q(\REGISTERS[28][21] ) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n1256), .CK(CLK), .Q(\REGISTERS[28][20] ) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n1255), .CK(CLK), .Q(\REGISTERS[28][19] ) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n1254), .CK(CLK), .Q(\REGISTERS[28][18] ) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n1253), .CK(CLK), .Q(\REGISTERS[28][17] ) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n1252), .CK(CLK), .Q(\REGISTERS[28][16] ) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n1251), .CK(CLK), .Q(\REGISTERS[28][15] ) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n1250), .CK(CLK), .Q(\REGISTERS[28][14] ) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n1249), .CK(CLK), .Q(\REGISTERS[28][13] ) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n1248), .CK(CLK), .Q(\REGISTERS[28][12] ) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n1247), .CK(CLK), .Q(\REGISTERS[28][11] ) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n1246), .CK(CLK), .Q(\REGISTERS[28][10] ) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n1245), .CK(CLK), .Q(\REGISTERS[28][9] )
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n1244), .CK(CLK), .Q(\REGISTERS[28][8] )
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n1243), .CK(CLK), .Q(\REGISTERS[28][7] )
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n1242), .CK(CLK), .Q(\REGISTERS[28][6] )
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n1241), .CK(CLK), .Q(\REGISTERS[28][5] )
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n1240), .CK(CLK), .Q(\REGISTERS[28][4] )
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n1239), .CK(CLK), .Q(\REGISTERS[28][3] )
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n1238), .CK(CLK), .Q(\REGISTERS[28][2] )
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n1237), .CK(CLK), .Q(\REGISTERS[28][1] )
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n1236), .CK(CLK), .Q(\REGISTERS[28][0] )
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n1235), .CK(CLK), .Q(\REGISTERS[29][31] ) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n1234), .CK(CLK), .Q(\REGISTERS[29][30] ) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n1233), .CK(CLK), .Q(\REGISTERS[29][29] ) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n1232), .CK(CLK), .Q(\REGISTERS[29][28] ) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n1231), .CK(CLK), .Q(\REGISTERS[29][27] ) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n1230), .CK(CLK), .Q(\REGISTERS[29][26] ) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n1229), .CK(CLK), .Q(\REGISTERS[29][25] ) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n1228), .CK(CLK), .Q(\REGISTERS[29][24] ) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n1227), .CK(CLK), .Q(\REGISTERS[29][23] ) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n1226), .CK(CLK), .Q(\REGISTERS[29][22] ) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n1225), .CK(CLK), .Q(\REGISTERS[29][21] ) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n1224), .CK(CLK), .Q(\REGISTERS[29][20] ) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n1223), .CK(CLK), .Q(\REGISTERS[29][19] ) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n1222), .CK(CLK), .Q(\REGISTERS[29][18] ) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n1221), .CK(CLK), .Q(\REGISTERS[29][17] ) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n1220), .CK(CLK), .Q(\REGISTERS[29][16] ) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n1219), .CK(CLK), .Q(\REGISTERS[29][15] ) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n1218), .CK(CLK), .Q(\REGISTERS[29][14] ) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n1217), .CK(CLK), .Q(\REGISTERS[29][13] ) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n1216), .CK(CLK), .Q(\REGISTERS[29][12] ) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n1215), .CK(CLK), .Q(\REGISTERS[29][11] ) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n1214), .CK(CLK), .Q(\REGISTERS[29][10] ) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n1213), .CK(CLK), .Q(\REGISTERS[29][9] )
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n1212), .CK(CLK), .Q(\REGISTERS[29][8] )
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n1211), .CK(CLK), .Q(\REGISTERS[29][7] )
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n1210), .CK(CLK), .Q(\REGISTERS[29][6] )
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n1209), .CK(CLK), .Q(\REGISTERS[29][5] )
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n1208), .CK(CLK), .Q(\REGISTERS[29][4] )
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n1207), .CK(CLK), .Q(\REGISTERS[29][3] )
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n1206), .CK(CLK), .Q(\REGISTERS[29][2] )
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n1205), .CK(CLK), .Q(\REGISTERS[29][1] )
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n1204), .CK(CLK), .Q(\REGISTERS[29][0] )
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n1203), .CK(CLK), .Q(\REGISTERS[30][31] ) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n1202), .CK(CLK), .Q(\REGISTERS[30][30] ) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n1201), .CK(CLK), .Q(\REGISTERS[30][29] ) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n1200), .CK(CLK), .Q(\REGISTERS[30][28] ) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n1199), .CK(CLK), .Q(\REGISTERS[30][27] ) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n1198), .CK(CLK), .Q(\REGISTERS[30][26] ) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n1197), .CK(CLK), .Q(\REGISTERS[30][25] ) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n1196), .CK(CLK), .Q(\REGISTERS[30][24] ) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n1195), .CK(CLK), .Q(\REGISTERS[30][23] ) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n1194), .CK(CLK), .Q(\REGISTERS[30][22] ) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n1193), .CK(CLK), .Q(\REGISTERS[30][21] ) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n1192), .CK(CLK), .Q(\REGISTERS[30][20] ) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n1191), .CK(CLK), .Q(\REGISTERS[30][19] ) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n1190), .CK(CLK), .Q(\REGISTERS[30][18] ) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n1189), .CK(CLK), .Q(\REGISTERS[30][17] ) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n1188), .CK(CLK), .Q(\REGISTERS[30][16] ) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n1187), .CK(CLK), .Q(\REGISTERS[30][15] ) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n1186), .CK(CLK), .Q(\REGISTERS[30][14] ) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n1185), .CK(CLK), .Q(\REGISTERS[30][13] ) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n1184), .CK(CLK), .Q(\REGISTERS[30][12] ) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n1183), .CK(CLK), .Q(\REGISTERS[30][11] ) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n1182), .CK(CLK), .Q(\REGISTERS[30][10] ) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n1181), .CK(CLK), .Q(\REGISTERS[30][9] )
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n1180), .CK(CLK), .Q(\REGISTERS[30][8] )
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n1179), .CK(CLK), .Q(\REGISTERS[30][7] )
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n1178), .CK(CLK), .Q(\REGISTERS[30][6] )
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n1177), .CK(CLK), .Q(\REGISTERS[30][5] )
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n1176), .CK(CLK), .Q(\REGISTERS[30][4] )
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n1175), .CK(CLK), .Q(\REGISTERS[30][3] )
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n1174), .CK(CLK), .Q(\REGISTERS[30][2] )
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n1173), .CK(CLK), .Q(\REGISTERS[30][1] )
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n1172), .CK(CLK), .Q(\REGISTERS[30][0] )
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n1171), .CK(CLK), .Q(\REGISTERS[31][31] ) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n1170), .CK(CLK), .Q(\REGISTERS[31][30] ) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n1169), .CK(CLK), .Q(\REGISTERS[31][29] ) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n1168), .CK(CLK), .Q(\REGISTERS[31][28] ) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n1167), .CK(CLK), .Q(\REGISTERS[31][27] ) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n1166), .CK(CLK), .Q(\REGISTERS[31][26] ) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n1165), .CK(CLK), .Q(\REGISTERS[31][25] ) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n1164), .CK(CLK), .Q(\REGISTERS[31][24] ) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n1163), .CK(CLK), .Q(\REGISTERS[31][23] ) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n1162), .CK(CLK), .Q(\REGISTERS[31][22] ) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n1161), .CK(CLK), .Q(\REGISTERS[31][21] ) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n1160), .CK(CLK), .Q(\REGISTERS[31][20] ) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n1159), .CK(CLK), .Q(\REGISTERS[31][19] ) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n1158), .CK(CLK), .Q(\REGISTERS[31][18] ) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n1157), .CK(CLK), .Q(\REGISTERS[31][17] ) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n1156), .CK(CLK), .Q(\REGISTERS[31][16] ) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n1155), .CK(CLK), .Q(\REGISTERS[31][15] ) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n1154), .CK(CLK), .Q(\REGISTERS[31][14] ) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n1153), .CK(CLK), .Q(\REGISTERS[31][13] ) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n1152), .CK(CLK), .Q(\REGISTERS[31][12] ) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n1151), .CK(CLK), .Q(\REGISTERS[31][11] ) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n1150), .CK(CLK), .Q(\REGISTERS[31][10] ) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n1149), .CK(CLK), .Q(\REGISTERS[31][9] )
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n1148), .CK(CLK), .Q(\REGISTERS[31][8] )
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n1147), .CK(CLK), .Q(\REGISTERS[31][7] )
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n1146), .CK(CLK), .Q(\REGISTERS[31][6] )
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n1145), .CK(CLK), .Q(\REGISTERS[31][5] )
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n1144), .CK(CLK), .Q(\REGISTERS[31][4] )
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n1143), .CK(CLK), .Q(\REGISTERS[31][3] )
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n1142), .CK(CLK), .Q(\REGISTERS[31][2] )
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n1141), .CK(CLK), .Q(\REGISTERS[31][1] )
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n1140), .CK(CLK), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT1_reg[31]  ( .G(N444), .D(N410), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N444), .D(N409), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N444), .D(N408), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N444), .D(N407), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N444), .D(N406), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N444), .D(N405), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N444), .D(N404), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N444), .D(N403), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N444), .D(N402), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N444), .D(N401), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N444), .D(N400), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N444), .D(N399), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N444), .D(N398), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N444), .D(N397), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N444), .D(N396), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N444), .D(N395), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N444), .D(N394), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N444), .D(N393), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N444), .D(N392), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N444), .D(N391), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N444), .D(N390), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N444), .D(N389), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N444), .D(N388), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N444), .D(N387), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N444), .D(N386), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N444), .D(N385), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N444), .D(N384), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N444), .D(N383), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N444), .D(N382), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N444), .D(N381), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N444), .D(N380), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N444), .D(N379), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N445), .D(N443), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N445), .D(N442), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N445), .D(N441), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N445), .D(N440), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N445), .D(N439), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N445), .D(N438), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N445), .D(N437), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N445), .D(N436), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N445), .D(N435), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N445), .D(N434), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N445), .D(N433), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N445), .D(N432), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N445), .D(N431), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N445), .D(N430), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N445), .D(N429), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N445), .D(N428), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N445), .D(N427), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N445), .D(N426), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N445), .D(N425), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N445), .D(N424), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N445), .D(N423), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N445), .D(N422), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N445), .D(N421), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N445), .D(N420), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N445), .D(N419), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N445), .D(N418), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N445), .D(N417), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N445), .D(N416), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N445), .D(N415), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N445), .D(N414), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N445), .D(N413), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N445), .D(N412), .Q(OUT2[0]) );
  INV_X1 U3 ( .A(n3083), .ZN(n1) );
  INV_X2 U4 ( .A(n1), .ZN(n2) );
  INV_X1 U5 ( .A(n3084), .ZN(n3) );
  INV_X2 U6 ( .A(n3), .ZN(n4) );
  INV_X1 U7 ( .A(n3085), .ZN(n5) );
  INV_X2 U8 ( .A(n5), .ZN(n6) );
  INV_X1 U9 ( .A(n3086), .ZN(n7) );
  INV_X2 U10 ( .A(n7), .ZN(n8) );
  INV_X1 U11 ( .A(n3087), .ZN(n9) );
  INV_X2 U12 ( .A(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n3088), .ZN(n11) );
  INV_X2 U14 ( .A(n11), .ZN(n12) );
  INV_X1 U15 ( .A(n3089), .ZN(n13) );
  INV_X2 U16 ( .A(n13), .ZN(n14) );
  INV_X1 U17 ( .A(n3077), .ZN(n15) );
  INV_X2 U18 ( .A(n15), .ZN(n16) );
  INV_X1 U19 ( .A(n3078), .ZN(n17) );
  INV_X2 U20 ( .A(n17), .ZN(n18) );
  INV_X1 U21 ( .A(n3075), .ZN(n19) );
  INV_X2 U22 ( .A(n19), .ZN(n20) );
  INV_X1 U23 ( .A(n3076), .ZN(n21) );
  INV_X2 U24 ( .A(n21), .ZN(n22) );
  INV_X1 U25 ( .A(n3073), .ZN(n23) );
  INV_X2 U26 ( .A(n23), .ZN(n24) );
  INV_X1 U27 ( .A(n3074), .ZN(n25) );
  INV_X2 U28 ( .A(n25), .ZN(n26) );
  INV_X1 U29 ( .A(n3071), .ZN(n27) );
  INV_X2 U30 ( .A(n27), .ZN(n28) );
  INV_X1 U31 ( .A(n3072), .ZN(n29) );
  INV_X2 U32 ( .A(n29), .ZN(n30) );
  INV_X1 U33 ( .A(n3068), .ZN(n31) );
  INV_X2 U34 ( .A(n31), .ZN(n32) );
  INV_X1 U35 ( .A(n3069), .ZN(n33) );
  INV_X2 U36 ( .A(n33), .ZN(n34) );
  INV_X1 U37 ( .A(n3066), .ZN(n35) );
  INV_X2 U38 ( .A(n35), .ZN(n36) );
  INV_X1 U39 ( .A(n3067), .ZN(n37) );
  INV_X2 U40 ( .A(n37), .ZN(n38) );
  INV_X1 U41 ( .A(n3064), .ZN(n39) );
  INV_X2 U42 ( .A(n39), .ZN(n40) );
  INV_X1 U43 ( .A(n3065), .ZN(n41) );
  INV_X2 U44 ( .A(n41), .ZN(n42) );
  INV_X1 U45 ( .A(n3062), .ZN(n43) );
  INV_X2 U46 ( .A(n43), .ZN(n44) );
  INV_X1 U47 ( .A(n3063), .ZN(n45) );
  INV_X2 U48 ( .A(n45), .ZN(n46) );
  INV_X1 U49 ( .A(n3055), .ZN(n47) );
  INV_X2 U50 ( .A(n47), .ZN(n48) );
  INV_X1 U51 ( .A(n3060), .ZN(n49) );
  INV_X2 U52 ( .A(n49), .ZN(n50) );
  INV_X1 U53 ( .A(n3051), .ZN(n51) );
  INV_X2 U54 ( .A(n51), .ZN(n52) );
  INV_X1 U55 ( .A(n3053), .ZN(n53) );
  INV_X2 U56 ( .A(n53), .ZN(n54) );
  INV_X1 U57 ( .A(n3047), .ZN(n55) );
  INV_X2 U58 ( .A(n55), .ZN(n56) );
  INV_X1 U59 ( .A(n3049), .ZN(n57) );
  INV_X2 U60 ( .A(n57), .ZN(n58) );
  INV_X1 U61 ( .A(n3043), .ZN(n59) );
  INV_X2 U62 ( .A(n59), .ZN(n60) );
  INV_X1 U63 ( .A(n3045), .ZN(n61) );
  INV_X2 U64 ( .A(n61), .ZN(n62) );
  OAI21_X4 U65 ( .B1(n3040), .B2(n3041), .A(n3042), .ZN(n3008) );
  INV_X4 U66 ( .A(RESET), .ZN(n3042) );
  MUX2_X1 U67 ( .A(\REGISTERS[15][0] ), .B(\REGISTERS[31][0] ), .S(ADD_RD2[4]), 
        .Z(n63) );
  MUX2_X1 U68 ( .A(\REGISTERS[7][0] ), .B(\REGISTERS[23][0] ), .S(ADD_RD2[4]), 
        .Z(n64) );
  MUX2_X1 U69 ( .A(n64), .B(n63), .S(ADD_RD2[3]), .Z(n65) );
  MUX2_X1 U70 ( .A(\REGISTERS[11][0] ), .B(\REGISTERS[27][0] ), .S(ADD_RD2[4]), 
        .Z(n66) );
  MUX2_X1 U71 ( .A(\REGISTERS[3][0] ), .B(\REGISTERS[19][0] ), .S(ADD_RD2[4]), 
        .Z(n67) );
  MUX2_X1 U72 ( .A(n67), .B(n66), .S(ADD_RD2[3]), .Z(n68) );
  MUX2_X1 U73 ( .A(n68), .B(n65), .S(ADD_RD2[2]), .Z(n69) );
  MUX2_X1 U74 ( .A(\REGISTERS[14][0] ), .B(\REGISTERS[30][0] ), .S(ADD_RD2[4]), 
        .Z(n70) );
  MUX2_X1 U75 ( .A(\REGISTERS[6][0] ), .B(\REGISTERS[22][0] ), .S(ADD_RD2[4]), 
        .Z(n71) );
  MUX2_X1 U76 ( .A(n71), .B(n70), .S(ADD_RD2[3]), .Z(n72) );
  MUX2_X1 U77 ( .A(\REGISTERS[10][0] ), .B(\REGISTERS[26][0] ), .S(ADD_RD2[4]), 
        .Z(n73) );
  MUX2_X1 U78 ( .A(\REGISTERS[2][0] ), .B(\REGISTERS[18][0] ), .S(ADD_RD2[4]), 
        .Z(n74) );
  MUX2_X1 U79 ( .A(n74), .B(n73), .S(ADD_RD2[3]), .Z(n75) );
  MUX2_X1 U80 ( .A(n75), .B(n72), .S(ADD_RD2[2]), .Z(n76) );
  MUX2_X1 U81 ( .A(n76), .B(n69), .S(ADD_RD2[0]), .Z(n77) );
  MUX2_X1 U82 ( .A(\REGISTERS[13][0] ), .B(\REGISTERS[29][0] ), .S(ADD_RD2[4]), 
        .Z(n78) );
  MUX2_X1 U83 ( .A(\REGISTERS[5][0] ), .B(\REGISTERS[21][0] ), .S(ADD_RD2[4]), 
        .Z(n79) );
  MUX2_X1 U84 ( .A(n79), .B(n78), .S(ADD_RD2[3]), .Z(n80) );
  MUX2_X1 U85 ( .A(\REGISTERS[9][0] ), .B(\REGISTERS[25][0] ), .S(ADD_RD2[4]), 
        .Z(n81) );
  MUX2_X1 U86 ( .A(\REGISTERS[1][0] ), .B(\REGISTERS[17][0] ), .S(ADD_RD2[4]), 
        .Z(n82) );
  MUX2_X1 U87 ( .A(n82), .B(n81), .S(ADD_RD2[3]), .Z(n83) );
  MUX2_X1 U88 ( .A(n83), .B(n80), .S(ADD_RD2[2]), .Z(n84) );
  MUX2_X1 U89 ( .A(\REGISTERS[12][0] ), .B(\REGISTERS[28][0] ), .S(ADD_RD2[4]), 
        .Z(n85) );
  MUX2_X1 U90 ( .A(\REGISTERS[4][0] ), .B(\REGISTERS[20][0] ), .S(ADD_RD2[4]), 
        .Z(n86) );
  MUX2_X1 U91 ( .A(n86), .B(n85), .S(ADD_RD2[3]), .Z(n87) );
  MUX2_X1 U92 ( .A(\REGISTERS[8][0] ), .B(\REGISTERS[24][0] ), .S(ADD_RD2[4]), 
        .Z(n88) );
  MUX2_X1 U93 ( .A(\REGISTERS[0][0] ), .B(\REGISTERS[16][0] ), .S(ADD_RD2[4]), 
        .Z(n89) );
  MUX2_X1 U94 ( .A(n89), .B(n88), .S(ADD_RD2[3]), .Z(n90) );
  MUX2_X1 U95 ( .A(n90), .B(n87), .S(ADD_RD2[2]), .Z(n91) );
  MUX2_X1 U96 ( .A(n91), .B(n84), .S(ADD_RD2[0]), .Z(n92) );
  MUX2_X1 U97 ( .A(n92), .B(n77), .S(ADD_RD2[1]), .Z(N412) );
  MUX2_X1 U98 ( .A(\REGISTERS[15][1] ), .B(\REGISTERS[31][1] ), .S(ADD_RD2[4]), 
        .Z(n93) );
  MUX2_X1 U99 ( .A(\REGISTERS[7][1] ), .B(\REGISTERS[23][1] ), .S(ADD_RD2[4]), 
        .Z(n94) );
  MUX2_X1 U100 ( .A(n94), .B(n93), .S(ADD_RD2[3]), .Z(n95) );
  MUX2_X1 U101 ( .A(\REGISTERS[11][1] ), .B(\REGISTERS[27][1] ), .S(ADD_RD2[4]), .Z(n96) );
  MUX2_X1 U102 ( .A(\REGISTERS[3][1] ), .B(\REGISTERS[19][1] ), .S(ADD_RD2[4]), 
        .Z(n97) );
  MUX2_X1 U103 ( .A(n97), .B(n96), .S(ADD_RD2[3]), .Z(n98) );
  MUX2_X1 U104 ( .A(n98), .B(n95), .S(ADD_RD2[2]), .Z(n99) );
  MUX2_X1 U105 ( .A(\REGISTERS[14][1] ), .B(\REGISTERS[30][1] ), .S(ADD_RD2[4]), .Z(n100) );
  MUX2_X1 U106 ( .A(\REGISTERS[6][1] ), .B(\REGISTERS[22][1] ), .S(ADD_RD2[4]), 
        .Z(n101) );
  MUX2_X1 U107 ( .A(n101), .B(n100), .S(ADD_RD2[3]), .Z(n102) );
  MUX2_X1 U108 ( .A(\REGISTERS[10][1] ), .B(\REGISTERS[26][1] ), .S(ADD_RD2[4]), .Z(n103) );
  MUX2_X1 U109 ( .A(\REGISTERS[2][1] ), .B(\REGISTERS[18][1] ), .S(ADD_RD2[4]), 
        .Z(n104) );
  MUX2_X1 U110 ( .A(n104), .B(n103), .S(ADD_RD2[3]), .Z(n105) );
  MUX2_X1 U111 ( .A(n105), .B(n102), .S(ADD_RD2[2]), .Z(n106) );
  MUX2_X1 U112 ( .A(n106), .B(n99), .S(ADD_RD2[0]), .Z(n107) );
  MUX2_X1 U113 ( .A(\REGISTERS[13][1] ), .B(\REGISTERS[29][1] ), .S(ADD_RD2[4]), .Z(n108) );
  MUX2_X1 U114 ( .A(\REGISTERS[5][1] ), .B(\REGISTERS[21][1] ), .S(ADD_RD2[4]), 
        .Z(n109) );
  MUX2_X1 U115 ( .A(n109), .B(n108), .S(ADD_RD2[3]), .Z(n110) );
  MUX2_X1 U116 ( .A(\REGISTERS[9][1] ), .B(\REGISTERS[25][1] ), .S(ADD_RD2[4]), 
        .Z(n111) );
  MUX2_X1 U117 ( .A(\REGISTERS[1][1] ), .B(\REGISTERS[17][1] ), .S(ADD_RD2[4]), 
        .Z(n112) );
  MUX2_X1 U118 ( .A(n112), .B(n111), .S(ADD_RD2[3]), .Z(n113) );
  MUX2_X1 U119 ( .A(n113), .B(n110), .S(ADD_RD2[2]), .Z(n114) );
  MUX2_X1 U120 ( .A(\REGISTERS[12][1] ), .B(\REGISTERS[28][1] ), .S(ADD_RD2[4]), .Z(n115) );
  MUX2_X1 U121 ( .A(\REGISTERS[4][1] ), .B(\REGISTERS[20][1] ), .S(ADD_RD2[4]), 
        .Z(n116) );
  MUX2_X1 U122 ( .A(n116), .B(n115), .S(ADD_RD2[3]), .Z(n117) );
  MUX2_X1 U123 ( .A(\REGISTERS[8][1] ), .B(\REGISTERS[24][1] ), .S(ADD_RD2[4]), 
        .Z(n118) );
  MUX2_X1 U124 ( .A(\REGISTERS[0][1] ), .B(\REGISTERS[16][1] ), .S(ADD_RD2[4]), 
        .Z(n119) );
  MUX2_X1 U125 ( .A(n119), .B(n118), .S(ADD_RD2[3]), .Z(n120) );
  MUX2_X1 U126 ( .A(n120), .B(n117), .S(ADD_RD2[2]), .Z(n121) );
  MUX2_X1 U127 ( .A(n121), .B(n114), .S(ADD_RD2[0]), .Z(n122) );
  MUX2_X1 U128 ( .A(n122), .B(n107), .S(ADD_RD2[1]), .Z(N413) );
  MUX2_X1 U129 ( .A(\REGISTERS[15][2] ), .B(\REGISTERS[31][2] ), .S(ADD_RD2[4]), .Z(n123) );
  MUX2_X1 U130 ( .A(\REGISTERS[7][2] ), .B(\REGISTERS[23][2] ), .S(ADD_RD2[4]), 
        .Z(n124) );
  MUX2_X1 U131 ( .A(n124), .B(n123), .S(ADD_RD2[3]), .Z(n125) );
  MUX2_X1 U132 ( .A(\REGISTERS[11][2] ), .B(\REGISTERS[27][2] ), .S(ADD_RD2[4]), .Z(n126) );
  MUX2_X1 U133 ( .A(\REGISTERS[3][2] ), .B(\REGISTERS[19][2] ), .S(ADD_RD2[4]), 
        .Z(n127) );
  MUX2_X1 U134 ( .A(n127), .B(n126), .S(ADD_RD2[3]), .Z(n128) );
  MUX2_X1 U135 ( .A(n128), .B(n125), .S(ADD_RD2[2]), .Z(n129) );
  MUX2_X1 U136 ( .A(\REGISTERS[14][2] ), .B(\REGISTERS[30][2] ), .S(ADD_RD2[4]), .Z(n130) );
  MUX2_X1 U137 ( .A(\REGISTERS[6][2] ), .B(\REGISTERS[22][2] ), .S(ADD_RD2[4]), 
        .Z(n131) );
  MUX2_X1 U138 ( .A(n131), .B(n130), .S(ADD_RD2[3]), .Z(n132) );
  MUX2_X1 U139 ( .A(\REGISTERS[10][2] ), .B(\REGISTERS[26][2] ), .S(ADD_RD2[4]), .Z(n133) );
  MUX2_X1 U140 ( .A(\REGISTERS[2][2] ), .B(\REGISTERS[18][2] ), .S(ADD_RD2[4]), 
        .Z(n134) );
  MUX2_X1 U141 ( .A(n134), .B(n133), .S(ADD_RD2[3]), .Z(n135) );
  MUX2_X1 U142 ( .A(n135), .B(n132), .S(ADD_RD2[2]), .Z(n136) );
  MUX2_X1 U143 ( .A(n136), .B(n129), .S(ADD_RD2[0]), .Z(n137) );
  MUX2_X1 U144 ( .A(\REGISTERS[13][2] ), .B(\REGISTERS[29][2] ), .S(ADD_RD2[4]), .Z(n138) );
  MUX2_X1 U145 ( .A(\REGISTERS[5][2] ), .B(\REGISTERS[21][2] ), .S(ADD_RD2[4]), 
        .Z(n139) );
  MUX2_X1 U146 ( .A(n139), .B(n138), .S(ADD_RD2[3]), .Z(n140) );
  MUX2_X1 U147 ( .A(\REGISTERS[9][2] ), .B(\REGISTERS[25][2] ), .S(ADD_RD2[4]), 
        .Z(n141) );
  MUX2_X1 U148 ( .A(\REGISTERS[1][2] ), .B(\REGISTERS[17][2] ), .S(ADD_RD2[4]), 
        .Z(n142) );
  MUX2_X1 U149 ( .A(n142), .B(n141), .S(ADD_RD2[3]), .Z(n143) );
  MUX2_X1 U150 ( .A(n143), .B(n140), .S(ADD_RD2[2]), .Z(n144) );
  MUX2_X1 U151 ( .A(\REGISTERS[12][2] ), .B(\REGISTERS[28][2] ), .S(ADD_RD2[4]), .Z(n145) );
  MUX2_X1 U152 ( .A(\REGISTERS[4][2] ), .B(\REGISTERS[20][2] ), .S(ADD_RD2[4]), 
        .Z(n146) );
  MUX2_X1 U153 ( .A(n146), .B(n145), .S(ADD_RD2[3]), .Z(n147) );
  MUX2_X1 U154 ( .A(\REGISTERS[8][2] ), .B(\REGISTERS[24][2] ), .S(ADD_RD2[4]), 
        .Z(n148) );
  MUX2_X1 U155 ( .A(\REGISTERS[0][2] ), .B(\REGISTERS[16][2] ), .S(ADD_RD2[4]), 
        .Z(n149) );
  MUX2_X1 U156 ( .A(n149), .B(n148), .S(ADD_RD2[3]), .Z(n150) );
  MUX2_X1 U157 ( .A(n150), .B(n147), .S(ADD_RD2[2]), .Z(n151) );
  MUX2_X1 U158 ( .A(n151), .B(n144), .S(ADD_RD2[0]), .Z(n152) );
  MUX2_X1 U159 ( .A(n152), .B(n137), .S(ADD_RD2[1]), .Z(N414) );
  MUX2_X1 U160 ( .A(\REGISTERS[15][3] ), .B(\REGISTERS[31][3] ), .S(ADD_RD2[4]), .Z(n153) );
  MUX2_X1 U161 ( .A(\REGISTERS[7][3] ), .B(\REGISTERS[23][3] ), .S(ADD_RD2[4]), 
        .Z(n154) );
  MUX2_X1 U162 ( .A(n154), .B(n153), .S(ADD_RD2[3]), .Z(n155) );
  MUX2_X1 U163 ( .A(\REGISTERS[11][3] ), .B(\REGISTERS[27][3] ), .S(ADD_RD2[4]), .Z(n156) );
  MUX2_X1 U164 ( .A(\REGISTERS[3][3] ), .B(\REGISTERS[19][3] ), .S(ADD_RD2[4]), 
        .Z(n157) );
  MUX2_X1 U165 ( .A(n157), .B(n156), .S(ADD_RD2[3]), .Z(n158) );
  MUX2_X1 U166 ( .A(n158), .B(n155), .S(ADD_RD2[2]), .Z(n159) );
  MUX2_X1 U167 ( .A(\REGISTERS[14][3] ), .B(\REGISTERS[30][3] ), .S(ADD_RD2[4]), .Z(n160) );
  MUX2_X1 U168 ( .A(\REGISTERS[6][3] ), .B(\REGISTERS[22][3] ), .S(ADD_RD2[4]), 
        .Z(n161) );
  MUX2_X1 U169 ( .A(n161), .B(n160), .S(ADD_RD2[3]), .Z(n162) );
  MUX2_X1 U170 ( .A(\REGISTERS[10][3] ), .B(\REGISTERS[26][3] ), .S(ADD_RD2[4]), .Z(n163) );
  MUX2_X1 U171 ( .A(\REGISTERS[2][3] ), .B(\REGISTERS[18][3] ), .S(ADD_RD2[4]), 
        .Z(n164) );
  MUX2_X1 U172 ( .A(n164), .B(n163), .S(ADD_RD2[3]), .Z(n165) );
  MUX2_X1 U173 ( .A(n165), .B(n162), .S(ADD_RD2[2]), .Z(n166) );
  MUX2_X1 U174 ( .A(n166), .B(n159), .S(ADD_RD2[0]), .Z(n167) );
  MUX2_X1 U175 ( .A(\REGISTERS[13][3] ), .B(\REGISTERS[29][3] ), .S(ADD_RD2[4]), .Z(n168) );
  MUX2_X1 U176 ( .A(\REGISTERS[5][3] ), .B(\REGISTERS[21][3] ), .S(ADD_RD2[4]), 
        .Z(n169) );
  MUX2_X1 U177 ( .A(n169), .B(n168), .S(ADD_RD2[3]), .Z(n170) );
  MUX2_X1 U178 ( .A(\REGISTERS[9][3] ), .B(\REGISTERS[25][3] ), .S(ADD_RD2[4]), 
        .Z(n171) );
  MUX2_X1 U179 ( .A(\REGISTERS[1][3] ), .B(\REGISTERS[17][3] ), .S(ADD_RD2[4]), 
        .Z(n172) );
  MUX2_X1 U180 ( .A(n172), .B(n171), .S(ADD_RD2[3]), .Z(n173) );
  MUX2_X1 U181 ( .A(n173), .B(n170), .S(ADD_RD2[2]), .Z(n174) );
  MUX2_X1 U182 ( .A(\REGISTERS[12][3] ), .B(\REGISTERS[28][3] ), .S(ADD_RD2[4]), .Z(n175) );
  MUX2_X1 U183 ( .A(\REGISTERS[4][3] ), .B(\REGISTERS[20][3] ), .S(ADD_RD2[4]), 
        .Z(n176) );
  MUX2_X1 U184 ( .A(n176), .B(n175), .S(ADD_RD2[3]), .Z(n177) );
  MUX2_X1 U185 ( .A(\REGISTERS[8][3] ), .B(\REGISTERS[24][3] ), .S(ADD_RD2[4]), 
        .Z(n178) );
  MUX2_X1 U186 ( .A(\REGISTERS[0][3] ), .B(\REGISTERS[16][3] ), .S(ADD_RD2[4]), 
        .Z(n179) );
  MUX2_X1 U187 ( .A(n179), .B(n178), .S(ADD_RD2[3]), .Z(n180) );
  MUX2_X1 U188 ( .A(n180), .B(n177), .S(ADD_RD2[2]), .Z(n181) );
  MUX2_X1 U189 ( .A(n181), .B(n174), .S(ADD_RD2[0]), .Z(n182) );
  MUX2_X1 U190 ( .A(n182), .B(n167), .S(ADD_RD2[1]), .Z(N415) );
  MUX2_X1 U191 ( .A(\REGISTERS[15][4] ), .B(\REGISTERS[31][4] ), .S(ADD_RD2[4]), .Z(n183) );
  MUX2_X1 U192 ( .A(\REGISTERS[7][4] ), .B(\REGISTERS[23][4] ), .S(ADD_RD2[4]), 
        .Z(n184) );
  MUX2_X1 U193 ( .A(n184), .B(n183), .S(ADD_RD2[3]), .Z(n185) );
  MUX2_X1 U194 ( .A(\REGISTERS[11][4] ), .B(\REGISTERS[27][4] ), .S(ADD_RD2[4]), .Z(n186) );
  MUX2_X1 U195 ( .A(\REGISTERS[3][4] ), .B(\REGISTERS[19][4] ), .S(ADD_RD2[4]), 
        .Z(n187) );
  MUX2_X1 U196 ( .A(n187), .B(n186), .S(ADD_RD2[3]), .Z(n188) );
  MUX2_X1 U197 ( .A(n188), .B(n185), .S(ADD_RD2[2]), .Z(n189) );
  MUX2_X1 U198 ( .A(\REGISTERS[14][4] ), .B(\REGISTERS[30][4] ), .S(ADD_RD2[4]), .Z(n190) );
  MUX2_X1 U199 ( .A(\REGISTERS[6][4] ), .B(\REGISTERS[22][4] ), .S(ADD_RD2[4]), 
        .Z(n191) );
  MUX2_X1 U200 ( .A(n191), .B(n190), .S(ADD_RD2[3]), .Z(n192) );
  MUX2_X1 U201 ( .A(\REGISTERS[10][4] ), .B(\REGISTERS[26][4] ), .S(ADD_RD2[4]), .Z(n193) );
  MUX2_X1 U202 ( .A(\REGISTERS[2][4] ), .B(\REGISTERS[18][4] ), .S(ADD_RD2[4]), 
        .Z(n194) );
  MUX2_X1 U203 ( .A(n194), .B(n193), .S(ADD_RD2[3]), .Z(n195) );
  MUX2_X1 U204 ( .A(n195), .B(n192), .S(ADD_RD2[2]), .Z(n196) );
  MUX2_X1 U205 ( .A(n196), .B(n189), .S(ADD_RD2[0]), .Z(n197) );
  MUX2_X1 U206 ( .A(\REGISTERS[13][4] ), .B(\REGISTERS[29][4] ), .S(ADD_RD2[4]), .Z(n198) );
  MUX2_X1 U207 ( .A(\REGISTERS[5][4] ), .B(\REGISTERS[21][4] ), .S(ADD_RD2[4]), 
        .Z(n199) );
  MUX2_X1 U208 ( .A(n199), .B(n198), .S(ADD_RD2[3]), .Z(n200) );
  MUX2_X1 U209 ( .A(\REGISTERS[9][4] ), .B(\REGISTERS[25][4] ), .S(ADD_RD2[4]), 
        .Z(n201) );
  MUX2_X1 U210 ( .A(\REGISTERS[1][4] ), .B(\REGISTERS[17][4] ), .S(ADD_RD2[4]), 
        .Z(n202) );
  MUX2_X1 U211 ( .A(n202), .B(n201), .S(ADD_RD2[3]), .Z(n203) );
  MUX2_X1 U212 ( .A(n203), .B(n200), .S(ADD_RD2[2]), .Z(n204) );
  MUX2_X1 U213 ( .A(\REGISTERS[12][4] ), .B(\REGISTERS[28][4] ), .S(ADD_RD2[4]), .Z(n205) );
  MUX2_X1 U214 ( .A(\REGISTERS[4][4] ), .B(\REGISTERS[20][4] ), .S(ADD_RD2[4]), 
        .Z(n206) );
  MUX2_X1 U215 ( .A(n206), .B(n205), .S(ADD_RD2[3]), .Z(n207) );
  MUX2_X1 U216 ( .A(\REGISTERS[8][4] ), .B(\REGISTERS[24][4] ), .S(ADD_RD2[4]), 
        .Z(n208) );
  MUX2_X1 U217 ( .A(\REGISTERS[0][4] ), .B(\REGISTERS[16][4] ), .S(ADD_RD2[4]), 
        .Z(n209) );
  MUX2_X1 U218 ( .A(n209), .B(n208), .S(ADD_RD2[3]), .Z(n210) );
  MUX2_X1 U219 ( .A(n210), .B(n207), .S(ADD_RD2[2]), .Z(n211) );
  MUX2_X1 U220 ( .A(n211), .B(n204), .S(ADD_RD2[0]), .Z(n212) );
  MUX2_X1 U221 ( .A(n212), .B(n197), .S(ADD_RD2[1]), .Z(N416) );
  MUX2_X1 U222 ( .A(\REGISTERS[15][5] ), .B(\REGISTERS[31][5] ), .S(ADD_RD2[4]), .Z(n213) );
  MUX2_X1 U223 ( .A(\REGISTERS[7][5] ), .B(\REGISTERS[23][5] ), .S(ADD_RD2[4]), 
        .Z(n214) );
  MUX2_X1 U224 ( .A(n214), .B(n213), .S(ADD_RD2[3]), .Z(n215) );
  MUX2_X1 U225 ( .A(\REGISTERS[11][5] ), .B(\REGISTERS[27][5] ), .S(ADD_RD2[4]), .Z(n216) );
  MUX2_X1 U226 ( .A(\REGISTERS[3][5] ), .B(\REGISTERS[19][5] ), .S(ADD_RD2[4]), 
        .Z(n217) );
  MUX2_X1 U227 ( .A(n217), .B(n216), .S(ADD_RD2[3]), .Z(n218) );
  MUX2_X1 U228 ( .A(n218), .B(n215), .S(ADD_RD2[2]), .Z(n219) );
  MUX2_X1 U229 ( .A(\REGISTERS[14][5] ), .B(\REGISTERS[30][5] ), .S(ADD_RD2[4]), .Z(n220) );
  MUX2_X1 U230 ( .A(\REGISTERS[6][5] ), .B(\REGISTERS[22][5] ), .S(ADD_RD2[4]), 
        .Z(n221) );
  MUX2_X1 U231 ( .A(n221), .B(n220), .S(ADD_RD2[3]), .Z(n222) );
  MUX2_X1 U232 ( .A(\REGISTERS[10][5] ), .B(\REGISTERS[26][5] ), .S(ADD_RD2[4]), .Z(n223) );
  MUX2_X1 U233 ( .A(\REGISTERS[2][5] ), .B(\REGISTERS[18][5] ), .S(ADD_RD2[4]), 
        .Z(n224) );
  MUX2_X1 U234 ( .A(n224), .B(n223), .S(ADD_RD2[3]), .Z(n225) );
  MUX2_X1 U235 ( .A(n225), .B(n222), .S(ADD_RD2[2]), .Z(n226) );
  MUX2_X1 U236 ( .A(n226), .B(n219), .S(ADD_RD2[0]), .Z(n227) );
  MUX2_X1 U237 ( .A(\REGISTERS[13][5] ), .B(\REGISTERS[29][5] ), .S(ADD_RD2[4]), .Z(n228) );
  MUX2_X1 U238 ( .A(\REGISTERS[5][5] ), .B(\REGISTERS[21][5] ), .S(ADD_RD2[4]), 
        .Z(n229) );
  MUX2_X1 U239 ( .A(n229), .B(n228), .S(ADD_RD2[3]), .Z(n230) );
  MUX2_X1 U240 ( .A(\REGISTERS[9][5] ), .B(\REGISTERS[25][5] ), .S(ADD_RD2[4]), 
        .Z(n231) );
  MUX2_X1 U241 ( .A(\REGISTERS[1][5] ), .B(\REGISTERS[17][5] ), .S(ADD_RD2[4]), 
        .Z(n232) );
  MUX2_X1 U242 ( .A(n232), .B(n231), .S(ADD_RD2[3]), .Z(n233) );
  MUX2_X1 U243 ( .A(n233), .B(n230), .S(ADD_RD2[2]), .Z(n234) );
  MUX2_X1 U244 ( .A(\REGISTERS[12][5] ), .B(\REGISTERS[28][5] ), .S(ADD_RD2[4]), .Z(n235) );
  MUX2_X1 U245 ( .A(\REGISTERS[4][5] ), .B(\REGISTERS[20][5] ), .S(ADD_RD2[4]), 
        .Z(n236) );
  MUX2_X1 U246 ( .A(n236), .B(n235), .S(ADD_RD2[3]), .Z(n237) );
  MUX2_X1 U247 ( .A(\REGISTERS[8][5] ), .B(\REGISTERS[24][5] ), .S(ADD_RD2[4]), 
        .Z(n238) );
  MUX2_X1 U248 ( .A(\REGISTERS[0][5] ), .B(\REGISTERS[16][5] ), .S(ADD_RD2[4]), 
        .Z(n239) );
  MUX2_X1 U249 ( .A(n239), .B(n238), .S(ADD_RD2[3]), .Z(n240) );
  MUX2_X1 U250 ( .A(n240), .B(n237), .S(ADD_RD2[2]), .Z(n241) );
  MUX2_X1 U251 ( .A(n241), .B(n234), .S(ADD_RD2[0]), .Z(n242) );
  MUX2_X1 U252 ( .A(n242), .B(n227), .S(ADD_RD2[1]), .Z(N417) );
  MUX2_X1 U253 ( .A(\REGISTERS[15][6] ), .B(\REGISTERS[31][6] ), .S(ADD_RD2[4]), .Z(n243) );
  MUX2_X1 U254 ( .A(\REGISTERS[7][6] ), .B(\REGISTERS[23][6] ), .S(ADD_RD2[4]), 
        .Z(n244) );
  MUX2_X1 U255 ( .A(n244), .B(n243), .S(ADD_RD2[3]), .Z(n245) );
  MUX2_X1 U256 ( .A(\REGISTERS[11][6] ), .B(\REGISTERS[27][6] ), .S(ADD_RD2[4]), .Z(n246) );
  MUX2_X1 U257 ( .A(\REGISTERS[3][6] ), .B(\REGISTERS[19][6] ), .S(ADD_RD2[4]), 
        .Z(n247) );
  MUX2_X1 U258 ( .A(n247), .B(n246), .S(ADD_RD2[3]), .Z(n248) );
  MUX2_X1 U259 ( .A(n248), .B(n245), .S(ADD_RD2[2]), .Z(n249) );
  MUX2_X1 U260 ( .A(\REGISTERS[14][6] ), .B(\REGISTERS[30][6] ), .S(ADD_RD2[4]), .Z(n250) );
  MUX2_X1 U261 ( .A(\REGISTERS[6][6] ), .B(\REGISTERS[22][6] ), .S(ADD_RD2[4]), 
        .Z(n251) );
  MUX2_X1 U262 ( .A(n251), .B(n250), .S(ADD_RD2[3]), .Z(n252) );
  MUX2_X1 U263 ( .A(\REGISTERS[10][6] ), .B(\REGISTERS[26][6] ), .S(ADD_RD2[4]), .Z(n253) );
  MUX2_X1 U264 ( .A(\REGISTERS[2][6] ), .B(\REGISTERS[18][6] ), .S(ADD_RD2[4]), 
        .Z(n254) );
  MUX2_X1 U265 ( .A(n254), .B(n253), .S(ADD_RD2[3]), .Z(n255) );
  MUX2_X1 U266 ( .A(n255), .B(n252), .S(ADD_RD2[2]), .Z(n256) );
  MUX2_X1 U267 ( .A(n256), .B(n249), .S(ADD_RD2[0]), .Z(n257) );
  MUX2_X1 U268 ( .A(\REGISTERS[13][6] ), .B(\REGISTERS[29][6] ), .S(ADD_RD2[4]), .Z(n258) );
  MUX2_X1 U269 ( .A(\REGISTERS[5][6] ), .B(\REGISTERS[21][6] ), .S(ADD_RD2[4]), 
        .Z(n259) );
  MUX2_X1 U270 ( .A(n259), .B(n258), .S(ADD_RD2[3]), .Z(n260) );
  MUX2_X1 U271 ( .A(\REGISTERS[9][6] ), .B(\REGISTERS[25][6] ), .S(ADD_RD2[4]), 
        .Z(n261) );
  MUX2_X1 U272 ( .A(\REGISTERS[1][6] ), .B(\REGISTERS[17][6] ), .S(ADD_RD2[4]), 
        .Z(n262) );
  MUX2_X1 U273 ( .A(n262), .B(n261), .S(ADD_RD2[3]), .Z(n263) );
  MUX2_X1 U274 ( .A(n263), .B(n260), .S(ADD_RD2[2]), .Z(n264) );
  MUX2_X1 U275 ( .A(\REGISTERS[12][6] ), .B(\REGISTERS[28][6] ), .S(ADD_RD2[4]), .Z(n265) );
  MUX2_X1 U276 ( .A(\REGISTERS[4][6] ), .B(\REGISTERS[20][6] ), .S(ADD_RD2[4]), 
        .Z(n266) );
  MUX2_X1 U277 ( .A(n266), .B(n265), .S(ADD_RD2[3]), .Z(n267) );
  MUX2_X1 U278 ( .A(\REGISTERS[8][6] ), .B(\REGISTERS[24][6] ), .S(ADD_RD2[4]), 
        .Z(n268) );
  MUX2_X1 U279 ( .A(\REGISTERS[0][6] ), .B(\REGISTERS[16][6] ), .S(ADD_RD2[4]), 
        .Z(n269) );
  MUX2_X1 U280 ( .A(n269), .B(n268), .S(ADD_RD2[3]), .Z(n270) );
  MUX2_X1 U281 ( .A(n270), .B(n267), .S(ADD_RD2[2]), .Z(n271) );
  MUX2_X1 U282 ( .A(n271), .B(n264), .S(ADD_RD2[0]), .Z(n272) );
  MUX2_X1 U283 ( .A(n272), .B(n257), .S(ADD_RD2[1]), .Z(N418) );
  MUX2_X1 U284 ( .A(\REGISTERS[15][7] ), .B(\REGISTERS[31][7] ), .S(ADD_RD2[4]), .Z(n273) );
  MUX2_X1 U285 ( .A(\REGISTERS[7][7] ), .B(\REGISTERS[23][7] ), .S(ADD_RD2[4]), 
        .Z(n274) );
  MUX2_X1 U286 ( .A(n274), .B(n273), .S(ADD_RD2[3]), .Z(n275) );
  MUX2_X1 U287 ( .A(\REGISTERS[11][7] ), .B(\REGISTERS[27][7] ), .S(ADD_RD2[4]), .Z(n276) );
  MUX2_X1 U288 ( .A(\REGISTERS[3][7] ), .B(\REGISTERS[19][7] ), .S(ADD_RD2[4]), 
        .Z(n277) );
  MUX2_X1 U289 ( .A(n277), .B(n276), .S(ADD_RD2[3]), .Z(n278) );
  MUX2_X1 U290 ( .A(n278), .B(n275), .S(ADD_RD2[2]), .Z(n279) );
  MUX2_X1 U291 ( .A(\REGISTERS[14][7] ), .B(\REGISTERS[30][7] ), .S(ADD_RD2[4]), .Z(n280) );
  MUX2_X1 U292 ( .A(\REGISTERS[6][7] ), .B(\REGISTERS[22][7] ), .S(ADD_RD2[4]), 
        .Z(n281) );
  MUX2_X1 U293 ( .A(n281), .B(n280), .S(ADD_RD2[3]), .Z(n282) );
  MUX2_X1 U294 ( .A(\REGISTERS[10][7] ), .B(\REGISTERS[26][7] ), .S(ADD_RD2[4]), .Z(n283) );
  MUX2_X1 U295 ( .A(\REGISTERS[2][7] ), .B(\REGISTERS[18][7] ), .S(ADD_RD2[4]), 
        .Z(n284) );
  MUX2_X1 U296 ( .A(n284), .B(n283), .S(ADD_RD2[3]), .Z(n285) );
  MUX2_X1 U297 ( .A(n285), .B(n282), .S(ADD_RD2[2]), .Z(n286) );
  MUX2_X1 U298 ( .A(n286), .B(n279), .S(ADD_RD2[0]), .Z(n287) );
  MUX2_X1 U299 ( .A(\REGISTERS[13][7] ), .B(\REGISTERS[29][7] ), .S(ADD_RD2[4]), .Z(n288) );
  MUX2_X1 U300 ( .A(\REGISTERS[5][7] ), .B(\REGISTERS[21][7] ), .S(ADD_RD2[4]), 
        .Z(n289) );
  MUX2_X1 U301 ( .A(n289), .B(n288), .S(ADD_RD2[3]), .Z(n290) );
  MUX2_X1 U302 ( .A(\REGISTERS[9][7] ), .B(\REGISTERS[25][7] ), .S(ADD_RD2[4]), 
        .Z(n291) );
  MUX2_X1 U303 ( .A(\REGISTERS[1][7] ), .B(\REGISTERS[17][7] ), .S(ADD_RD2[4]), 
        .Z(n292) );
  MUX2_X1 U304 ( .A(n292), .B(n291), .S(ADD_RD2[3]), .Z(n293) );
  MUX2_X1 U305 ( .A(n293), .B(n290), .S(ADD_RD2[2]), .Z(n294) );
  MUX2_X1 U306 ( .A(\REGISTERS[12][7] ), .B(\REGISTERS[28][7] ), .S(ADD_RD2[4]), .Z(n295) );
  MUX2_X1 U307 ( .A(\REGISTERS[4][7] ), .B(\REGISTERS[20][7] ), .S(ADD_RD2[4]), 
        .Z(n296) );
  MUX2_X1 U308 ( .A(n296), .B(n295), .S(ADD_RD2[3]), .Z(n297) );
  MUX2_X1 U309 ( .A(\REGISTERS[8][7] ), .B(\REGISTERS[24][7] ), .S(ADD_RD2[4]), 
        .Z(n298) );
  MUX2_X1 U310 ( .A(\REGISTERS[0][7] ), .B(\REGISTERS[16][7] ), .S(ADD_RD2[4]), 
        .Z(n299) );
  MUX2_X1 U311 ( .A(n299), .B(n298), .S(ADD_RD2[3]), .Z(n300) );
  MUX2_X1 U312 ( .A(n300), .B(n297), .S(ADD_RD2[2]), .Z(n301) );
  MUX2_X1 U313 ( .A(n301), .B(n294), .S(ADD_RD2[0]), .Z(n302) );
  MUX2_X1 U314 ( .A(n302), .B(n287), .S(ADD_RD2[1]), .Z(N419) );
  MUX2_X1 U315 ( .A(\REGISTERS[15][8] ), .B(\REGISTERS[31][8] ), .S(ADD_RD2[4]), .Z(n303) );
  MUX2_X1 U316 ( .A(\REGISTERS[7][8] ), .B(\REGISTERS[23][8] ), .S(ADD_RD2[4]), 
        .Z(n304) );
  MUX2_X1 U317 ( .A(n304), .B(n303), .S(ADD_RD2[3]), .Z(n305) );
  MUX2_X1 U318 ( .A(\REGISTERS[11][8] ), .B(\REGISTERS[27][8] ), .S(ADD_RD2[4]), .Z(n306) );
  MUX2_X1 U319 ( .A(\REGISTERS[3][8] ), .B(\REGISTERS[19][8] ), .S(ADD_RD2[4]), 
        .Z(n307) );
  MUX2_X1 U320 ( .A(n307), .B(n306), .S(ADD_RD2[3]), .Z(n308) );
  MUX2_X1 U321 ( .A(n308), .B(n305), .S(ADD_RD2[2]), .Z(n309) );
  MUX2_X1 U322 ( .A(\REGISTERS[14][8] ), .B(\REGISTERS[30][8] ), .S(ADD_RD2[4]), .Z(n310) );
  MUX2_X1 U323 ( .A(\REGISTERS[6][8] ), .B(\REGISTERS[22][8] ), .S(ADD_RD2[4]), 
        .Z(n311) );
  MUX2_X1 U324 ( .A(n311), .B(n310), .S(ADD_RD2[3]), .Z(n312) );
  MUX2_X1 U325 ( .A(\REGISTERS[10][8] ), .B(\REGISTERS[26][8] ), .S(ADD_RD2[4]), .Z(n313) );
  MUX2_X1 U326 ( .A(\REGISTERS[2][8] ), .B(\REGISTERS[18][8] ), .S(ADD_RD2[4]), 
        .Z(n314) );
  MUX2_X1 U327 ( .A(n314), .B(n313), .S(ADD_RD2[3]), .Z(n315) );
  MUX2_X1 U328 ( .A(n315), .B(n312), .S(ADD_RD2[2]), .Z(n316) );
  MUX2_X1 U329 ( .A(n316), .B(n309), .S(ADD_RD2[0]), .Z(n317) );
  MUX2_X1 U330 ( .A(\REGISTERS[13][8] ), .B(\REGISTERS[29][8] ), .S(ADD_RD2[4]), .Z(n318) );
  MUX2_X1 U331 ( .A(\REGISTERS[5][8] ), .B(\REGISTERS[21][8] ), .S(ADD_RD2[4]), 
        .Z(n319) );
  MUX2_X1 U332 ( .A(n319), .B(n318), .S(ADD_RD2[3]), .Z(n320) );
  MUX2_X1 U333 ( .A(\REGISTERS[9][8] ), .B(\REGISTERS[25][8] ), .S(ADD_RD2[4]), 
        .Z(n321) );
  MUX2_X1 U334 ( .A(\REGISTERS[1][8] ), .B(\REGISTERS[17][8] ), .S(ADD_RD2[4]), 
        .Z(n322) );
  MUX2_X1 U335 ( .A(n322), .B(n321), .S(ADD_RD2[3]), .Z(n323) );
  MUX2_X1 U336 ( .A(n323), .B(n320), .S(ADD_RD2[2]), .Z(n324) );
  MUX2_X1 U337 ( .A(\REGISTERS[12][8] ), .B(\REGISTERS[28][8] ), .S(ADD_RD2[4]), .Z(n325) );
  MUX2_X1 U338 ( .A(\REGISTERS[4][8] ), .B(\REGISTERS[20][8] ), .S(ADD_RD2[4]), 
        .Z(n326) );
  MUX2_X1 U339 ( .A(n326), .B(n325), .S(ADD_RD2[3]), .Z(n327) );
  MUX2_X1 U340 ( .A(\REGISTERS[8][8] ), .B(\REGISTERS[24][8] ), .S(ADD_RD2[4]), 
        .Z(n328) );
  MUX2_X1 U341 ( .A(\REGISTERS[0][8] ), .B(\REGISTERS[16][8] ), .S(ADD_RD2[4]), 
        .Z(n329) );
  MUX2_X1 U342 ( .A(n329), .B(n328), .S(ADD_RD2[3]), .Z(n330) );
  MUX2_X1 U343 ( .A(n330), .B(n327), .S(ADD_RD2[2]), .Z(n331) );
  MUX2_X1 U344 ( .A(n331), .B(n324), .S(ADD_RD2[0]), .Z(n332) );
  MUX2_X1 U345 ( .A(n332), .B(n317), .S(ADD_RD2[1]), .Z(N420) );
  MUX2_X1 U346 ( .A(\REGISTERS[15][9] ), .B(\REGISTERS[31][9] ), .S(ADD_RD2[4]), .Z(n333) );
  MUX2_X1 U347 ( .A(\REGISTERS[7][9] ), .B(\REGISTERS[23][9] ), .S(ADD_RD2[4]), 
        .Z(n334) );
  MUX2_X1 U348 ( .A(n334), .B(n333), .S(ADD_RD2[3]), .Z(n335) );
  MUX2_X1 U349 ( .A(\REGISTERS[11][9] ), .B(\REGISTERS[27][9] ), .S(ADD_RD2[4]), .Z(n336) );
  MUX2_X1 U350 ( .A(\REGISTERS[3][9] ), .B(\REGISTERS[19][9] ), .S(ADD_RD2[4]), 
        .Z(n337) );
  MUX2_X1 U351 ( .A(n337), .B(n336), .S(ADD_RD2[3]), .Z(n338) );
  MUX2_X1 U352 ( .A(n338), .B(n335), .S(ADD_RD2[2]), .Z(n339) );
  MUX2_X1 U353 ( .A(\REGISTERS[14][9] ), .B(\REGISTERS[30][9] ), .S(ADD_RD2[4]), .Z(n340) );
  MUX2_X1 U354 ( .A(\REGISTERS[6][9] ), .B(\REGISTERS[22][9] ), .S(ADD_RD2[4]), 
        .Z(n341) );
  MUX2_X1 U355 ( .A(n341), .B(n340), .S(ADD_RD2[3]), .Z(n342) );
  MUX2_X1 U356 ( .A(\REGISTERS[10][9] ), .B(\REGISTERS[26][9] ), .S(ADD_RD2[4]), .Z(n343) );
  MUX2_X1 U357 ( .A(\REGISTERS[2][9] ), .B(\REGISTERS[18][9] ), .S(ADD_RD2[4]), 
        .Z(n344) );
  MUX2_X1 U358 ( .A(n344), .B(n343), .S(ADD_RD2[3]), .Z(n345) );
  MUX2_X1 U359 ( .A(n345), .B(n342), .S(ADD_RD2[2]), .Z(n346) );
  MUX2_X1 U360 ( .A(n346), .B(n339), .S(ADD_RD2[0]), .Z(n347) );
  MUX2_X1 U361 ( .A(\REGISTERS[13][9] ), .B(\REGISTERS[29][9] ), .S(ADD_RD2[4]), .Z(n348) );
  MUX2_X1 U362 ( .A(\REGISTERS[5][9] ), .B(\REGISTERS[21][9] ), .S(ADD_RD2[4]), 
        .Z(n349) );
  MUX2_X1 U363 ( .A(n349), .B(n348), .S(ADD_RD2[3]), .Z(n350) );
  MUX2_X1 U364 ( .A(\REGISTERS[9][9] ), .B(\REGISTERS[25][9] ), .S(ADD_RD2[4]), 
        .Z(n351) );
  MUX2_X1 U365 ( .A(\REGISTERS[1][9] ), .B(\REGISTERS[17][9] ), .S(ADD_RD2[4]), 
        .Z(n352) );
  MUX2_X1 U366 ( .A(n352), .B(n351), .S(ADD_RD2[3]), .Z(n353) );
  MUX2_X1 U367 ( .A(n353), .B(n350), .S(ADD_RD2[2]), .Z(n354) );
  MUX2_X1 U368 ( .A(\REGISTERS[12][9] ), .B(\REGISTERS[28][9] ), .S(ADD_RD2[4]), .Z(n355) );
  MUX2_X1 U369 ( .A(\REGISTERS[4][9] ), .B(\REGISTERS[20][9] ), .S(ADD_RD2[4]), 
        .Z(n356) );
  MUX2_X1 U370 ( .A(n356), .B(n355), .S(ADD_RD2[3]), .Z(n357) );
  MUX2_X1 U371 ( .A(\REGISTERS[8][9] ), .B(\REGISTERS[24][9] ), .S(ADD_RD2[4]), 
        .Z(n358) );
  MUX2_X1 U372 ( .A(\REGISTERS[0][9] ), .B(\REGISTERS[16][9] ), .S(ADD_RD2[4]), 
        .Z(n359) );
  MUX2_X1 U373 ( .A(n359), .B(n358), .S(ADD_RD2[3]), .Z(n360) );
  MUX2_X1 U374 ( .A(n360), .B(n357), .S(ADD_RD2[2]), .Z(n361) );
  MUX2_X1 U375 ( .A(n361), .B(n354), .S(ADD_RD2[0]), .Z(n362) );
  MUX2_X1 U376 ( .A(n362), .B(n347), .S(ADD_RD2[1]), .Z(N421) );
  MUX2_X1 U377 ( .A(\REGISTERS[15][10] ), .B(\REGISTERS[31][10] ), .S(
        ADD_RD2[4]), .Z(n363) );
  MUX2_X1 U378 ( .A(\REGISTERS[7][10] ), .B(\REGISTERS[23][10] ), .S(
        ADD_RD2[4]), .Z(n364) );
  MUX2_X1 U379 ( .A(n364), .B(n363), .S(ADD_RD2[3]), .Z(n365) );
  MUX2_X1 U380 ( .A(\REGISTERS[11][10] ), .B(\REGISTERS[27][10] ), .S(
        ADD_RD2[4]), .Z(n366) );
  MUX2_X1 U381 ( .A(\REGISTERS[3][10] ), .B(\REGISTERS[19][10] ), .S(
        ADD_RD2[4]), .Z(n367) );
  MUX2_X1 U382 ( .A(n367), .B(n366), .S(ADD_RD2[3]), .Z(n368) );
  MUX2_X1 U383 ( .A(n368), .B(n365), .S(ADD_RD2[2]), .Z(n369) );
  MUX2_X1 U384 ( .A(\REGISTERS[14][10] ), .B(\REGISTERS[30][10] ), .S(
        ADD_RD2[4]), .Z(n370) );
  MUX2_X1 U385 ( .A(\REGISTERS[6][10] ), .B(\REGISTERS[22][10] ), .S(
        ADD_RD2[4]), .Z(n371) );
  MUX2_X1 U386 ( .A(n371), .B(n370), .S(ADD_RD2[3]), .Z(n372) );
  MUX2_X1 U387 ( .A(\REGISTERS[10][10] ), .B(\REGISTERS[26][10] ), .S(
        ADD_RD2[4]), .Z(n373) );
  MUX2_X1 U388 ( .A(\REGISTERS[2][10] ), .B(\REGISTERS[18][10] ), .S(
        ADD_RD2[4]), .Z(n374) );
  MUX2_X1 U389 ( .A(n374), .B(n373), .S(ADD_RD2[3]), .Z(n375) );
  MUX2_X1 U390 ( .A(n375), .B(n372), .S(ADD_RD2[2]), .Z(n376) );
  MUX2_X1 U391 ( .A(n376), .B(n369), .S(ADD_RD2[0]), .Z(n377) );
  MUX2_X1 U392 ( .A(\REGISTERS[13][10] ), .B(\REGISTERS[29][10] ), .S(
        ADD_RD2[4]), .Z(n378) );
  MUX2_X1 U393 ( .A(\REGISTERS[5][10] ), .B(\REGISTERS[21][10] ), .S(
        ADD_RD2[4]), .Z(n379) );
  MUX2_X1 U394 ( .A(n379), .B(n378), .S(ADD_RD2[3]), .Z(n380) );
  MUX2_X1 U395 ( .A(\REGISTERS[9][10] ), .B(\REGISTERS[25][10] ), .S(
        ADD_RD2[4]), .Z(n381) );
  MUX2_X1 U396 ( .A(\REGISTERS[1][10] ), .B(\REGISTERS[17][10] ), .S(
        ADD_RD2[4]), .Z(n382) );
  MUX2_X1 U397 ( .A(n382), .B(n381), .S(ADD_RD2[3]), .Z(n383) );
  MUX2_X1 U398 ( .A(n383), .B(n380), .S(ADD_RD2[2]), .Z(n384) );
  MUX2_X1 U399 ( .A(\REGISTERS[12][10] ), .B(\REGISTERS[28][10] ), .S(
        ADD_RD2[4]), .Z(n385) );
  MUX2_X1 U400 ( .A(\REGISTERS[4][10] ), .B(\REGISTERS[20][10] ), .S(
        ADD_RD2[4]), .Z(n386) );
  MUX2_X1 U401 ( .A(n386), .B(n385), .S(ADD_RD2[3]), .Z(n387) );
  MUX2_X1 U402 ( .A(\REGISTERS[8][10] ), .B(\REGISTERS[24][10] ), .S(
        ADD_RD2[4]), .Z(n388) );
  MUX2_X1 U403 ( .A(\REGISTERS[0][10] ), .B(\REGISTERS[16][10] ), .S(
        ADD_RD2[4]), .Z(n389) );
  MUX2_X1 U404 ( .A(n389), .B(n388), .S(ADD_RD2[3]), .Z(n390) );
  MUX2_X1 U405 ( .A(n390), .B(n387), .S(ADD_RD2[2]), .Z(n391) );
  MUX2_X1 U406 ( .A(n391), .B(n384), .S(ADD_RD2[0]), .Z(n392) );
  MUX2_X1 U407 ( .A(n392), .B(n377), .S(ADD_RD2[1]), .Z(N422) );
  MUX2_X1 U408 ( .A(\REGISTERS[15][11] ), .B(\REGISTERS[31][11] ), .S(
        ADD_RD2[4]), .Z(n393) );
  MUX2_X1 U409 ( .A(\REGISTERS[7][11] ), .B(\REGISTERS[23][11] ), .S(
        ADD_RD2[4]), .Z(n394) );
  MUX2_X1 U410 ( .A(n394), .B(n393), .S(ADD_RD2[3]), .Z(n395) );
  MUX2_X1 U411 ( .A(\REGISTERS[11][11] ), .B(\REGISTERS[27][11] ), .S(
        ADD_RD2[4]), .Z(n396) );
  MUX2_X1 U412 ( .A(\REGISTERS[3][11] ), .B(\REGISTERS[19][11] ), .S(
        ADD_RD2[4]), .Z(n397) );
  MUX2_X1 U413 ( .A(n397), .B(n396), .S(ADD_RD2[3]), .Z(n398) );
  MUX2_X1 U414 ( .A(n398), .B(n395), .S(ADD_RD2[2]), .Z(n399) );
  MUX2_X1 U415 ( .A(\REGISTERS[14][11] ), .B(\REGISTERS[30][11] ), .S(
        ADD_RD2[4]), .Z(n400) );
  MUX2_X1 U416 ( .A(\REGISTERS[6][11] ), .B(\REGISTERS[22][11] ), .S(
        ADD_RD2[4]), .Z(n401) );
  MUX2_X1 U417 ( .A(n401), .B(n400), .S(ADD_RD2[3]), .Z(n402) );
  MUX2_X1 U418 ( .A(\REGISTERS[10][11] ), .B(\REGISTERS[26][11] ), .S(
        ADD_RD2[4]), .Z(n403) );
  MUX2_X1 U419 ( .A(\REGISTERS[2][11] ), .B(\REGISTERS[18][11] ), .S(
        ADD_RD2[4]), .Z(n404) );
  MUX2_X1 U420 ( .A(n404), .B(n403), .S(ADD_RD2[3]), .Z(n405) );
  MUX2_X1 U421 ( .A(n405), .B(n402), .S(ADD_RD2[2]), .Z(n406) );
  MUX2_X1 U422 ( .A(n406), .B(n399), .S(ADD_RD2[0]), .Z(n407) );
  MUX2_X1 U423 ( .A(\REGISTERS[13][11] ), .B(\REGISTERS[29][11] ), .S(
        ADD_RD2[4]), .Z(n408) );
  MUX2_X1 U424 ( .A(\REGISTERS[5][11] ), .B(\REGISTERS[21][11] ), .S(
        ADD_RD2[4]), .Z(n409) );
  MUX2_X1 U425 ( .A(n409), .B(n408), .S(ADD_RD2[3]), .Z(n410) );
  MUX2_X1 U426 ( .A(\REGISTERS[9][11] ), .B(\REGISTERS[25][11] ), .S(
        ADD_RD2[4]), .Z(n411) );
  MUX2_X1 U427 ( .A(\REGISTERS[1][11] ), .B(\REGISTERS[17][11] ), .S(
        ADD_RD2[4]), .Z(n412) );
  MUX2_X1 U428 ( .A(n412), .B(n411), .S(ADD_RD2[3]), .Z(n413) );
  MUX2_X1 U429 ( .A(n413), .B(n410), .S(ADD_RD2[2]), .Z(n414) );
  MUX2_X1 U430 ( .A(\REGISTERS[12][11] ), .B(\REGISTERS[28][11] ), .S(
        ADD_RD2[4]), .Z(n415) );
  MUX2_X1 U431 ( .A(\REGISTERS[4][11] ), .B(\REGISTERS[20][11] ), .S(
        ADD_RD2[4]), .Z(n416) );
  MUX2_X1 U432 ( .A(n416), .B(n415), .S(ADD_RD2[3]), .Z(n417) );
  MUX2_X1 U433 ( .A(\REGISTERS[8][11] ), .B(\REGISTERS[24][11] ), .S(
        ADD_RD2[4]), .Z(n418) );
  MUX2_X1 U434 ( .A(\REGISTERS[0][11] ), .B(\REGISTERS[16][11] ), .S(
        ADD_RD2[4]), .Z(n419) );
  MUX2_X1 U435 ( .A(n419), .B(n418), .S(ADD_RD2[3]), .Z(n420) );
  MUX2_X1 U436 ( .A(n420), .B(n417), .S(ADD_RD2[2]), .Z(n421) );
  MUX2_X1 U437 ( .A(n421), .B(n414), .S(ADD_RD2[0]), .Z(n422) );
  MUX2_X1 U438 ( .A(n422), .B(n407), .S(ADD_RD2[1]), .Z(N423) );
  MUX2_X1 U439 ( .A(\REGISTERS[15][12] ), .B(\REGISTERS[31][12] ), .S(
        ADD_RD2[4]), .Z(n423) );
  MUX2_X1 U440 ( .A(\REGISTERS[7][12] ), .B(\REGISTERS[23][12] ), .S(
        ADD_RD2[4]), .Z(n424) );
  MUX2_X1 U441 ( .A(n424), .B(n423), .S(ADD_RD2[3]), .Z(n425) );
  MUX2_X1 U442 ( .A(\REGISTERS[11][12] ), .B(\REGISTERS[27][12] ), .S(
        ADD_RD2[4]), .Z(n426) );
  MUX2_X1 U443 ( .A(\REGISTERS[3][12] ), .B(\REGISTERS[19][12] ), .S(
        ADD_RD2[4]), .Z(n427) );
  MUX2_X1 U444 ( .A(n427), .B(n426), .S(ADD_RD2[3]), .Z(n428) );
  MUX2_X1 U445 ( .A(n428), .B(n425), .S(ADD_RD2[2]), .Z(n429) );
  MUX2_X1 U446 ( .A(\REGISTERS[14][12] ), .B(\REGISTERS[30][12] ), .S(
        ADD_RD2[4]), .Z(n430) );
  MUX2_X1 U447 ( .A(\REGISTERS[6][12] ), .B(\REGISTERS[22][12] ), .S(
        ADD_RD2[4]), .Z(n431) );
  MUX2_X1 U448 ( .A(n431), .B(n430), .S(ADD_RD2[3]), .Z(n432) );
  MUX2_X1 U449 ( .A(\REGISTERS[10][12] ), .B(\REGISTERS[26][12] ), .S(
        ADD_RD2[4]), .Z(n433) );
  MUX2_X1 U450 ( .A(\REGISTERS[2][12] ), .B(\REGISTERS[18][12] ), .S(
        ADD_RD2[4]), .Z(n434) );
  MUX2_X1 U451 ( .A(n434), .B(n433), .S(ADD_RD2[3]), .Z(n435) );
  MUX2_X1 U452 ( .A(n435), .B(n432), .S(ADD_RD2[2]), .Z(n436) );
  MUX2_X1 U453 ( .A(n436), .B(n429), .S(ADD_RD2[0]), .Z(n437) );
  MUX2_X1 U454 ( .A(\REGISTERS[13][12] ), .B(\REGISTERS[29][12] ), .S(
        ADD_RD2[4]), .Z(n438) );
  MUX2_X1 U455 ( .A(\REGISTERS[5][12] ), .B(\REGISTERS[21][12] ), .S(
        ADD_RD2[4]), .Z(n439) );
  MUX2_X1 U456 ( .A(n439), .B(n438), .S(ADD_RD2[3]), .Z(n440) );
  MUX2_X1 U457 ( .A(\REGISTERS[9][12] ), .B(\REGISTERS[25][12] ), .S(
        ADD_RD2[4]), .Z(n441) );
  MUX2_X1 U458 ( .A(\REGISTERS[1][12] ), .B(\REGISTERS[17][12] ), .S(
        ADD_RD2[4]), .Z(n442) );
  MUX2_X1 U459 ( .A(n442), .B(n441), .S(ADD_RD2[3]), .Z(n443) );
  MUX2_X1 U460 ( .A(n443), .B(n440), .S(ADD_RD2[2]), .Z(n444) );
  MUX2_X1 U461 ( .A(\REGISTERS[12][12] ), .B(\REGISTERS[28][12] ), .S(
        ADD_RD2[4]), .Z(n445) );
  MUX2_X1 U462 ( .A(\REGISTERS[4][12] ), .B(\REGISTERS[20][12] ), .S(
        ADD_RD2[4]), .Z(n446) );
  MUX2_X1 U463 ( .A(n446), .B(n445), .S(ADD_RD2[3]), .Z(n447) );
  MUX2_X1 U464 ( .A(\REGISTERS[8][12] ), .B(\REGISTERS[24][12] ), .S(
        ADD_RD2[4]), .Z(n448) );
  MUX2_X1 U465 ( .A(\REGISTERS[0][12] ), .B(\REGISTERS[16][12] ), .S(
        ADD_RD2[4]), .Z(n449) );
  MUX2_X1 U466 ( .A(n449), .B(n448), .S(ADD_RD2[3]), .Z(n450) );
  MUX2_X1 U467 ( .A(n450), .B(n447), .S(ADD_RD2[2]), .Z(n451) );
  MUX2_X1 U468 ( .A(n451), .B(n444), .S(ADD_RD2[0]), .Z(n452) );
  MUX2_X1 U469 ( .A(n452), .B(n437), .S(ADD_RD2[1]), .Z(N424) );
  MUX2_X1 U470 ( .A(\REGISTERS[15][13] ), .B(\REGISTERS[31][13] ), .S(
        ADD_RD2[4]), .Z(n453) );
  MUX2_X1 U471 ( .A(\REGISTERS[7][13] ), .B(\REGISTERS[23][13] ), .S(
        ADD_RD2[4]), .Z(n454) );
  MUX2_X1 U472 ( .A(n454), .B(n453), .S(ADD_RD2[3]), .Z(n455) );
  MUX2_X1 U473 ( .A(\REGISTERS[11][13] ), .B(\REGISTERS[27][13] ), .S(
        ADD_RD2[4]), .Z(n456) );
  MUX2_X1 U474 ( .A(\REGISTERS[3][13] ), .B(\REGISTERS[19][13] ), .S(
        ADD_RD2[4]), .Z(n457) );
  MUX2_X1 U475 ( .A(n457), .B(n456), .S(ADD_RD2[3]), .Z(n458) );
  MUX2_X1 U476 ( .A(n458), .B(n455), .S(ADD_RD2[2]), .Z(n459) );
  MUX2_X1 U477 ( .A(\REGISTERS[14][13] ), .B(\REGISTERS[30][13] ), .S(
        ADD_RD2[4]), .Z(n460) );
  MUX2_X1 U478 ( .A(\REGISTERS[6][13] ), .B(\REGISTERS[22][13] ), .S(
        ADD_RD2[4]), .Z(n461) );
  MUX2_X1 U479 ( .A(n461), .B(n460), .S(ADD_RD2[3]), .Z(n462) );
  MUX2_X1 U480 ( .A(\REGISTERS[10][13] ), .B(\REGISTERS[26][13] ), .S(
        ADD_RD2[4]), .Z(n463) );
  MUX2_X1 U481 ( .A(\REGISTERS[2][13] ), .B(\REGISTERS[18][13] ), .S(
        ADD_RD2[4]), .Z(n464) );
  MUX2_X1 U482 ( .A(n464), .B(n463), .S(ADD_RD2[3]), .Z(n465) );
  MUX2_X1 U483 ( .A(n465), .B(n462), .S(ADD_RD2[2]), .Z(n466) );
  MUX2_X1 U484 ( .A(n466), .B(n459), .S(ADD_RD2[0]), .Z(n467) );
  MUX2_X1 U485 ( .A(\REGISTERS[13][13] ), .B(\REGISTERS[29][13] ), .S(
        ADD_RD2[4]), .Z(n468) );
  MUX2_X1 U486 ( .A(\REGISTERS[5][13] ), .B(\REGISTERS[21][13] ), .S(
        ADD_RD2[4]), .Z(n469) );
  MUX2_X1 U487 ( .A(n469), .B(n468), .S(ADD_RD2[3]), .Z(n470) );
  MUX2_X1 U488 ( .A(\REGISTERS[9][13] ), .B(\REGISTERS[25][13] ), .S(
        ADD_RD2[4]), .Z(n471) );
  MUX2_X1 U489 ( .A(\REGISTERS[1][13] ), .B(\REGISTERS[17][13] ), .S(
        ADD_RD2[4]), .Z(n472) );
  MUX2_X1 U490 ( .A(n472), .B(n471), .S(ADD_RD2[3]), .Z(n473) );
  MUX2_X1 U491 ( .A(n473), .B(n470), .S(ADD_RD2[2]), .Z(n474) );
  MUX2_X1 U492 ( .A(\REGISTERS[12][13] ), .B(\REGISTERS[28][13] ), .S(
        ADD_RD2[4]), .Z(n475) );
  MUX2_X1 U493 ( .A(\REGISTERS[4][13] ), .B(\REGISTERS[20][13] ), .S(
        ADD_RD2[4]), .Z(n476) );
  MUX2_X1 U494 ( .A(n476), .B(n475), .S(ADD_RD2[3]), .Z(n477) );
  MUX2_X1 U495 ( .A(\REGISTERS[8][13] ), .B(\REGISTERS[24][13] ), .S(
        ADD_RD2[4]), .Z(n478) );
  MUX2_X1 U496 ( .A(\REGISTERS[0][13] ), .B(\REGISTERS[16][13] ), .S(
        ADD_RD2[4]), .Z(n479) );
  MUX2_X1 U497 ( .A(n479), .B(n478), .S(ADD_RD2[3]), .Z(n480) );
  MUX2_X1 U498 ( .A(n480), .B(n477), .S(ADD_RD2[2]), .Z(n481) );
  MUX2_X1 U499 ( .A(n481), .B(n474), .S(ADD_RD2[0]), .Z(n482) );
  MUX2_X1 U500 ( .A(n482), .B(n467), .S(ADD_RD2[1]), .Z(N425) );
  MUX2_X1 U501 ( .A(\REGISTERS[15][14] ), .B(\REGISTERS[31][14] ), .S(
        ADD_RD2[4]), .Z(n483) );
  MUX2_X1 U502 ( .A(\REGISTERS[7][14] ), .B(\REGISTERS[23][14] ), .S(
        ADD_RD2[4]), .Z(n484) );
  MUX2_X1 U503 ( .A(n484), .B(n483), .S(ADD_RD2[3]), .Z(n485) );
  MUX2_X1 U504 ( .A(\REGISTERS[11][14] ), .B(\REGISTERS[27][14] ), .S(
        ADD_RD2[4]), .Z(n486) );
  MUX2_X1 U505 ( .A(\REGISTERS[3][14] ), .B(\REGISTERS[19][14] ), .S(
        ADD_RD2[4]), .Z(n487) );
  MUX2_X1 U506 ( .A(n487), .B(n486), .S(ADD_RD2[3]), .Z(n488) );
  MUX2_X1 U507 ( .A(n488), .B(n485), .S(ADD_RD2[2]), .Z(n489) );
  MUX2_X1 U508 ( .A(\REGISTERS[14][14] ), .B(\REGISTERS[30][14] ), .S(
        ADD_RD2[4]), .Z(n490) );
  MUX2_X1 U509 ( .A(\REGISTERS[6][14] ), .B(\REGISTERS[22][14] ), .S(
        ADD_RD2[4]), .Z(n491) );
  MUX2_X1 U510 ( .A(n491), .B(n490), .S(ADD_RD2[3]), .Z(n492) );
  MUX2_X1 U511 ( .A(\REGISTERS[10][14] ), .B(\REGISTERS[26][14] ), .S(
        ADD_RD2[4]), .Z(n493) );
  MUX2_X1 U512 ( .A(\REGISTERS[2][14] ), .B(\REGISTERS[18][14] ), .S(
        ADD_RD2[4]), .Z(n494) );
  MUX2_X1 U513 ( .A(n494), .B(n493), .S(ADD_RD2[3]), .Z(n495) );
  MUX2_X1 U514 ( .A(n495), .B(n492), .S(ADD_RD2[2]), .Z(n496) );
  MUX2_X1 U515 ( .A(n496), .B(n489), .S(ADD_RD2[0]), .Z(n497) );
  MUX2_X1 U516 ( .A(\REGISTERS[13][14] ), .B(\REGISTERS[29][14] ), .S(
        ADD_RD2[4]), .Z(n498) );
  MUX2_X1 U517 ( .A(\REGISTERS[5][14] ), .B(\REGISTERS[21][14] ), .S(
        ADD_RD2[4]), .Z(n499) );
  MUX2_X1 U518 ( .A(n499), .B(n498), .S(ADD_RD2[3]), .Z(n500) );
  MUX2_X1 U519 ( .A(\REGISTERS[9][14] ), .B(\REGISTERS[25][14] ), .S(
        ADD_RD2[4]), .Z(n501) );
  MUX2_X1 U520 ( .A(\REGISTERS[1][14] ), .B(\REGISTERS[17][14] ), .S(
        ADD_RD2[4]), .Z(n502) );
  MUX2_X1 U521 ( .A(n502), .B(n501), .S(ADD_RD2[3]), .Z(n503) );
  MUX2_X1 U522 ( .A(n503), .B(n500), .S(ADD_RD2[2]), .Z(n504) );
  MUX2_X1 U523 ( .A(\REGISTERS[12][14] ), .B(\REGISTERS[28][14] ), .S(
        ADD_RD2[4]), .Z(n505) );
  MUX2_X1 U524 ( .A(\REGISTERS[4][14] ), .B(\REGISTERS[20][14] ), .S(
        ADD_RD2[4]), .Z(n506) );
  MUX2_X1 U525 ( .A(n506), .B(n505), .S(ADD_RD2[3]), .Z(n507) );
  MUX2_X1 U526 ( .A(\REGISTERS[8][14] ), .B(\REGISTERS[24][14] ), .S(
        ADD_RD2[4]), .Z(n508) );
  MUX2_X1 U527 ( .A(\REGISTERS[0][14] ), .B(\REGISTERS[16][14] ), .S(
        ADD_RD2[4]), .Z(n509) );
  MUX2_X1 U528 ( .A(n509), .B(n508), .S(ADD_RD2[3]), .Z(n510) );
  MUX2_X1 U529 ( .A(n510), .B(n507), .S(ADD_RD2[2]), .Z(n511) );
  MUX2_X1 U530 ( .A(n511), .B(n504), .S(ADD_RD2[0]), .Z(n512) );
  MUX2_X1 U531 ( .A(n512), .B(n497), .S(ADD_RD2[1]), .Z(N426) );
  MUX2_X1 U532 ( .A(\REGISTERS[15][15] ), .B(\REGISTERS[31][15] ), .S(
        ADD_RD2[4]), .Z(n513) );
  MUX2_X1 U533 ( .A(\REGISTERS[7][15] ), .B(\REGISTERS[23][15] ), .S(
        ADD_RD2[4]), .Z(n514) );
  MUX2_X1 U534 ( .A(n514), .B(n513), .S(ADD_RD2[3]), .Z(n515) );
  MUX2_X1 U535 ( .A(\REGISTERS[11][15] ), .B(\REGISTERS[27][15] ), .S(
        ADD_RD2[4]), .Z(n516) );
  MUX2_X1 U536 ( .A(\REGISTERS[3][15] ), .B(\REGISTERS[19][15] ), .S(
        ADD_RD2[4]), .Z(n517) );
  MUX2_X1 U537 ( .A(n517), .B(n516), .S(ADD_RD2[3]), .Z(n518) );
  MUX2_X1 U538 ( .A(n518), .B(n515), .S(ADD_RD2[2]), .Z(n519) );
  MUX2_X1 U539 ( .A(\REGISTERS[14][15] ), .B(\REGISTERS[30][15] ), .S(
        ADD_RD2[4]), .Z(n520) );
  MUX2_X1 U540 ( .A(\REGISTERS[6][15] ), .B(\REGISTERS[22][15] ), .S(
        ADD_RD2[4]), .Z(n521) );
  MUX2_X1 U541 ( .A(n521), .B(n520), .S(ADD_RD2[3]), .Z(n522) );
  MUX2_X1 U542 ( .A(\REGISTERS[10][15] ), .B(\REGISTERS[26][15] ), .S(
        ADD_RD2[4]), .Z(n523) );
  MUX2_X1 U543 ( .A(\REGISTERS[2][15] ), .B(\REGISTERS[18][15] ), .S(
        ADD_RD2[4]), .Z(n524) );
  MUX2_X1 U544 ( .A(n524), .B(n523), .S(ADD_RD2[3]), .Z(n525) );
  MUX2_X1 U545 ( .A(n525), .B(n522), .S(ADD_RD2[2]), .Z(n526) );
  MUX2_X1 U546 ( .A(n526), .B(n519), .S(ADD_RD2[0]), .Z(n527) );
  MUX2_X1 U547 ( .A(\REGISTERS[13][15] ), .B(\REGISTERS[29][15] ), .S(
        ADD_RD2[4]), .Z(n528) );
  MUX2_X1 U548 ( .A(\REGISTERS[5][15] ), .B(\REGISTERS[21][15] ), .S(
        ADD_RD2[4]), .Z(n529) );
  MUX2_X1 U549 ( .A(n529), .B(n528), .S(ADD_RD2[3]), .Z(n530) );
  MUX2_X1 U550 ( .A(\REGISTERS[9][15] ), .B(\REGISTERS[25][15] ), .S(
        ADD_RD2[4]), .Z(n531) );
  MUX2_X1 U551 ( .A(\REGISTERS[1][15] ), .B(\REGISTERS[17][15] ), .S(
        ADD_RD2[4]), .Z(n532) );
  MUX2_X1 U552 ( .A(n532), .B(n531), .S(ADD_RD2[3]), .Z(n533) );
  MUX2_X1 U553 ( .A(n533), .B(n530), .S(ADD_RD2[2]), .Z(n534) );
  MUX2_X1 U554 ( .A(\REGISTERS[12][15] ), .B(\REGISTERS[28][15] ), .S(
        ADD_RD2[4]), .Z(n535) );
  MUX2_X1 U555 ( .A(\REGISTERS[4][15] ), .B(\REGISTERS[20][15] ), .S(
        ADD_RD2[4]), .Z(n536) );
  MUX2_X1 U556 ( .A(n536), .B(n535), .S(ADD_RD2[3]), .Z(n537) );
  MUX2_X1 U557 ( .A(\REGISTERS[8][15] ), .B(\REGISTERS[24][15] ), .S(
        ADD_RD2[4]), .Z(n538) );
  MUX2_X1 U558 ( .A(\REGISTERS[0][15] ), .B(\REGISTERS[16][15] ), .S(
        ADD_RD2[4]), .Z(n539) );
  MUX2_X1 U559 ( .A(n539), .B(n538), .S(ADD_RD2[3]), .Z(n540) );
  MUX2_X1 U560 ( .A(n540), .B(n537), .S(ADD_RD2[2]), .Z(n541) );
  MUX2_X1 U561 ( .A(n541), .B(n534), .S(ADD_RD2[0]), .Z(n542) );
  MUX2_X1 U562 ( .A(n542), .B(n527), .S(ADD_RD2[1]), .Z(N427) );
  MUX2_X1 U563 ( .A(\REGISTERS[15][16] ), .B(\REGISTERS[31][16] ), .S(
        ADD_RD2[4]), .Z(n543) );
  MUX2_X1 U564 ( .A(\REGISTERS[7][16] ), .B(\REGISTERS[23][16] ), .S(
        ADD_RD2[4]), .Z(n544) );
  MUX2_X1 U565 ( .A(n544), .B(n543), .S(ADD_RD2[3]), .Z(n545) );
  MUX2_X1 U566 ( .A(\REGISTERS[11][16] ), .B(\REGISTERS[27][16] ), .S(
        ADD_RD2[4]), .Z(n546) );
  MUX2_X1 U567 ( .A(\REGISTERS[3][16] ), .B(\REGISTERS[19][16] ), .S(
        ADD_RD2[4]), .Z(n547) );
  MUX2_X1 U568 ( .A(n547), .B(n546), .S(ADD_RD2[3]), .Z(n548) );
  MUX2_X1 U569 ( .A(n548), .B(n545), .S(ADD_RD2[2]), .Z(n549) );
  MUX2_X1 U570 ( .A(\REGISTERS[14][16] ), .B(\REGISTERS[30][16] ), .S(
        ADD_RD2[4]), .Z(n550) );
  MUX2_X1 U571 ( .A(\REGISTERS[6][16] ), .B(\REGISTERS[22][16] ), .S(
        ADD_RD2[4]), .Z(n551) );
  MUX2_X1 U572 ( .A(n551), .B(n550), .S(ADD_RD2[3]), .Z(n552) );
  MUX2_X1 U573 ( .A(\REGISTERS[10][16] ), .B(\REGISTERS[26][16] ), .S(
        ADD_RD2[4]), .Z(n553) );
  MUX2_X1 U574 ( .A(\REGISTERS[2][16] ), .B(\REGISTERS[18][16] ), .S(
        ADD_RD2[4]), .Z(n554) );
  MUX2_X1 U575 ( .A(n554), .B(n553), .S(ADD_RD2[3]), .Z(n555) );
  MUX2_X1 U576 ( .A(n555), .B(n552), .S(ADD_RD2[2]), .Z(n556) );
  MUX2_X1 U577 ( .A(n556), .B(n549), .S(ADD_RD2[0]), .Z(n557) );
  MUX2_X1 U578 ( .A(\REGISTERS[13][16] ), .B(\REGISTERS[29][16] ), .S(
        ADD_RD2[4]), .Z(n558) );
  MUX2_X1 U579 ( .A(\REGISTERS[5][16] ), .B(\REGISTERS[21][16] ), .S(
        ADD_RD2[4]), .Z(n559) );
  MUX2_X1 U580 ( .A(n559), .B(n558), .S(ADD_RD2[3]), .Z(n560) );
  MUX2_X1 U581 ( .A(\REGISTERS[9][16] ), .B(\REGISTERS[25][16] ), .S(
        ADD_RD2[4]), .Z(n561) );
  MUX2_X1 U582 ( .A(\REGISTERS[1][16] ), .B(\REGISTERS[17][16] ), .S(
        ADD_RD2[4]), .Z(n562) );
  MUX2_X1 U583 ( .A(n562), .B(n561), .S(ADD_RD2[3]), .Z(n563) );
  MUX2_X1 U584 ( .A(n563), .B(n560), .S(ADD_RD2[2]), .Z(n564) );
  MUX2_X1 U585 ( .A(\REGISTERS[12][16] ), .B(\REGISTERS[28][16] ), .S(
        ADD_RD2[4]), .Z(n565) );
  MUX2_X1 U586 ( .A(\REGISTERS[4][16] ), .B(\REGISTERS[20][16] ), .S(
        ADD_RD2[4]), .Z(n566) );
  MUX2_X1 U587 ( .A(n566), .B(n565), .S(ADD_RD2[3]), .Z(n567) );
  MUX2_X1 U588 ( .A(\REGISTERS[8][16] ), .B(\REGISTERS[24][16] ), .S(
        ADD_RD2[4]), .Z(n568) );
  MUX2_X1 U589 ( .A(\REGISTERS[0][16] ), .B(\REGISTERS[16][16] ), .S(
        ADD_RD2[4]), .Z(n569) );
  MUX2_X1 U590 ( .A(n569), .B(n568), .S(ADD_RD2[3]), .Z(n570) );
  MUX2_X1 U591 ( .A(n570), .B(n567), .S(ADD_RD2[2]), .Z(n571) );
  MUX2_X1 U592 ( .A(n571), .B(n564), .S(ADD_RD2[0]), .Z(n572) );
  MUX2_X1 U593 ( .A(n572), .B(n557), .S(ADD_RD2[1]), .Z(N428) );
  MUX2_X1 U594 ( .A(\REGISTERS[15][17] ), .B(\REGISTERS[31][17] ), .S(
        ADD_RD2[4]), .Z(n573) );
  MUX2_X1 U595 ( .A(\REGISTERS[7][17] ), .B(\REGISTERS[23][17] ), .S(
        ADD_RD2[4]), .Z(n574) );
  MUX2_X1 U596 ( .A(n574), .B(n573), .S(ADD_RD2[3]), .Z(n575) );
  MUX2_X1 U597 ( .A(\REGISTERS[11][17] ), .B(\REGISTERS[27][17] ), .S(
        ADD_RD2[4]), .Z(n576) );
  MUX2_X1 U598 ( .A(\REGISTERS[3][17] ), .B(\REGISTERS[19][17] ), .S(
        ADD_RD2[4]), .Z(n577) );
  MUX2_X1 U599 ( .A(n577), .B(n576), .S(ADD_RD2[3]), .Z(n578) );
  MUX2_X1 U600 ( .A(n578), .B(n575), .S(ADD_RD2[2]), .Z(n579) );
  MUX2_X1 U601 ( .A(\REGISTERS[14][17] ), .B(\REGISTERS[30][17] ), .S(
        ADD_RD2[4]), .Z(n580) );
  MUX2_X1 U602 ( .A(\REGISTERS[6][17] ), .B(\REGISTERS[22][17] ), .S(
        ADD_RD2[4]), .Z(n581) );
  MUX2_X1 U603 ( .A(n581), .B(n580), .S(ADD_RD2[3]), .Z(n582) );
  MUX2_X1 U604 ( .A(\REGISTERS[10][17] ), .B(\REGISTERS[26][17] ), .S(
        ADD_RD2[4]), .Z(n583) );
  MUX2_X1 U605 ( .A(\REGISTERS[2][17] ), .B(\REGISTERS[18][17] ), .S(
        ADD_RD2[4]), .Z(n584) );
  MUX2_X1 U606 ( .A(n584), .B(n583), .S(ADD_RD2[3]), .Z(n585) );
  MUX2_X1 U607 ( .A(n585), .B(n582), .S(ADD_RD2[2]), .Z(n586) );
  MUX2_X1 U608 ( .A(n586), .B(n579), .S(ADD_RD2[0]), .Z(n587) );
  MUX2_X1 U609 ( .A(\REGISTERS[13][17] ), .B(\REGISTERS[29][17] ), .S(
        ADD_RD2[4]), .Z(n588) );
  MUX2_X1 U610 ( .A(\REGISTERS[5][17] ), .B(\REGISTERS[21][17] ), .S(
        ADD_RD2[4]), .Z(n589) );
  MUX2_X1 U611 ( .A(n589), .B(n588), .S(ADD_RD2[3]), .Z(n590) );
  MUX2_X1 U612 ( .A(\REGISTERS[9][17] ), .B(\REGISTERS[25][17] ), .S(
        ADD_RD2[4]), .Z(n591) );
  MUX2_X1 U613 ( .A(\REGISTERS[1][17] ), .B(\REGISTERS[17][17] ), .S(
        ADD_RD2[4]), .Z(n592) );
  MUX2_X1 U614 ( .A(n592), .B(n591), .S(ADD_RD2[3]), .Z(n593) );
  MUX2_X1 U615 ( .A(n593), .B(n590), .S(ADD_RD2[2]), .Z(n594) );
  MUX2_X1 U616 ( .A(\REGISTERS[12][17] ), .B(\REGISTERS[28][17] ), .S(
        ADD_RD2[4]), .Z(n595) );
  MUX2_X1 U617 ( .A(\REGISTERS[4][17] ), .B(\REGISTERS[20][17] ), .S(
        ADD_RD2[4]), .Z(n596) );
  MUX2_X1 U618 ( .A(n596), .B(n595), .S(ADD_RD2[3]), .Z(n597) );
  MUX2_X1 U619 ( .A(\REGISTERS[8][17] ), .B(\REGISTERS[24][17] ), .S(
        ADD_RD2[4]), .Z(n598) );
  MUX2_X1 U620 ( .A(\REGISTERS[0][17] ), .B(\REGISTERS[16][17] ), .S(
        ADD_RD2[4]), .Z(n599) );
  MUX2_X1 U621 ( .A(n599), .B(n598), .S(ADD_RD2[3]), .Z(n600) );
  MUX2_X1 U622 ( .A(n600), .B(n597), .S(ADD_RD2[2]), .Z(n601) );
  MUX2_X1 U623 ( .A(n601), .B(n594), .S(ADD_RD2[0]), .Z(n602) );
  MUX2_X1 U624 ( .A(n602), .B(n587), .S(ADD_RD2[1]), .Z(N429) );
  MUX2_X1 U625 ( .A(\REGISTERS[15][18] ), .B(\REGISTERS[31][18] ), .S(
        ADD_RD2[4]), .Z(n603) );
  MUX2_X1 U626 ( .A(\REGISTERS[7][18] ), .B(\REGISTERS[23][18] ), .S(
        ADD_RD2[4]), .Z(n604) );
  MUX2_X1 U627 ( .A(n604), .B(n603), .S(ADD_RD2[3]), .Z(n605) );
  MUX2_X1 U628 ( .A(\REGISTERS[11][18] ), .B(\REGISTERS[27][18] ), .S(
        ADD_RD2[4]), .Z(n606) );
  MUX2_X1 U629 ( .A(\REGISTERS[3][18] ), .B(\REGISTERS[19][18] ), .S(
        ADD_RD2[4]), .Z(n607) );
  MUX2_X1 U630 ( .A(n607), .B(n606), .S(ADD_RD2[3]), .Z(n608) );
  MUX2_X1 U631 ( .A(n608), .B(n605), .S(ADD_RD2[2]), .Z(n609) );
  MUX2_X1 U632 ( .A(\REGISTERS[14][18] ), .B(\REGISTERS[30][18] ), .S(
        ADD_RD2[4]), .Z(n610) );
  MUX2_X1 U633 ( .A(\REGISTERS[6][18] ), .B(\REGISTERS[22][18] ), .S(
        ADD_RD2[4]), .Z(n611) );
  MUX2_X1 U634 ( .A(n611), .B(n610), .S(ADD_RD2[3]), .Z(n612) );
  MUX2_X1 U635 ( .A(\REGISTERS[10][18] ), .B(\REGISTERS[26][18] ), .S(
        ADD_RD2[4]), .Z(n613) );
  MUX2_X1 U636 ( .A(\REGISTERS[2][18] ), .B(\REGISTERS[18][18] ), .S(
        ADD_RD2[4]), .Z(n614) );
  MUX2_X1 U637 ( .A(n614), .B(n613), .S(ADD_RD2[3]), .Z(n615) );
  MUX2_X1 U638 ( .A(n615), .B(n612), .S(ADD_RD2[2]), .Z(n616) );
  MUX2_X1 U639 ( .A(n616), .B(n609), .S(ADD_RD2[0]), .Z(n617) );
  MUX2_X1 U640 ( .A(\REGISTERS[13][18] ), .B(\REGISTERS[29][18] ), .S(
        ADD_RD2[4]), .Z(n618) );
  MUX2_X1 U641 ( .A(\REGISTERS[5][18] ), .B(\REGISTERS[21][18] ), .S(
        ADD_RD2[4]), .Z(n619) );
  MUX2_X1 U642 ( .A(n619), .B(n618), .S(ADD_RD2[3]), .Z(n620) );
  MUX2_X1 U643 ( .A(\REGISTERS[9][18] ), .B(\REGISTERS[25][18] ), .S(
        ADD_RD2[4]), .Z(n621) );
  MUX2_X1 U644 ( .A(\REGISTERS[1][18] ), .B(\REGISTERS[17][18] ), .S(
        ADD_RD2[4]), .Z(n622) );
  MUX2_X1 U645 ( .A(n622), .B(n621), .S(ADD_RD2[3]), .Z(n623) );
  MUX2_X1 U646 ( .A(n623), .B(n620), .S(ADD_RD2[2]), .Z(n624) );
  MUX2_X1 U647 ( .A(\REGISTERS[12][18] ), .B(\REGISTERS[28][18] ), .S(
        ADD_RD2[4]), .Z(n625) );
  MUX2_X1 U648 ( .A(\REGISTERS[4][18] ), .B(\REGISTERS[20][18] ), .S(
        ADD_RD2[4]), .Z(n626) );
  MUX2_X1 U649 ( .A(n626), .B(n625), .S(ADD_RD2[3]), .Z(n627) );
  MUX2_X1 U650 ( .A(\REGISTERS[8][18] ), .B(\REGISTERS[24][18] ), .S(
        ADD_RD2[4]), .Z(n628) );
  MUX2_X1 U651 ( .A(\REGISTERS[0][18] ), .B(\REGISTERS[16][18] ), .S(
        ADD_RD2[4]), .Z(n629) );
  MUX2_X1 U652 ( .A(n629), .B(n628), .S(ADD_RD2[3]), .Z(n630) );
  MUX2_X1 U653 ( .A(n630), .B(n627), .S(ADD_RD2[2]), .Z(n631) );
  MUX2_X1 U654 ( .A(n631), .B(n624), .S(ADD_RD2[0]), .Z(n632) );
  MUX2_X1 U655 ( .A(n632), .B(n617), .S(ADD_RD2[1]), .Z(N430) );
  MUX2_X1 U656 ( .A(\REGISTERS[15][19] ), .B(\REGISTERS[31][19] ), .S(
        ADD_RD2[4]), .Z(n633) );
  MUX2_X1 U657 ( .A(\REGISTERS[7][19] ), .B(\REGISTERS[23][19] ), .S(
        ADD_RD2[4]), .Z(n634) );
  MUX2_X1 U658 ( .A(n634), .B(n633), .S(ADD_RD2[3]), .Z(n635) );
  MUX2_X1 U659 ( .A(\REGISTERS[11][19] ), .B(\REGISTERS[27][19] ), .S(
        ADD_RD2[4]), .Z(n636) );
  MUX2_X1 U660 ( .A(\REGISTERS[3][19] ), .B(\REGISTERS[19][19] ), .S(
        ADD_RD2[4]), .Z(n637) );
  MUX2_X1 U661 ( .A(n637), .B(n636), .S(ADD_RD2[3]), .Z(n638) );
  MUX2_X1 U662 ( .A(n638), .B(n635), .S(ADD_RD2[2]), .Z(n639) );
  MUX2_X1 U663 ( .A(\REGISTERS[14][19] ), .B(\REGISTERS[30][19] ), .S(
        ADD_RD2[4]), .Z(n640) );
  MUX2_X1 U664 ( .A(\REGISTERS[6][19] ), .B(\REGISTERS[22][19] ), .S(
        ADD_RD2[4]), .Z(n641) );
  MUX2_X1 U665 ( .A(n641), .B(n640), .S(ADD_RD2[3]), .Z(n642) );
  MUX2_X1 U666 ( .A(\REGISTERS[10][19] ), .B(\REGISTERS[26][19] ), .S(
        ADD_RD2[4]), .Z(n643) );
  MUX2_X1 U667 ( .A(\REGISTERS[2][19] ), .B(\REGISTERS[18][19] ), .S(
        ADD_RD2[4]), .Z(n644) );
  MUX2_X1 U668 ( .A(n644), .B(n643), .S(ADD_RD2[3]), .Z(n645) );
  MUX2_X1 U669 ( .A(n645), .B(n642), .S(ADD_RD2[2]), .Z(n646) );
  MUX2_X1 U670 ( .A(n646), .B(n639), .S(ADD_RD2[0]), .Z(n647) );
  MUX2_X1 U671 ( .A(\REGISTERS[13][19] ), .B(\REGISTERS[29][19] ), .S(
        ADD_RD2[4]), .Z(n648) );
  MUX2_X1 U672 ( .A(\REGISTERS[5][19] ), .B(\REGISTERS[21][19] ), .S(
        ADD_RD2[4]), .Z(n649) );
  MUX2_X1 U673 ( .A(n649), .B(n648), .S(ADD_RD2[3]), .Z(n650) );
  MUX2_X1 U674 ( .A(\REGISTERS[9][19] ), .B(\REGISTERS[25][19] ), .S(
        ADD_RD2[4]), .Z(n651) );
  MUX2_X1 U675 ( .A(\REGISTERS[1][19] ), .B(\REGISTERS[17][19] ), .S(
        ADD_RD2[4]), .Z(n652) );
  MUX2_X1 U676 ( .A(n652), .B(n651), .S(ADD_RD2[3]), .Z(n653) );
  MUX2_X1 U677 ( .A(n653), .B(n650), .S(ADD_RD2[2]), .Z(n654) );
  MUX2_X1 U678 ( .A(\REGISTERS[12][19] ), .B(\REGISTERS[28][19] ), .S(
        ADD_RD2[4]), .Z(n655) );
  MUX2_X1 U679 ( .A(\REGISTERS[4][19] ), .B(\REGISTERS[20][19] ), .S(
        ADD_RD2[4]), .Z(n656) );
  MUX2_X1 U680 ( .A(n656), .B(n655), .S(ADD_RD2[3]), .Z(n657) );
  MUX2_X1 U681 ( .A(\REGISTERS[8][19] ), .B(\REGISTERS[24][19] ), .S(
        ADD_RD2[4]), .Z(n658) );
  MUX2_X1 U682 ( .A(\REGISTERS[0][19] ), .B(\REGISTERS[16][19] ), .S(
        ADD_RD2[4]), .Z(n659) );
  MUX2_X1 U683 ( .A(n659), .B(n658), .S(ADD_RD2[3]), .Z(n660) );
  MUX2_X1 U684 ( .A(n660), .B(n657), .S(ADD_RD2[2]), .Z(n661) );
  MUX2_X1 U685 ( .A(n661), .B(n654), .S(ADD_RD2[0]), .Z(n662) );
  MUX2_X1 U686 ( .A(n662), .B(n647), .S(ADD_RD2[1]), .Z(N431) );
  MUX2_X1 U687 ( .A(\REGISTERS[15][20] ), .B(\REGISTERS[31][20] ), .S(
        ADD_RD2[4]), .Z(n663) );
  MUX2_X1 U688 ( .A(\REGISTERS[7][20] ), .B(\REGISTERS[23][20] ), .S(
        ADD_RD2[4]), .Z(n664) );
  MUX2_X1 U689 ( .A(n664), .B(n663), .S(ADD_RD2[3]), .Z(n665) );
  MUX2_X1 U690 ( .A(\REGISTERS[11][20] ), .B(\REGISTERS[27][20] ), .S(
        ADD_RD2[4]), .Z(n666) );
  MUX2_X1 U691 ( .A(\REGISTERS[3][20] ), .B(\REGISTERS[19][20] ), .S(
        ADD_RD2[4]), .Z(n667) );
  MUX2_X1 U692 ( .A(n667), .B(n666), .S(ADD_RD2[3]), .Z(n668) );
  MUX2_X1 U693 ( .A(n668), .B(n665), .S(ADD_RD2[2]), .Z(n669) );
  MUX2_X1 U694 ( .A(\REGISTERS[14][20] ), .B(\REGISTERS[30][20] ), .S(
        ADD_RD2[4]), .Z(n670) );
  MUX2_X1 U695 ( .A(\REGISTERS[6][20] ), .B(\REGISTERS[22][20] ), .S(
        ADD_RD2[4]), .Z(n671) );
  MUX2_X1 U696 ( .A(n671), .B(n670), .S(ADD_RD2[3]), .Z(n672) );
  MUX2_X1 U697 ( .A(\REGISTERS[10][20] ), .B(\REGISTERS[26][20] ), .S(
        ADD_RD2[4]), .Z(n673) );
  MUX2_X1 U698 ( .A(\REGISTERS[2][20] ), .B(\REGISTERS[18][20] ), .S(
        ADD_RD2[4]), .Z(n674) );
  MUX2_X1 U699 ( .A(n674), .B(n673), .S(ADD_RD2[3]), .Z(n675) );
  MUX2_X1 U700 ( .A(n675), .B(n672), .S(ADD_RD2[2]), .Z(n676) );
  MUX2_X1 U701 ( .A(n676), .B(n669), .S(ADD_RD2[0]), .Z(n677) );
  MUX2_X1 U702 ( .A(\REGISTERS[13][20] ), .B(\REGISTERS[29][20] ), .S(
        ADD_RD2[4]), .Z(n678) );
  MUX2_X1 U703 ( .A(\REGISTERS[5][20] ), .B(\REGISTERS[21][20] ), .S(
        ADD_RD2[4]), .Z(n679) );
  MUX2_X1 U704 ( .A(n679), .B(n678), .S(ADD_RD2[3]), .Z(n680) );
  MUX2_X1 U705 ( .A(\REGISTERS[9][20] ), .B(\REGISTERS[25][20] ), .S(
        ADD_RD2[4]), .Z(n681) );
  MUX2_X1 U706 ( .A(\REGISTERS[1][20] ), .B(\REGISTERS[17][20] ), .S(
        ADD_RD2[4]), .Z(n682) );
  MUX2_X1 U707 ( .A(n682), .B(n681), .S(ADD_RD2[3]), .Z(n683) );
  MUX2_X1 U708 ( .A(n683), .B(n680), .S(ADD_RD2[2]), .Z(n684) );
  MUX2_X1 U709 ( .A(\REGISTERS[12][20] ), .B(\REGISTERS[28][20] ), .S(
        ADD_RD2[4]), .Z(n685) );
  MUX2_X1 U710 ( .A(\REGISTERS[4][20] ), .B(\REGISTERS[20][20] ), .S(
        ADD_RD2[4]), .Z(n686) );
  MUX2_X1 U711 ( .A(n686), .B(n685), .S(ADD_RD2[3]), .Z(n687) );
  MUX2_X1 U712 ( .A(\REGISTERS[8][20] ), .B(\REGISTERS[24][20] ), .S(
        ADD_RD2[4]), .Z(n688) );
  MUX2_X1 U713 ( .A(\REGISTERS[0][20] ), .B(\REGISTERS[16][20] ), .S(
        ADD_RD2[4]), .Z(n689) );
  MUX2_X1 U714 ( .A(n689), .B(n688), .S(ADD_RD2[3]), .Z(n690) );
  MUX2_X1 U715 ( .A(n690), .B(n687), .S(ADD_RD2[2]), .Z(n691) );
  MUX2_X1 U716 ( .A(n691), .B(n684), .S(ADD_RD2[0]), .Z(n692) );
  MUX2_X1 U717 ( .A(n692), .B(n677), .S(ADD_RD2[1]), .Z(N432) );
  MUX2_X1 U718 ( .A(\REGISTERS[15][21] ), .B(\REGISTERS[31][21] ), .S(
        ADD_RD2[4]), .Z(n693) );
  MUX2_X1 U719 ( .A(\REGISTERS[7][21] ), .B(\REGISTERS[23][21] ), .S(
        ADD_RD2[4]), .Z(n694) );
  MUX2_X1 U720 ( .A(n694), .B(n693), .S(ADD_RD2[3]), .Z(n695) );
  MUX2_X1 U721 ( .A(\REGISTERS[11][21] ), .B(\REGISTERS[27][21] ), .S(
        ADD_RD2[4]), .Z(n696) );
  MUX2_X1 U722 ( .A(\REGISTERS[3][21] ), .B(\REGISTERS[19][21] ), .S(
        ADD_RD2[4]), .Z(n697) );
  MUX2_X1 U723 ( .A(n697), .B(n696), .S(ADD_RD2[3]), .Z(n698) );
  MUX2_X1 U724 ( .A(n698), .B(n695), .S(ADD_RD2[2]), .Z(n699) );
  MUX2_X1 U725 ( .A(\REGISTERS[14][21] ), .B(\REGISTERS[30][21] ), .S(
        ADD_RD2[4]), .Z(n700) );
  MUX2_X1 U726 ( .A(\REGISTERS[6][21] ), .B(\REGISTERS[22][21] ), .S(
        ADD_RD2[4]), .Z(n701) );
  MUX2_X1 U727 ( .A(n701), .B(n700), .S(ADD_RD2[3]), .Z(n702) );
  MUX2_X1 U728 ( .A(\REGISTERS[10][21] ), .B(\REGISTERS[26][21] ), .S(
        ADD_RD2[4]), .Z(n703) );
  MUX2_X1 U729 ( .A(\REGISTERS[2][21] ), .B(\REGISTERS[18][21] ), .S(
        ADD_RD2[4]), .Z(n704) );
  MUX2_X1 U730 ( .A(n704), .B(n703), .S(ADD_RD2[3]), .Z(n705) );
  MUX2_X1 U731 ( .A(n705), .B(n702), .S(ADD_RD2[2]), .Z(n706) );
  MUX2_X1 U732 ( .A(n706), .B(n699), .S(ADD_RD2[0]), .Z(n707) );
  MUX2_X1 U733 ( .A(\REGISTERS[13][21] ), .B(\REGISTERS[29][21] ), .S(
        ADD_RD2[4]), .Z(n708) );
  MUX2_X1 U734 ( .A(\REGISTERS[5][21] ), .B(\REGISTERS[21][21] ), .S(
        ADD_RD2[4]), .Z(n709) );
  MUX2_X1 U735 ( .A(n709), .B(n708), .S(ADD_RD2[3]), .Z(n710) );
  MUX2_X1 U736 ( .A(\REGISTERS[9][21] ), .B(\REGISTERS[25][21] ), .S(
        ADD_RD2[4]), .Z(n711) );
  MUX2_X1 U737 ( .A(\REGISTERS[1][21] ), .B(\REGISTERS[17][21] ), .S(
        ADD_RD2[4]), .Z(n712) );
  MUX2_X1 U738 ( .A(n712), .B(n711), .S(ADD_RD2[3]), .Z(n713) );
  MUX2_X1 U739 ( .A(n713), .B(n710), .S(ADD_RD2[2]), .Z(n714) );
  MUX2_X1 U740 ( .A(\REGISTERS[12][21] ), .B(\REGISTERS[28][21] ), .S(
        ADD_RD2[4]), .Z(n715) );
  MUX2_X1 U741 ( .A(\REGISTERS[4][21] ), .B(\REGISTERS[20][21] ), .S(
        ADD_RD2[4]), .Z(n716) );
  MUX2_X1 U742 ( .A(n716), .B(n715), .S(ADD_RD2[3]), .Z(n717) );
  MUX2_X1 U743 ( .A(\REGISTERS[8][21] ), .B(\REGISTERS[24][21] ), .S(
        ADD_RD2[4]), .Z(n718) );
  MUX2_X1 U744 ( .A(\REGISTERS[0][21] ), .B(\REGISTERS[16][21] ), .S(
        ADD_RD2[4]), .Z(n719) );
  MUX2_X1 U745 ( .A(n719), .B(n718), .S(ADD_RD2[3]), .Z(n720) );
  MUX2_X1 U746 ( .A(n720), .B(n717), .S(ADD_RD2[2]), .Z(n721) );
  MUX2_X1 U747 ( .A(n721), .B(n714), .S(ADD_RD2[0]), .Z(n722) );
  MUX2_X1 U748 ( .A(n722), .B(n707), .S(ADD_RD2[1]), .Z(N433) );
  MUX2_X1 U749 ( .A(\REGISTERS[15][22] ), .B(\REGISTERS[31][22] ), .S(
        ADD_RD2[4]), .Z(n723) );
  MUX2_X1 U750 ( .A(\REGISTERS[7][22] ), .B(\REGISTERS[23][22] ), .S(
        ADD_RD2[4]), .Z(n724) );
  MUX2_X1 U751 ( .A(n724), .B(n723), .S(ADD_RD2[3]), .Z(n725) );
  MUX2_X1 U752 ( .A(\REGISTERS[11][22] ), .B(\REGISTERS[27][22] ), .S(
        ADD_RD2[4]), .Z(n726) );
  MUX2_X1 U753 ( .A(\REGISTERS[3][22] ), .B(\REGISTERS[19][22] ), .S(
        ADD_RD2[4]), .Z(n727) );
  MUX2_X1 U754 ( .A(n727), .B(n726), .S(ADD_RD2[3]), .Z(n728) );
  MUX2_X1 U755 ( .A(n728), .B(n725), .S(ADD_RD2[2]), .Z(n729) );
  MUX2_X1 U756 ( .A(\REGISTERS[14][22] ), .B(\REGISTERS[30][22] ), .S(
        ADD_RD2[4]), .Z(n730) );
  MUX2_X1 U757 ( .A(\REGISTERS[6][22] ), .B(\REGISTERS[22][22] ), .S(
        ADD_RD2[4]), .Z(n731) );
  MUX2_X1 U758 ( .A(n731), .B(n730), .S(ADD_RD2[3]), .Z(n732) );
  MUX2_X1 U759 ( .A(\REGISTERS[10][22] ), .B(\REGISTERS[26][22] ), .S(
        ADD_RD2[4]), .Z(n733) );
  MUX2_X1 U760 ( .A(\REGISTERS[2][22] ), .B(\REGISTERS[18][22] ), .S(
        ADD_RD2[4]), .Z(n734) );
  MUX2_X1 U761 ( .A(n734), .B(n733), .S(ADD_RD2[3]), .Z(n735) );
  MUX2_X1 U762 ( .A(n735), .B(n732), .S(ADD_RD2[2]), .Z(n736) );
  MUX2_X1 U763 ( .A(n736), .B(n729), .S(ADD_RD2[0]), .Z(n737) );
  MUX2_X1 U764 ( .A(\REGISTERS[13][22] ), .B(\REGISTERS[29][22] ), .S(
        ADD_RD2[4]), .Z(n738) );
  MUX2_X1 U765 ( .A(\REGISTERS[5][22] ), .B(\REGISTERS[21][22] ), .S(
        ADD_RD2[4]), .Z(n739) );
  MUX2_X1 U766 ( .A(n739), .B(n738), .S(ADD_RD2[3]), .Z(n740) );
  MUX2_X1 U767 ( .A(\REGISTERS[9][22] ), .B(\REGISTERS[25][22] ), .S(
        ADD_RD2[4]), .Z(n741) );
  MUX2_X1 U768 ( .A(\REGISTERS[1][22] ), .B(\REGISTERS[17][22] ), .S(
        ADD_RD2[4]), .Z(n742) );
  MUX2_X1 U769 ( .A(n742), .B(n741), .S(ADD_RD2[3]), .Z(n743) );
  MUX2_X1 U770 ( .A(n743), .B(n740), .S(ADD_RD2[2]), .Z(n744) );
  MUX2_X1 U771 ( .A(\REGISTERS[12][22] ), .B(\REGISTERS[28][22] ), .S(
        ADD_RD2[4]), .Z(n745) );
  MUX2_X1 U772 ( .A(\REGISTERS[4][22] ), .B(\REGISTERS[20][22] ), .S(
        ADD_RD2[4]), .Z(n746) );
  MUX2_X1 U773 ( .A(n746), .B(n745), .S(ADD_RD2[3]), .Z(n747) );
  MUX2_X1 U774 ( .A(\REGISTERS[8][22] ), .B(\REGISTERS[24][22] ), .S(
        ADD_RD2[4]), .Z(n748) );
  MUX2_X1 U775 ( .A(\REGISTERS[0][22] ), .B(\REGISTERS[16][22] ), .S(
        ADD_RD2[4]), .Z(n749) );
  MUX2_X1 U776 ( .A(n749), .B(n748), .S(ADD_RD2[3]), .Z(n750) );
  MUX2_X1 U777 ( .A(n750), .B(n747), .S(ADD_RD2[2]), .Z(n751) );
  MUX2_X1 U778 ( .A(n751), .B(n744), .S(ADD_RD2[0]), .Z(n752) );
  MUX2_X1 U779 ( .A(n752), .B(n737), .S(ADD_RD2[1]), .Z(N434) );
  MUX2_X1 U780 ( .A(\REGISTERS[15][23] ), .B(\REGISTERS[31][23] ), .S(
        ADD_RD2[4]), .Z(n753) );
  MUX2_X1 U781 ( .A(\REGISTERS[7][23] ), .B(\REGISTERS[23][23] ), .S(
        ADD_RD2[4]), .Z(n754) );
  MUX2_X1 U782 ( .A(n754), .B(n753), .S(ADD_RD2[3]), .Z(n755) );
  MUX2_X1 U783 ( .A(\REGISTERS[11][23] ), .B(\REGISTERS[27][23] ), .S(
        ADD_RD2[4]), .Z(n756) );
  MUX2_X1 U784 ( .A(\REGISTERS[3][23] ), .B(\REGISTERS[19][23] ), .S(
        ADD_RD2[4]), .Z(n757) );
  MUX2_X1 U785 ( .A(n757), .B(n756), .S(ADD_RD2[3]), .Z(n758) );
  MUX2_X1 U786 ( .A(n758), .B(n755), .S(ADD_RD2[2]), .Z(n759) );
  MUX2_X1 U787 ( .A(\REGISTERS[14][23] ), .B(\REGISTERS[30][23] ), .S(
        ADD_RD2[4]), .Z(n760) );
  MUX2_X1 U788 ( .A(\REGISTERS[6][23] ), .B(\REGISTERS[22][23] ), .S(
        ADD_RD2[4]), .Z(n761) );
  MUX2_X1 U789 ( .A(n761), .B(n760), .S(ADD_RD2[3]), .Z(n762) );
  MUX2_X1 U790 ( .A(\REGISTERS[10][23] ), .B(\REGISTERS[26][23] ), .S(
        ADD_RD2[4]), .Z(n763) );
  MUX2_X1 U791 ( .A(\REGISTERS[2][23] ), .B(\REGISTERS[18][23] ), .S(
        ADD_RD2[4]), .Z(n764) );
  MUX2_X1 U792 ( .A(n764), .B(n763), .S(ADD_RD2[3]), .Z(n765) );
  MUX2_X1 U793 ( .A(n765), .B(n762), .S(ADD_RD2[2]), .Z(n766) );
  MUX2_X1 U794 ( .A(n766), .B(n759), .S(ADD_RD2[0]), .Z(n767) );
  MUX2_X1 U795 ( .A(\REGISTERS[13][23] ), .B(\REGISTERS[29][23] ), .S(
        ADD_RD2[4]), .Z(n768) );
  MUX2_X1 U796 ( .A(\REGISTERS[5][23] ), .B(\REGISTERS[21][23] ), .S(
        ADD_RD2[4]), .Z(n769) );
  MUX2_X1 U797 ( .A(n769), .B(n768), .S(ADD_RD2[3]), .Z(n770) );
  MUX2_X1 U798 ( .A(\REGISTERS[9][23] ), .B(\REGISTERS[25][23] ), .S(
        ADD_RD2[4]), .Z(n771) );
  MUX2_X1 U799 ( .A(\REGISTERS[1][23] ), .B(\REGISTERS[17][23] ), .S(
        ADD_RD2[4]), .Z(n772) );
  MUX2_X1 U800 ( .A(n772), .B(n771), .S(ADD_RD2[3]), .Z(n773) );
  MUX2_X1 U801 ( .A(n773), .B(n770), .S(ADD_RD2[2]), .Z(n774) );
  MUX2_X1 U802 ( .A(\REGISTERS[12][23] ), .B(\REGISTERS[28][23] ), .S(
        ADD_RD2[4]), .Z(n775) );
  MUX2_X1 U803 ( .A(\REGISTERS[4][23] ), .B(\REGISTERS[20][23] ), .S(
        ADD_RD2[4]), .Z(n776) );
  MUX2_X1 U804 ( .A(n776), .B(n775), .S(ADD_RD2[3]), .Z(n777) );
  MUX2_X1 U805 ( .A(\REGISTERS[8][23] ), .B(\REGISTERS[24][23] ), .S(
        ADD_RD2[4]), .Z(n778) );
  MUX2_X1 U806 ( .A(\REGISTERS[0][23] ), .B(\REGISTERS[16][23] ), .S(
        ADD_RD2[4]), .Z(n779) );
  MUX2_X1 U807 ( .A(n779), .B(n778), .S(ADD_RD2[3]), .Z(n780) );
  MUX2_X1 U808 ( .A(n780), .B(n777), .S(ADD_RD2[2]), .Z(n781) );
  MUX2_X1 U809 ( .A(n781), .B(n774), .S(ADD_RD2[0]), .Z(n782) );
  MUX2_X1 U810 ( .A(n782), .B(n767), .S(ADD_RD2[1]), .Z(N435) );
  MUX2_X1 U811 ( .A(\REGISTERS[15][24] ), .B(\REGISTERS[31][24] ), .S(
        ADD_RD2[4]), .Z(n783) );
  MUX2_X1 U812 ( .A(\REGISTERS[7][24] ), .B(\REGISTERS[23][24] ), .S(
        ADD_RD2[4]), .Z(n784) );
  MUX2_X1 U813 ( .A(n784), .B(n783), .S(ADD_RD2[3]), .Z(n785) );
  MUX2_X1 U814 ( .A(\REGISTERS[11][24] ), .B(\REGISTERS[27][24] ), .S(
        ADD_RD2[4]), .Z(n786) );
  MUX2_X1 U815 ( .A(\REGISTERS[3][24] ), .B(\REGISTERS[19][24] ), .S(
        ADD_RD2[4]), .Z(n787) );
  MUX2_X1 U816 ( .A(n787), .B(n786), .S(ADD_RD2[3]), .Z(n788) );
  MUX2_X1 U817 ( .A(n788), .B(n785), .S(ADD_RD2[2]), .Z(n789) );
  MUX2_X1 U818 ( .A(\REGISTERS[14][24] ), .B(\REGISTERS[30][24] ), .S(
        ADD_RD2[4]), .Z(n790) );
  MUX2_X1 U819 ( .A(\REGISTERS[6][24] ), .B(\REGISTERS[22][24] ), .S(
        ADD_RD2[4]), .Z(n791) );
  MUX2_X1 U820 ( .A(n791), .B(n790), .S(ADD_RD2[3]), .Z(n792) );
  MUX2_X1 U821 ( .A(\REGISTERS[10][24] ), .B(\REGISTERS[26][24] ), .S(
        ADD_RD2[4]), .Z(n793) );
  MUX2_X1 U822 ( .A(\REGISTERS[2][24] ), .B(\REGISTERS[18][24] ), .S(
        ADD_RD2[4]), .Z(n794) );
  MUX2_X1 U823 ( .A(n794), .B(n793), .S(ADD_RD2[3]), .Z(n795) );
  MUX2_X1 U824 ( .A(n795), .B(n792), .S(ADD_RD2[2]), .Z(n796) );
  MUX2_X1 U825 ( .A(n796), .B(n789), .S(ADD_RD2[0]), .Z(n797) );
  MUX2_X1 U826 ( .A(\REGISTERS[13][24] ), .B(\REGISTERS[29][24] ), .S(
        ADD_RD2[4]), .Z(n798) );
  MUX2_X1 U827 ( .A(\REGISTERS[5][24] ), .B(\REGISTERS[21][24] ), .S(
        ADD_RD2[4]), .Z(n799) );
  MUX2_X1 U828 ( .A(n799), .B(n798), .S(ADD_RD2[3]), .Z(n800) );
  MUX2_X1 U829 ( .A(\REGISTERS[9][24] ), .B(\REGISTERS[25][24] ), .S(
        ADD_RD2[4]), .Z(n801) );
  MUX2_X1 U830 ( .A(\REGISTERS[1][24] ), .B(\REGISTERS[17][24] ), .S(
        ADD_RD2[4]), .Z(n802) );
  MUX2_X1 U831 ( .A(n802), .B(n801), .S(ADD_RD2[3]), .Z(n803) );
  MUX2_X1 U832 ( .A(n803), .B(n800), .S(ADD_RD2[2]), .Z(n804) );
  MUX2_X1 U833 ( .A(\REGISTERS[12][24] ), .B(\REGISTERS[28][24] ), .S(
        ADD_RD2[4]), .Z(n805) );
  MUX2_X1 U834 ( .A(\REGISTERS[4][24] ), .B(\REGISTERS[20][24] ), .S(
        ADD_RD2[4]), .Z(n806) );
  MUX2_X1 U835 ( .A(n806), .B(n805), .S(ADD_RD2[3]), .Z(n807) );
  MUX2_X1 U836 ( .A(\REGISTERS[8][24] ), .B(\REGISTERS[24][24] ), .S(
        ADD_RD2[4]), .Z(n808) );
  MUX2_X1 U837 ( .A(\REGISTERS[0][24] ), .B(\REGISTERS[16][24] ), .S(
        ADD_RD2[4]), .Z(n809) );
  MUX2_X1 U838 ( .A(n809), .B(n808), .S(ADD_RD2[3]), .Z(n810) );
  MUX2_X1 U839 ( .A(n810), .B(n807), .S(ADD_RD2[2]), .Z(n811) );
  MUX2_X1 U840 ( .A(n811), .B(n804), .S(ADD_RD2[0]), .Z(n812) );
  MUX2_X1 U841 ( .A(n812), .B(n797), .S(ADD_RD2[1]), .Z(N436) );
  MUX2_X1 U842 ( .A(\REGISTERS[15][25] ), .B(\REGISTERS[31][25] ), .S(
        ADD_RD2[4]), .Z(n813) );
  MUX2_X1 U843 ( .A(\REGISTERS[7][25] ), .B(\REGISTERS[23][25] ), .S(
        ADD_RD2[4]), .Z(n814) );
  MUX2_X1 U844 ( .A(n814), .B(n813), .S(ADD_RD2[3]), .Z(n815) );
  MUX2_X1 U845 ( .A(\REGISTERS[11][25] ), .B(\REGISTERS[27][25] ), .S(
        ADD_RD2[4]), .Z(n816) );
  MUX2_X1 U846 ( .A(\REGISTERS[3][25] ), .B(\REGISTERS[19][25] ), .S(
        ADD_RD2[4]), .Z(n817) );
  MUX2_X1 U847 ( .A(n817), .B(n816), .S(ADD_RD2[3]), .Z(n818) );
  MUX2_X1 U848 ( .A(n818), .B(n815), .S(ADD_RD2[2]), .Z(n819) );
  MUX2_X1 U849 ( .A(\REGISTERS[14][25] ), .B(\REGISTERS[30][25] ), .S(
        ADD_RD2[4]), .Z(n820) );
  MUX2_X1 U850 ( .A(\REGISTERS[6][25] ), .B(\REGISTERS[22][25] ), .S(
        ADD_RD2[4]), .Z(n821) );
  MUX2_X1 U851 ( .A(n821), .B(n820), .S(ADD_RD2[3]), .Z(n822) );
  MUX2_X1 U852 ( .A(\REGISTERS[10][25] ), .B(\REGISTERS[26][25] ), .S(
        ADD_RD2[4]), .Z(n823) );
  MUX2_X1 U853 ( .A(\REGISTERS[2][25] ), .B(\REGISTERS[18][25] ), .S(
        ADD_RD2[4]), .Z(n824) );
  MUX2_X1 U854 ( .A(n824), .B(n823), .S(ADD_RD2[3]), .Z(n825) );
  MUX2_X1 U855 ( .A(n825), .B(n822), .S(ADD_RD2[2]), .Z(n826) );
  MUX2_X1 U856 ( .A(n826), .B(n819), .S(ADD_RD2[0]), .Z(n827) );
  MUX2_X1 U857 ( .A(\REGISTERS[13][25] ), .B(\REGISTERS[29][25] ), .S(
        ADD_RD2[4]), .Z(n828) );
  MUX2_X1 U858 ( .A(\REGISTERS[5][25] ), .B(\REGISTERS[21][25] ), .S(
        ADD_RD2[4]), .Z(n829) );
  MUX2_X1 U859 ( .A(n829), .B(n828), .S(ADD_RD2[3]), .Z(n830) );
  MUX2_X1 U860 ( .A(\REGISTERS[9][25] ), .B(\REGISTERS[25][25] ), .S(
        ADD_RD2[4]), .Z(n831) );
  MUX2_X1 U861 ( .A(\REGISTERS[1][25] ), .B(\REGISTERS[17][25] ), .S(
        ADD_RD2[4]), .Z(n832) );
  MUX2_X1 U862 ( .A(n832), .B(n831), .S(ADD_RD2[3]), .Z(n833) );
  MUX2_X1 U863 ( .A(n833), .B(n830), .S(ADD_RD2[2]), .Z(n834) );
  MUX2_X1 U864 ( .A(\REGISTERS[12][25] ), .B(\REGISTERS[28][25] ), .S(
        ADD_RD2[4]), .Z(n835) );
  MUX2_X1 U865 ( .A(\REGISTERS[4][25] ), .B(\REGISTERS[20][25] ), .S(
        ADD_RD2[4]), .Z(n836) );
  MUX2_X1 U866 ( .A(n836), .B(n835), .S(ADD_RD2[3]), .Z(n837) );
  MUX2_X1 U867 ( .A(\REGISTERS[8][25] ), .B(\REGISTERS[24][25] ), .S(
        ADD_RD2[4]), .Z(n838) );
  MUX2_X1 U868 ( .A(\REGISTERS[0][25] ), .B(\REGISTERS[16][25] ), .S(
        ADD_RD2[4]), .Z(n839) );
  MUX2_X1 U869 ( .A(n839), .B(n838), .S(ADD_RD2[3]), .Z(n840) );
  MUX2_X1 U870 ( .A(n840), .B(n837), .S(ADD_RD2[2]), .Z(n841) );
  MUX2_X1 U871 ( .A(n841), .B(n834), .S(ADD_RD2[0]), .Z(n842) );
  MUX2_X1 U872 ( .A(n842), .B(n827), .S(ADD_RD2[1]), .Z(N437) );
  MUX2_X1 U873 ( .A(\REGISTERS[15][26] ), .B(\REGISTERS[31][26] ), .S(
        ADD_RD2[4]), .Z(n843) );
  MUX2_X1 U874 ( .A(\REGISTERS[7][26] ), .B(\REGISTERS[23][26] ), .S(
        ADD_RD2[4]), .Z(n844) );
  MUX2_X1 U875 ( .A(n844), .B(n843), .S(ADD_RD2[3]), .Z(n845) );
  MUX2_X1 U876 ( .A(\REGISTERS[11][26] ), .B(\REGISTERS[27][26] ), .S(
        ADD_RD2[4]), .Z(n846) );
  MUX2_X1 U877 ( .A(\REGISTERS[3][26] ), .B(\REGISTERS[19][26] ), .S(
        ADD_RD2[4]), .Z(n847) );
  MUX2_X1 U878 ( .A(n847), .B(n846), .S(ADD_RD2[3]), .Z(n848) );
  MUX2_X1 U879 ( .A(n848), .B(n845), .S(ADD_RD2[2]), .Z(n849) );
  MUX2_X1 U880 ( .A(\REGISTERS[14][26] ), .B(\REGISTERS[30][26] ), .S(
        ADD_RD2[4]), .Z(n850) );
  MUX2_X1 U881 ( .A(\REGISTERS[6][26] ), .B(\REGISTERS[22][26] ), .S(
        ADD_RD2[4]), .Z(n851) );
  MUX2_X1 U882 ( .A(n851), .B(n850), .S(ADD_RD2[3]), .Z(n852) );
  MUX2_X1 U883 ( .A(\REGISTERS[10][26] ), .B(\REGISTERS[26][26] ), .S(
        ADD_RD2[4]), .Z(n853) );
  MUX2_X1 U884 ( .A(\REGISTERS[2][26] ), .B(\REGISTERS[18][26] ), .S(
        ADD_RD2[4]), .Z(n854) );
  MUX2_X1 U885 ( .A(n854), .B(n853), .S(ADD_RD2[3]), .Z(n855) );
  MUX2_X1 U886 ( .A(n855), .B(n852), .S(ADD_RD2[2]), .Z(n856) );
  MUX2_X1 U887 ( .A(n856), .B(n849), .S(ADD_RD2[0]), .Z(n857) );
  MUX2_X1 U888 ( .A(\REGISTERS[13][26] ), .B(\REGISTERS[29][26] ), .S(
        ADD_RD2[4]), .Z(n858) );
  MUX2_X1 U889 ( .A(\REGISTERS[5][26] ), .B(\REGISTERS[21][26] ), .S(
        ADD_RD2[4]), .Z(n859) );
  MUX2_X1 U890 ( .A(n859), .B(n858), .S(ADD_RD2[3]), .Z(n860) );
  MUX2_X1 U891 ( .A(\REGISTERS[9][26] ), .B(\REGISTERS[25][26] ), .S(
        ADD_RD2[4]), .Z(n861) );
  MUX2_X1 U892 ( .A(\REGISTERS[1][26] ), .B(\REGISTERS[17][26] ), .S(
        ADD_RD2[4]), .Z(n862) );
  MUX2_X1 U893 ( .A(n862), .B(n861), .S(ADD_RD2[3]), .Z(n863) );
  MUX2_X1 U894 ( .A(n863), .B(n860), .S(ADD_RD2[2]), .Z(n864) );
  MUX2_X1 U895 ( .A(\REGISTERS[12][26] ), .B(\REGISTERS[28][26] ), .S(
        ADD_RD2[4]), .Z(n865) );
  MUX2_X1 U896 ( .A(\REGISTERS[4][26] ), .B(\REGISTERS[20][26] ), .S(
        ADD_RD2[4]), .Z(n866) );
  MUX2_X1 U897 ( .A(n866), .B(n865), .S(ADD_RD2[3]), .Z(n867) );
  MUX2_X1 U898 ( .A(\REGISTERS[8][26] ), .B(\REGISTERS[24][26] ), .S(
        ADD_RD2[4]), .Z(n868) );
  MUX2_X1 U899 ( .A(\REGISTERS[0][26] ), .B(\REGISTERS[16][26] ), .S(
        ADD_RD2[4]), .Z(n869) );
  MUX2_X1 U900 ( .A(n869), .B(n868), .S(ADD_RD2[3]), .Z(n870) );
  MUX2_X1 U901 ( .A(n870), .B(n867), .S(ADD_RD2[2]), .Z(n871) );
  MUX2_X1 U902 ( .A(n871), .B(n864), .S(ADD_RD2[0]), .Z(n872) );
  MUX2_X1 U903 ( .A(n872), .B(n857), .S(ADD_RD2[1]), .Z(N438) );
  MUX2_X1 U904 ( .A(\REGISTERS[15][27] ), .B(\REGISTERS[31][27] ), .S(
        ADD_RD2[4]), .Z(n873) );
  MUX2_X1 U905 ( .A(\REGISTERS[7][27] ), .B(\REGISTERS[23][27] ), .S(
        ADD_RD2[4]), .Z(n874) );
  MUX2_X1 U906 ( .A(n874), .B(n873), .S(ADD_RD2[3]), .Z(n875) );
  MUX2_X1 U907 ( .A(\REGISTERS[11][27] ), .B(\REGISTERS[27][27] ), .S(
        ADD_RD2[4]), .Z(n876) );
  MUX2_X1 U908 ( .A(\REGISTERS[3][27] ), .B(\REGISTERS[19][27] ), .S(
        ADD_RD2[4]), .Z(n877) );
  MUX2_X1 U909 ( .A(n877), .B(n876), .S(ADD_RD2[3]), .Z(n878) );
  MUX2_X1 U910 ( .A(n878), .B(n875), .S(ADD_RD2[2]), .Z(n879) );
  MUX2_X1 U911 ( .A(\REGISTERS[14][27] ), .B(\REGISTERS[30][27] ), .S(
        ADD_RD2[4]), .Z(n880) );
  MUX2_X1 U912 ( .A(\REGISTERS[6][27] ), .B(\REGISTERS[22][27] ), .S(
        ADD_RD2[4]), .Z(n881) );
  MUX2_X1 U913 ( .A(n881), .B(n880), .S(ADD_RD2[3]), .Z(n882) );
  MUX2_X1 U914 ( .A(\REGISTERS[10][27] ), .B(\REGISTERS[26][27] ), .S(
        ADD_RD2[4]), .Z(n883) );
  MUX2_X1 U915 ( .A(\REGISTERS[2][27] ), .B(\REGISTERS[18][27] ), .S(
        ADD_RD2[4]), .Z(n884) );
  MUX2_X1 U916 ( .A(n884), .B(n883), .S(ADD_RD2[3]), .Z(n885) );
  MUX2_X1 U917 ( .A(n885), .B(n882), .S(ADD_RD2[2]), .Z(n886) );
  MUX2_X1 U918 ( .A(n886), .B(n879), .S(ADD_RD2[0]), .Z(n887) );
  MUX2_X1 U919 ( .A(\REGISTERS[13][27] ), .B(\REGISTERS[29][27] ), .S(
        ADD_RD2[4]), .Z(n888) );
  MUX2_X1 U920 ( .A(\REGISTERS[5][27] ), .B(\REGISTERS[21][27] ), .S(
        ADD_RD2[4]), .Z(n889) );
  MUX2_X1 U921 ( .A(n889), .B(n888), .S(ADD_RD2[3]), .Z(n890) );
  MUX2_X1 U922 ( .A(\REGISTERS[9][27] ), .B(\REGISTERS[25][27] ), .S(
        ADD_RD2[4]), .Z(n891) );
  MUX2_X1 U923 ( .A(\REGISTERS[1][27] ), .B(\REGISTERS[17][27] ), .S(
        ADD_RD2[4]), .Z(n892) );
  MUX2_X1 U924 ( .A(n892), .B(n891), .S(ADD_RD2[3]), .Z(n893) );
  MUX2_X1 U925 ( .A(n893), .B(n890), .S(ADD_RD2[2]), .Z(n894) );
  MUX2_X1 U926 ( .A(\REGISTERS[12][27] ), .B(\REGISTERS[28][27] ), .S(
        ADD_RD2[4]), .Z(n895) );
  MUX2_X1 U927 ( .A(\REGISTERS[4][27] ), .B(\REGISTERS[20][27] ), .S(
        ADD_RD2[4]), .Z(n896) );
  MUX2_X1 U928 ( .A(n896), .B(n895), .S(ADD_RD2[3]), .Z(n897) );
  MUX2_X1 U929 ( .A(\REGISTERS[8][27] ), .B(\REGISTERS[24][27] ), .S(
        ADD_RD2[4]), .Z(n898) );
  MUX2_X1 U930 ( .A(\REGISTERS[0][27] ), .B(\REGISTERS[16][27] ), .S(
        ADD_RD2[4]), .Z(n899) );
  MUX2_X1 U931 ( .A(n899), .B(n898), .S(ADD_RD2[3]), .Z(n900) );
  MUX2_X1 U932 ( .A(n900), .B(n897), .S(ADD_RD2[2]), .Z(n901) );
  MUX2_X1 U933 ( .A(n901), .B(n894), .S(ADD_RD2[0]), .Z(n902) );
  MUX2_X1 U934 ( .A(n902), .B(n887), .S(ADD_RD2[1]), .Z(N439) );
  MUX2_X1 U935 ( .A(\REGISTERS[15][28] ), .B(\REGISTERS[31][28] ), .S(
        ADD_RD2[4]), .Z(n903) );
  MUX2_X1 U936 ( .A(\REGISTERS[7][28] ), .B(\REGISTERS[23][28] ), .S(
        ADD_RD2[4]), .Z(n904) );
  MUX2_X1 U937 ( .A(n904), .B(n903), .S(ADD_RD2[3]), .Z(n905) );
  MUX2_X1 U938 ( .A(\REGISTERS[11][28] ), .B(\REGISTERS[27][28] ), .S(
        ADD_RD2[4]), .Z(n906) );
  MUX2_X1 U939 ( .A(\REGISTERS[3][28] ), .B(\REGISTERS[19][28] ), .S(
        ADD_RD2[4]), .Z(n907) );
  MUX2_X1 U940 ( .A(n907), .B(n906), .S(ADD_RD2[3]), .Z(n908) );
  MUX2_X1 U941 ( .A(n908), .B(n905), .S(ADD_RD2[2]), .Z(n909) );
  MUX2_X1 U942 ( .A(\REGISTERS[14][28] ), .B(\REGISTERS[30][28] ), .S(
        ADD_RD2[4]), .Z(n910) );
  MUX2_X1 U943 ( .A(\REGISTERS[6][28] ), .B(\REGISTERS[22][28] ), .S(
        ADD_RD2[4]), .Z(n911) );
  MUX2_X1 U944 ( .A(n911), .B(n910), .S(ADD_RD2[3]), .Z(n912) );
  MUX2_X1 U945 ( .A(\REGISTERS[10][28] ), .B(\REGISTERS[26][28] ), .S(
        ADD_RD2[4]), .Z(n913) );
  MUX2_X1 U946 ( .A(\REGISTERS[2][28] ), .B(\REGISTERS[18][28] ), .S(
        ADD_RD2[4]), .Z(n914) );
  MUX2_X1 U947 ( .A(n914), .B(n913), .S(ADD_RD2[3]), .Z(n915) );
  MUX2_X1 U948 ( .A(n915), .B(n912), .S(ADD_RD2[2]), .Z(n916) );
  MUX2_X1 U949 ( .A(n916), .B(n909), .S(ADD_RD2[0]), .Z(n917) );
  MUX2_X1 U950 ( .A(\REGISTERS[13][28] ), .B(\REGISTERS[29][28] ), .S(
        ADD_RD2[4]), .Z(n918) );
  MUX2_X1 U951 ( .A(\REGISTERS[5][28] ), .B(\REGISTERS[21][28] ), .S(
        ADD_RD2[4]), .Z(n919) );
  MUX2_X1 U952 ( .A(n919), .B(n918), .S(ADD_RD2[3]), .Z(n920) );
  MUX2_X1 U953 ( .A(\REGISTERS[9][28] ), .B(\REGISTERS[25][28] ), .S(
        ADD_RD2[4]), .Z(n921) );
  MUX2_X1 U954 ( .A(\REGISTERS[1][28] ), .B(\REGISTERS[17][28] ), .S(
        ADD_RD2[4]), .Z(n922) );
  MUX2_X1 U955 ( .A(n922), .B(n921), .S(ADD_RD2[3]), .Z(n923) );
  MUX2_X1 U956 ( .A(n923), .B(n920), .S(ADD_RD2[2]), .Z(n924) );
  MUX2_X1 U957 ( .A(\REGISTERS[12][28] ), .B(\REGISTERS[28][28] ), .S(
        ADD_RD2[4]), .Z(n925) );
  MUX2_X1 U958 ( .A(\REGISTERS[4][28] ), .B(\REGISTERS[20][28] ), .S(
        ADD_RD2[4]), .Z(n926) );
  MUX2_X1 U959 ( .A(n926), .B(n925), .S(ADD_RD2[3]), .Z(n927) );
  MUX2_X1 U960 ( .A(\REGISTERS[8][28] ), .B(\REGISTERS[24][28] ), .S(
        ADD_RD2[4]), .Z(n928) );
  MUX2_X1 U961 ( .A(\REGISTERS[0][28] ), .B(\REGISTERS[16][28] ), .S(
        ADD_RD2[4]), .Z(n929) );
  MUX2_X1 U962 ( .A(n929), .B(n928), .S(ADD_RD2[3]), .Z(n930) );
  MUX2_X1 U963 ( .A(n930), .B(n927), .S(ADD_RD2[2]), .Z(n931) );
  MUX2_X1 U964 ( .A(n931), .B(n924), .S(ADD_RD2[0]), .Z(n932) );
  MUX2_X1 U965 ( .A(n932), .B(n917), .S(ADD_RD2[1]), .Z(N440) );
  MUX2_X1 U966 ( .A(\REGISTERS[15][29] ), .B(\REGISTERS[31][29] ), .S(
        ADD_RD2[4]), .Z(n933) );
  MUX2_X1 U967 ( .A(\REGISTERS[7][29] ), .B(\REGISTERS[23][29] ), .S(
        ADD_RD2[4]), .Z(n934) );
  MUX2_X1 U968 ( .A(n934), .B(n933), .S(ADD_RD2[3]), .Z(n935) );
  MUX2_X1 U969 ( .A(\REGISTERS[11][29] ), .B(\REGISTERS[27][29] ), .S(
        ADD_RD2[4]), .Z(n936) );
  MUX2_X1 U970 ( .A(\REGISTERS[3][29] ), .B(\REGISTERS[19][29] ), .S(
        ADD_RD2[4]), .Z(n937) );
  MUX2_X1 U971 ( .A(n937), .B(n936), .S(ADD_RD2[3]), .Z(n938) );
  MUX2_X1 U972 ( .A(n938), .B(n935), .S(ADD_RD2[2]), .Z(n939) );
  MUX2_X1 U973 ( .A(\REGISTERS[14][29] ), .B(\REGISTERS[30][29] ), .S(
        ADD_RD2[4]), .Z(n940) );
  MUX2_X1 U974 ( .A(\REGISTERS[6][29] ), .B(\REGISTERS[22][29] ), .S(
        ADD_RD2[4]), .Z(n941) );
  MUX2_X1 U975 ( .A(n941), .B(n940), .S(ADD_RD2[3]), .Z(n942) );
  MUX2_X1 U976 ( .A(\REGISTERS[10][29] ), .B(\REGISTERS[26][29] ), .S(
        ADD_RD2[4]), .Z(n943) );
  MUX2_X1 U977 ( .A(\REGISTERS[2][29] ), .B(\REGISTERS[18][29] ), .S(
        ADD_RD2[4]), .Z(n944) );
  MUX2_X1 U978 ( .A(n944), .B(n943), .S(ADD_RD2[3]), .Z(n945) );
  MUX2_X1 U979 ( .A(n945), .B(n942), .S(ADD_RD2[2]), .Z(n946) );
  MUX2_X1 U980 ( .A(n946), .B(n939), .S(ADD_RD2[0]), .Z(n947) );
  MUX2_X1 U981 ( .A(\REGISTERS[13][29] ), .B(\REGISTERS[29][29] ), .S(
        ADD_RD2[4]), .Z(n948) );
  MUX2_X1 U982 ( .A(\REGISTERS[5][29] ), .B(\REGISTERS[21][29] ), .S(
        ADD_RD2[4]), .Z(n949) );
  MUX2_X1 U983 ( .A(n949), .B(n948), .S(ADD_RD2[3]), .Z(n950) );
  MUX2_X1 U984 ( .A(\REGISTERS[9][29] ), .B(\REGISTERS[25][29] ), .S(
        ADD_RD2[4]), .Z(n951) );
  MUX2_X1 U985 ( .A(\REGISTERS[1][29] ), .B(\REGISTERS[17][29] ), .S(
        ADD_RD2[4]), .Z(n952) );
  MUX2_X1 U986 ( .A(n952), .B(n951), .S(ADD_RD2[3]), .Z(n953) );
  MUX2_X1 U987 ( .A(n953), .B(n950), .S(ADD_RD2[2]), .Z(n954) );
  MUX2_X1 U988 ( .A(\REGISTERS[12][29] ), .B(\REGISTERS[28][29] ), .S(
        ADD_RD2[4]), .Z(n955) );
  MUX2_X1 U989 ( .A(\REGISTERS[4][29] ), .B(\REGISTERS[20][29] ), .S(
        ADD_RD2[4]), .Z(n956) );
  MUX2_X1 U990 ( .A(n956), .B(n955), .S(ADD_RD2[3]), .Z(n957) );
  MUX2_X1 U991 ( .A(\REGISTERS[8][29] ), .B(\REGISTERS[24][29] ), .S(
        ADD_RD2[4]), .Z(n958) );
  MUX2_X1 U992 ( .A(\REGISTERS[0][29] ), .B(\REGISTERS[16][29] ), .S(
        ADD_RD2[4]), .Z(n959) );
  MUX2_X1 U993 ( .A(n959), .B(n958), .S(ADD_RD2[3]), .Z(n960) );
  MUX2_X1 U994 ( .A(n960), .B(n957), .S(ADD_RD2[2]), .Z(n961) );
  MUX2_X1 U995 ( .A(n961), .B(n954), .S(ADD_RD2[0]), .Z(n962) );
  MUX2_X1 U996 ( .A(n962), .B(n947), .S(ADD_RD2[1]), .Z(N441) );
  MUX2_X1 U997 ( .A(\REGISTERS[15][30] ), .B(\REGISTERS[31][30] ), .S(
        ADD_RD2[4]), .Z(n963) );
  MUX2_X1 U998 ( .A(\REGISTERS[7][30] ), .B(\REGISTERS[23][30] ), .S(
        ADD_RD2[4]), .Z(n964) );
  MUX2_X1 U999 ( .A(n964), .B(n963), .S(ADD_RD2[3]), .Z(n965) );
  MUX2_X1 U1000 ( .A(\REGISTERS[11][30] ), .B(\REGISTERS[27][30] ), .S(
        ADD_RD2[4]), .Z(n966) );
  MUX2_X1 U1001 ( .A(\REGISTERS[3][30] ), .B(\REGISTERS[19][30] ), .S(
        ADD_RD2[4]), .Z(n967) );
  MUX2_X1 U1002 ( .A(n967), .B(n966), .S(ADD_RD2[3]), .Z(n968) );
  MUX2_X1 U1003 ( .A(n968), .B(n965), .S(ADD_RD2[2]), .Z(n969) );
  MUX2_X1 U1004 ( .A(\REGISTERS[14][30] ), .B(\REGISTERS[30][30] ), .S(
        ADD_RD2[4]), .Z(n970) );
  MUX2_X1 U1005 ( .A(\REGISTERS[6][30] ), .B(\REGISTERS[22][30] ), .S(
        ADD_RD2[4]), .Z(n971) );
  MUX2_X1 U1006 ( .A(n971), .B(n970), .S(ADD_RD2[3]), .Z(n972) );
  MUX2_X1 U1007 ( .A(\REGISTERS[10][30] ), .B(\REGISTERS[26][30] ), .S(
        ADD_RD2[4]), .Z(n973) );
  MUX2_X1 U1008 ( .A(\REGISTERS[2][30] ), .B(\REGISTERS[18][30] ), .S(
        ADD_RD2[4]), .Z(n974) );
  MUX2_X1 U1009 ( .A(n974), .B(n973), .S(ADD_RD2[3]), .Z(n975) );
  MUX2_X1 U1010 ( .A(n975), .B(n972), .S(ADD_RD2[2]), .Z(n976) );
  MUX2_X1 U1011 ( .A(n976), .B(n969), .S(ADD_RD2[0]), .Z(n977) );
  MUX2_X1 U1012 ( .A(\REGISTERS[13][30] ), .B(\REGISTERS[29][30] ), .S(
        ADD_RD2[4]), .Z(n978) );
  MUX2_X1 U1013 ( .A(\REGISTERS[5][30] ), .B(\REGISTERS[21][30] ), .S(
        ADD_RD2[4]), .Z(n979) );
  MUX2_X1 U1014 ( .A(n979), .B(n978), .S(ADD_RD2[3]), .Z(n980) );
  MUX2_X1 U1015 ( .A(\REGISTERS[9][30] ), .B(\REGISTERS[25][30] ), .S(
        ADD_RD2[4]), .Z(n981) );
  MUX2_X1 U1016 ( .A(\REGISTERS[1][30] ), .B(\REGISTERS[17][30] ), .S(
        ADD_RD2[4]), .Z(n982) );
  MUX2_X1 U1017 ( .A(n982), .B(n981), .S(ADD_RD2[3]), .Z(n983) );
  MUX2_X1 U1018 ( .A(n983), .B(n980), .S(ADD_RD2[2]), .Z(n984) );
  MUX2_X1 U1019 ( .A(\REGISTERS[12][30] ), .B(\REGISTERS[28][30] ), .S(
        ADD_RD2[4]), .Z(n985) );
  MUX2_X1 U1020 ( .A(\REGISTERS[4][30] ), .B(\REGISTERS[20][30] ), .S(
        ADD_RD2[4]), .Z(n986) );
  MUX2_X1 U1021 ( .A(n986), .B(n985), .S(ADD_RD2[3]), .Z(n987) );
  MUX2_X1 U1022 ( .A(\REGISTERS[8][30] ), .B(\REGISTERS[24][30] ), .S(
        ADD_RD2[4]), .Z(n988) );
  MUX2_X1 U1023 ( .A(\REGISTERS[0][30] ), .B(\REGISTERS[16][30] ), .S(
        ADD_RD2[4]), .Z(n989) );
  MUX2_X1 U1024 ( .A(n989), .B(n988), .S(ADD_RD2[3]), .Z(n990) );
  MUX2_X1 U1025 ( .A(n990), .B(n987), .S(ADD_RD2[2]), .Z(n991) );
  MUX2_X1 U1026 ( .A(n991), .B(n984), .S(ADD_RD2[0]), .Z(n992) );
  MUX2_X1 U1027 ( .A(n992), .B(n977), .S(ADD_RD2[1]), .Z(N442) );
  MUX2_X1 U1028 ( .A(\REGISTERS[15][31] ), .B(\REGISTERS[31][31] ), .S(
        ADD_RD2[4]), .Z(n993) );
  MUX2_X1 U1029 ( .A(\REGISTERS[7][31] ), .B(\REGISTERS[23][31] ), .S(
        ADD_RD2[4]), .Z(n994) );
  MUX2_X1 U1030 ( .A(n994), .B(n993), .S(ADD_RD2[3]), .Z(n995) );
  MUX2_X1 U1031 ( .A(\REGISTERS[11][31] ), .B(\REGISTERS[27][31] ), .S(
        ADD_RD2[4]), .Z(n996) );
  MUX2_X1 U1032 ( .A(\REGISTERS[3][31] ), .B(\REGISTERS[19][31] ), .S(
        ADD_RD2[4]), .Z(n997) );
  MUX2_X1 U1033 ( .A(n997), .B(n996), .S(ADD_RD2[3]), .Z(n998) );
  MUX2_X1 U1034 ( .A(n998), .B(n995), .S(ADD_RD2[2]), .Z(n999) );
  MUX2_X1 U1035 ( .A(\REGISTERS[14][31] ), .B(\REGISTERS[30][31] ), .S(
        ADD_RD2[4]), .Z(n1000) );
  MUX2_X1 U1036 ( .A(\REGISTERS[6][31] ), .B(\REGISTERS[22][31] ), .S(
        ADD_RD2[4]), .Z(n1001) );
  MUX2_X1 U1037 ( .A(n1001), .B(n1000), .S(ADD_RD2[3]), .Z(n1002) );
  MUX2_X1 U1038 ( .A(\REGISTERS[10][31] ), .B(\REGISTERS[26][31] ), .S(
        ADD_RD2[4]), .Z(n1003) );
  MUX2_X1 U1039 ( .A(\REGISTERS[2][31] ), .B(\REGISTERS[18][31] ), .S(
        ADD_RD2[4]), .Z(n1004) );
  MUX2_X1 U1040 ( .A(n1004), .B(n1003), .S(ADD_RD2[3]), .Z(n1005) );
  MUX2_X1 U1041 ( .A(n1005), .B(n1002), .S(ADD_RD2[2]), .Z(n1006) );
  MUX2_X1 U1042 ( .A(n1006), .B(n999), .S(ADD_RD2[0]), .Z(n1007) );
  MUX2_X1 U1043 ( .A(\REGISTERS[13][31] ), .B(\REGISTERS[29][31] ), .S(
        ADD_RD2[4]), .Z(n1008) );
  MUX2_X1 U1044 ( .A(\REGISTERS[5][31] ), .B(\REGISTERS[21][31] ), .S(
        ADD_RD2[4]), .Z(n1009) );
  MUX2_X1 U1045 ( .A(n1009), .B(n1008), .S(ADD_RD2[3]), .Z(n1010) );
  MUX2_X1 U1046 ( .A(\REGISTERS[9][31] ), .B(\REGISTERS[25][31] ), .S(
        ADD_RD2[4]), .Z(n1011) );
  MUX2_X1 U1047 ( .A(\REGISTERS[1][31] ), .B(\REGISTERS[17][31] ), .S(
        ADD_RD2[4]), .Z(n1012) );
  MUX2_X1 U1048 ( .A(n1012), .B(n1011), .S(ADD_RD2[3]), .Z(n1013) );
  MUX2_X1 U1049 ( .A(n1013), .B(n1010), .S(ADD_RD2[2]), .Z(n1014) );
  MUX2_X1 U1050 ( .A(\REGISTERS[12][31] ), .B(\REGISTERS[28][31] ), .S(
        ADD_RD2[4]), .Z(n1015) );
  MUX2_X1 U1051 ( .A(\REGISTERS[4][31] ), .B(\REGISTERS[20][31] ), .S(
        ADD_RD2[4]), .Z(n1016) );
  MUX2_X1 U1052 ( .A(n1016), .B(n1015), .S(ADD_RD2[3]), .Z(n1017) );
  MUX2_X1 U1053 ( .A(\REGISTERS[8][31] ), .B(\REGISTERS[24][31] ), .S(
        ADD_RD2[4]), .Z(n1018) );
  MUX2_X1 U1054 ( .A(\REGISTERS[0][31] ), .B(\REGISTERS[16][31] ), .S(
        ADD_RD2[4]), .Z(n1019) );
  MUX2_X1 U1055 ( .A(n1019), .B(n1018), .S(ADD_RD2[3]), .Z(n1020) );
  MUX2_X1 U1056 ( .A(n1020), .B(n1017), .S(ADD_RD2[2]), .Z(n1021) );
  MUX2_X1 U1057 ( .A(n1021), .B(n1014), .S(ADD_RD2[0]), .Z(n1022) );
  MUX2_X1 U1058 ( .A(n1022), .B(n1007), .S(ADD_RD2[1]), .Z(N443) );
  MUX2_X1 U1059 ( .A(\REGISTERS[15][0] ), .B(\REGISTERS[31][0] ), .S(
        ADD_RD1[4]), .Z(n1023) );
  MUX2_X1 U1060 ( .A(\REGISTERS[7][0] ), .B(\REGISTERS[23][0] ), .S(ADD_RD1[4]), .Z(n1024) );
  MUX2_X1 U1061 ( .A(n1024), .B(n1023), .S(ADD_RD1[3]), .Z(n1025) );
  MUX2_X1 U1062 ( .A(\REGISTERS[11][0] ), .B(\REGISTERS[27][0] ), .S(
        ADD_RD1[4]), .Z(n1026) );
  MUX2_X1 U1063 ( .A(\REGISTERS[3][0] ), .B(\REGISTERS[19][0] ), .S(ADD_RD1[4]), .Z(n1027) );
  MUX2_X1 U1064 ( .A(n1027), .B(n1026), .S(ADD_RD1[3]), .Z(n1028) );
  MUX2_X1 U1065 ( .A(n1028), .B(n1025), .S(ADD_RD1[2]), .Z(n1029) );
  MUX2_X1 U1066 ( .A(\REGISTERS[14][0] ), .B(\REGISTERS[30][0] ), .S(
        ADD_RD1[4]), .Z(n1030) );
  MUX2_X1 U1067 ( .A(\REGISTERS[6][0] ), .B(\REGISTERS[22][0] ), .S(ADD_RD1[4]), .Z(n1031) );
  MUX2_X1 U1068 ( .A(n1031), .B(n1030), .S(ADD_RD1[3]), .Z(n1032) );
  MUX2_X1 U1069 ( .A(\REGISTERS[10][0] ), .B(\REGISTERS[26][0] ), .S(
        ADD_RD1[4]), .Z(n1033) );
  MUX2_X1 U1070 ( .A(\REGISTERS[2][0] ), .B(\REGISTERS[18][0] ), .S(ADD_RD1[4]), .Z(n1034) );
  MUX2_X1 U1071 ( .A(n1034), .B(n1033), .S(ADD_RD1[3]), .Z(n1035) );
  MUX2_X1 U1072 ( .A(n1035), .B(n1032), .S(ADD_RD1[2]), .Z(n1036) );
  MUX2_X1 U1073 ( .A(n1036), .B(n1029), .S(ADD_RD1[0]), .Z(n1037) );
  MUX2_X1 U1074 ( .A(\REGISTERS[13][0] ), .B(\REGISTERS[29][0] ), .S(
        ADD_RD1[4]), .Z(n1038) );
  MUX2_X1 U1075 ( .A(\REGISTERS[5][0] ), .B(\REGISTERS[21][0] ), .S(ADD_RD1[4]), .Z(n1039) );
  MUX2_X1 U1076 ( .A(n1039), .B(n1038), .S(ADD_RD1[3]), .Z(n1040) );
  MUX2_X1 U1077 ( .A(\REGISTERS[9][0] ), .B(\REGISTERS[25][0] ), .S(ADD_RD1[4]), .Z(n1041) );
  MUX2_X1 U1078 ( .A(\REGISTERS[1][0] ), .B(\REGISTERS[17][0] ), .S(ADD_RD1[4]), .Z(n1042) );
  MUX2_X1 U1079 ( .A(n1042), .B(n1041), .S(ADD_RD1[3]), .Z(n1043) );
  MUX2_X1 U1080 ( .A(n1043), .B(n1040), .S(ADD_RD1[2]), .Z(n1044) );
  MUX2_X1 U1081 ( .A(\REGISTERS[12][0] ), .B(\REGISTERS[28][0] ), .S(
        ADD_RD1[4]), .Z(n1045) );
  MUX2_X1 U1082 ( .A(\REGISTERS[4][0] ), .B(\REGISTERS[20][0] ), .S(ADD_RD1[4]), .Z(n1046) );
  MUX2_X1 U1083 ( .A(n1046), .B(n1045), .S(ADD_RD1[3]), .Z(n1047) );
  MUX2_X1 U1084 ( .A(\REGISTERS[8][0] ), .B(\REGISTERS[24][0] ), .S(ADD_RD1[4]), .Z(n1048) );
  MUX2_X1 U1085 ( .A(\REGISTERS[0][0] ), .B(\REGISTERS[16][0] ), .S(ADD_RD1[4]), .Z(n1049) );
  MUX2_X1 U1086 ( .A(n1049), .B(n1048), .S(ADD_RD1[3]), .Z(n1050) );
  MUX2_X1 U1087 ( .A(n1050), .B(n1047), .S(ADD_RD1[2]), .Z(n1051) );
  MUX2_X1 U1088 ( .A(n1051), .B(n1044), .S(ADD_RD1[0]), .Z(n1052) );
  MUX2_X1 U1089 ( .A(n1052), .B(n1037), .S(ADD_RD1[1]), .Z(N379) );
  MUX2_X1 U1090 ( .A(\REGISTERS[15][1] ), .B(\REGISTERS[31][1] ), .S(
        ADD_RD1[4]), .Z(n1053) );
  MUX2_X1 U1091 ( .A(\REGISTERS[7][1] ), .B(\REGISTERS[23][1] ), .S(ADD_RD1[4]), .Z(n1054) );
  MUX2_X1 U1092 ( .A(n1054), .B(n1053), .S(ADD_RD1[3]), .Z(n1055) );
  MUX2_X1 U1093 ( .A(\REGISTERS[11][1] ), .B(\REGISTERS[27][1] ), .S(
        ADD_RD1[4]), .Z(n1056) );
  MUX2_X1 U1094 ( .A(\REGISTERS[3][1] ), .B(\REGISTERS[19][1] ), .S(ADD_RD1[4]), .Z(n1057) );
  MUX2_X1 U1095 ( .A(n1057), .B(n1056), .S(ADD_RD1[3]), .Z(n1058) );
  MUX2_X1 U1096 ( .A(n1058), .B(n1055), .S(ADD_RD1[2]), .Z(n1059) );
  MUX2_X1 U1097 ( .A(\REGISTERS[14][1] ), .B(\REGISTERS[30][1] ), .S(
        ADD_RD1[4]), .Z(n1060) );
  MUX2_X1 U1098 ( .A(\REGISTERS[6][1] ), .B(\REGISTERS[22][1] ), .S(ADD_RD1[4]), .Z(n1061) );
  MUX2_X1 U1099 ( .A(n1061), .B(n1060), .S(ADD_RD1[3]), .Z(n1062) );
  MUX2_X1 U1100 ( .A(\REGISTERS[10][1] ), .B(\REGISTERS[26][1] ), .S(
        ADD_RD1[4]), .Z(n1063) );
  MUX2_X1 U1101 ( .A(\REGISTERS[2][1] ), .B(\REGISTERS[18][1] ), .S(ADD_RD1[4]), .Z(n1064) );
  MUX2_X1 U1102 ( .A(n1064), .B(n1063), .S(ADD_RD1[3]), .Z(n1065) );
  MUX2_X1 U1103 ( .A(n1065), .B(n1062), .S(ADD_RD1[2]), .Z(n1066) );
  MUX2_X1 U1104 ( .A(n1066), .B(n1059), .S(ADD_RD1[0]), .Z(n1067) );
  MUX2_X1 U1105 ( .A(\REGISTERS[13][1] ), .B(\REGISTERS[29][1] ), .S(
        ADD_RD1[4]), .Z(n1068) );
  MUX2_X1 U1106 ( .A(\REGISTERS[5][1] ), .B(\REGISTERS[21][1] ), .S(ADD_RD1[4]), .Z(n1069) );
  MUX2_X1 U1107 ( .A(n1069), .B(n1068), .S(ADD_RD1[3]), .Z(n1070) );
  MUX2_X1 U1108 ( .A(\REGISTERS[9][1] ), .B(\REGISTERS[25][1] ), .S(ADD_RD1[4]), .Z(n1071) );
  MUX2_X1 U1109 ( .A(\REGISTERS[1][1] ), .B(\REGISTERS[17][1] ), .S(ADD_RD1[4]), .Z(n1072) );
  MUX2_X1 U1110 ( .A(n1072), .B(n1071), .S(ADD_RD1[3]), .Z(n1073) );
  MUX2_X1 U1111 ( .A(n1073), .B(n1070), .S(ADD_RD1[2]), .Z(n1074) );
  MUX2_X1 U1112 ( .A(\REGISTERS[12][1] ), .B(\REGISTERS[28][1] ), .S(
        ADD_RD1[4]), .Z(n1075) );
  MUX2_X1 U1113 ( .A(\REGISTERS[4][1] ), .B(\REGISTERS[20][1] ), .S(ADD_RD1[4]), .Z(n1076) );
  MUX2_X1 U1114 ( .A(n1076), .B(n1075), .S(ADD_RD1[3]), .Z(n1077) );
  MUX2_X1 U1115 ( .A(\REGISTERS[8][1] ), .B(\REGISTERS[24][1] ), .S(ADD_RD1[4]), .Z(n1078) );
  MUX2_X1 U1116 ( .A(\REGISTERS[0][1] ), .B(\REGISTERS[16][1] ), .S(ADD_RD1[4]), .Z(n1079) );
  MUX2_X1 U1117 ( .A(n1079), .B(n1078), .S(ADD_RD1[3]), .Z(n1080) );
  MUX2_X1 U1118 ( .A(n1080), .B(n1077), .S(ADD_RD1[2]), .Z(n1081) );
  MUX2_X1 U1119 ( .A(n1081), .B(n1074), .S(ADD_RD1[0]), .Z(n1082) );
  MUX2_X1 U1120 ( .A(n1082), .B(n1067), .S(ADD_RD1[1]), .Z(N380) );
  MUX2_X1 U1121 ( .A(\REGISTERS[15][2] ), .B(\REGISTERS[31][2] ), .S(
        ADD_RD1[4]), .Z(n1083) );
  MUX2_X1 U1122 ( .A(\REGISTERS[7][2] ), .B(\REGISTERS[23][2] ), .S(ADD_RD1[4]), .Z(n1084) );
  MUX2_X1 U1123 ( .A(n1084), .B(n1083), .S(ADD_RD1[3]), .Z(n1085) );
  MUX2_X1 U1124 ( .A(\REGISTERS[11][2] ), .B(\REGISTERS[27][2] ), .S(
        ADD_RD1[4]), .Z(n1086) );
  MUX2_X1 U1125 ( .A(\REGISTERS[3][2] ), .B(\REGISTERS[19][2] ), .S(ADD_RD1[4]), .Z(n1087) );
  MUX2_X1 U1126 ( .A(n1087), .B(n1086), .S(ADD_RD1[3]), .Z(n1088) );
  MUX2_X1 U1127 ( .A(n1088), .B(n1085), .S(ADD_RD1[2]), .Z(n1089) );
  MUX2_X1 U1128 ( .A(\REGISTERS[14][2] ), .B(\REGISTERS[30][2] ), .S(
        ADD_RD1[4]), .Z(n1090) );
  MUX2_X1 U1129 ( .A(\REGISTERS[6][2] ), .B(\REGISTERS[22][2] ), .S(ADD_RD1[4]), .Z(n1091) );
  MUX2_X1 U1130 ( .A(n1091), .B(n1090), .S(ADD_RD1[3]), .Z(n1092) );
  MUX2_X1 U1131 ( .A(\REGISTERS[10][2] ), .B(\REGISTERS[26][2] ), .S(
        ADD_RD1[4]), .Z(n1093) );
  MUX2_X1 U1132 ( .A(\REGISTERS[2][2] ), .B(\REGISTERS[18][2] ), .S(ADD_RD1[4]), .Z(n1094) );
  MUX2_X1 U1133 ( .A(n1094), .B(n1093), .S(ADD_RD1[3]), .Z(n1095) );
  MUX2_X1 U1134 ( .A(n1095), .B(n1092), .S(ADD_RD1[2]), .Z(n1096) );
  MUX2_X1 U1135 ( .A(n1096), .B(n1089), .S(ADD_RD1[0]), .Z(n1097) );
  MUX2_X1 U1136 ( .A(\REGISTERS[13][2] ), .B(\REGISTERS[29][2] ), .S(
        ADD_RD1[4]), .Z(n1098) );
  MUX2_X1 U1137 ( .A(\REGISTERS[5][2] ), .B(\REGISTERS[21][2] ), .S(ADD_RD1[4]), .Z(n1099) );
  MUX2_X1 U1138 ( .A(n1099), .B(n1098), .S(ADD_RD1[3]), .Z(n1100) );
  MUX2_X1 U1139 ( .A(\REGISTERS[9][2] ), .B(\REGISTERS[25][2] ), .S(ADD_RD1[4]), .Z(n1101) );
  MUX2_X1 U1140 ( .A(\REGISTERS[1][2] ), .B(\REGISTERS[17][2] ), .S(ADD_RD1[4]), .Z(n1102) );
  MUX2_X1 U1141 ( .A(n1102), .B(n1101), .S(ADD_RD1[3]), .Z(n1103) );
  MUX2_X1 U1142 ( .A(n1103), .B(n1100), .S(ADD_RD1[2]), .Z(n1104) );
  MUX2_X1 U1143 ( .A(\REGISTERS[12][2] ), .B(\REGISTERS[28][2] ), .S(
        ADD_RD1[4]), .Z(n1105) );
  MUX2_X1 U1144 ( .A(\REGISTERS[4][2] ), .B(\REGISTERS[20][2] ), .S(ADD_RD1[4]), .Z(n1106) );
  MUX2_X1 U1145 ( .A(n1106), .B(n1105), .S(ADD_RD1[3]), .Z(n1107) );
  MUX2_X1 U1146 ( .A(\REGISTERS[8][2] ), .B(\REGISTERS[24][2] ), .S(ADD_RD1[4]), .Z(n1108) );
  MUX2_X1 U1147 ( .A(\REGISTERS[0][2] ), .B(\REGISTERS[16][2] ), .S(ADD_RD1[4]), .Z(n1109) );
  MUX2_X1 U1148 ( .A(n1109), .B(n1108), .S(ADD_RD1[3]), .Z(n1110) );
  MUX2_X1 U1149 ( .A(n1110), .B(n1107), .S(ADD_RD1[2]), .Z(n1111) );
  MUX2_X1 U1150 ( .A(n1111), .B(n1104), .S(ADD_RD1[0]), .Z(n1112) );
  MUX2_X1 U1151 ( .A(n1112), .B(n1097), .S(ADD_RD1[1]), .Z(N381) );
  MUX2_X1 U1152 ( .A(\REGISTERS[15][3] ), .B(\REGISTERS[31][3] ), .S(
        ADD_RD1[4]), .Z(n1113) );
  MUX2_X1 U1153 ( .A(\REGISTERS[7][3] ), .B(\REGISTERS[23][3] ), .S(ADD_RD1[4]), .Z(n1114) );
  MUX2_X1 U1154 ( .A(n1114), .B(n1113), .S(ADD_RD1[3]), .Z(n1115) );
  MUX2_X1 U1155 ( .A(\REGISTERS[11][3] ), .B(\REGISTERS[27][3] ), .S(
        ADD_RD1[4]), .Z(n1116) );
  MUX2_X1 U1156 ( .A(\REGISTERS[3][3] ), .B(\REGISTERS[19][3] ), .S(ADD_RD1[4]), .Z(n1117) );
  MUX2_X1 U1157 ( .A(n1117), .B(n1116), .S(ADD_RD1[3]), .Z(n1118) );
  MUX2_X1 U1158 ( .A(n1118), .B(n1115), .S(ADD_RD1[2]), .Z(n1119) );
  MUX2_X1 U1159 ( .A(\REGISTERS[14][3] ), .B(\REGISTERS[30][3] ), .S(
        ADD_RD1[4]), .Z(n1120) );
  MUX2_X1 U1160 ( .A(\REGISTERS[6][3] ), .B(\REGISTERS[22][3] ), .S(ADD_RD1[4]), .Z(n1121) );
  MUX2_X1 U1161 ( .A(n1121), .B(n1120), .S(ADD_RD1[3]), .Z(n1122) );
  MUX2_X1 U1162 ( .A(\REGISTERS[10][3] ), .B(\REGISTERS[26][3] ), .S(
        ADD_RD1[4]), .Z(n1123) );
  MUX2_X1 U1163 ( .A(\REGISTERS[2][3] ), .B(\REGISTERS[18][3] ), .S(ADD_RD1[4]), .Z(n1124) );
  MUX2_X1 U1164 ( .A(n1124), .B(n1123), .S(ADD_RD1[3]), .Z(n1125) );
  MUX2_X1 U1165 ( .A(n1125), .B(n1122), .S(ADD_RD1[2]), .Z(n1126) );
  MUX2_X1 U1166 ( .A(n1126), .B(n1119), .S(ADD_RD1[0]), .Z(n1127) );
  MUX2_X1 U1167 ( .A(\REGISTERS[13][3] ), .B(\REGISTERS[29][3] ), .S(
        ADD_RD1[4]), .Z(n1128) );
  MUX2_X1 U1168 ( .A(\REGISTERS[5][3] ), .B(\REGISTERS[21][3] ), .S(ADD_RD1[4]), .Z(n1129) );
  MUX2_X1 U1169 ( .A(n1129), .B(n1128), .S(ADD_RD1[3]), .Z(n1130) );
  MUX2_X1 U1170 ( .A(\REGISTERS[9][3] ), .B(\REGISTERS[25][3] ), .S(ADD_RD1[4]), .Z(n1131) );
  MUX2_X1 U1171 ( .A(\REGISTERS[1][3] ), .B(\REGISTERS[17][3] ), .S(ADD_RD1[4]), .Z(n1132) );
  MUX2_X1 U1172 ( .A(n1132), .B(n1131), .S(ADD_RD1[3]), .Z(n1133) );
  MUX2_X1 U1173 ( .A(n1133), .B(n1130), .S(ADD_RD1[2]), .Z(n1134) );
  MUX2_X1 U1174 ( .A(\REGISTERS[12][3] ), .B(\REGISTERS[28][3] ), .S(
        ADD_RD1[4]), .Z(n1135) );
  MUX2_X1 U1175 ( .A(\REGISTERS[4][3] ), .B(\REGISTERS[20][3] ), .S(ADD_RD1[4]), .Z(n1136) );
  MUX2_X1 U1176 ( .A(n1136), .B(n1135), .S(ADD_RD1[3]), .Z(n1137) );
  MUX2_X1 U1177 ( .A(\REGISTERS[8][3] ), .B(\REGISTERS[24][3] ), .S(ADD_RD1[4]), .Z(n1138) );
  MUX2_X1 U1178 ( .A(\REGISTERS[0][3] ), .B(\REGISTERS[16][3] ), .S(ADD_RD1[4]), .Z(n1139) );
  MUX2_X1 U1179 ( .A(n1139), .B(n1138), .S(ADD_RD1[3]), .Z(n2164) );
  MUX2_X1 U1180 ( .A(n2164), .B(n1137), .S(ADD_RD1[2]), .Z(n2165) );
  MUX2_X1 U1181 ( .A(n2165), .B(n1134), .S(ADD_RD1[0]), .Z(n2166) );
  MUX2_X1 U1182 ( .A(n2166), .B(n1127), .S(ADD_RD1[1]), .Z(N382) );
  MUX2_X1 U1183 ( .A(\REGISTERS[15][4] ), .B(\REGISTERS[31][4] ), .S(
        ADD_RD1[4]), .Z(n2167) );
  MUX2_X1 U1184 ( .A(\REGISTERS[7][4] ), .B(\REGISTERS[23][4] ), .S(ADD_RD1[4]), .Z(n2168) );
  MUX2_X1 U1185 ( .A(n2168), .B(n2167), .S(ADD_RD1[3]), .Z(n2169) );
  MUX2_X1 U1186 ( .A(\REGISTERS[11][4] ), .B(\REGISTERS[27][4] ), .S(
        ADD_RD1[4]), .Z(n2170) );
  MUX2_X1 U1187 ( .A(\REGISTERS[3][4] ), .B(\REGISTERS[19][4] ), .S(ADD_RD1[4]), .Z(n2171) );
  MUX2_X1 U1188 ( .A(n2171), .B(n2170), .S(ADD_RD1[3]), .Z(n2172) );
  MUX2_X1 U1189 ( .A(n2172), .B(n2169), .S(ADD_RD1[2]), .Z(n2173) );
  MUX2_X1 U1190 ( .A(\REGISTERS[14][4] ), .B(\REGISTERS[30][4] ), .S(
        ADD_RD1[4]), .Z(n2174) );
  MUX2_X1 U1191 ( .A(\REGISTERS[6][4] ), .B(\REGISTERS[22][4] ), .S(ADD_RD1[4]), .Z(n2175) );
  MUX2_X1 U1192 ( .A(n2175), .B(n2174), .S(ADD_RD1[3]), .Z(n2176) );
  MUX2_X1 U1193 ( .A(\REGISTERS[10][4] ), .B(\REGISTERS[26][4] ), .S(
        ADD_RD1[4]), .Z(n2177) );
  MUX2_X1 U1194 ( .A(\REGISTERS[2][4] ), .B(\REGISTERS[18][4] ), .S(ADD_RD1[4]), .Z(n2178) );
  MUX2_X1 U1195 ( .A(n2178), .B(n2177), .S(ADD_RD1[3]), .Z(n2179) );
  MUX2_X1 U1196 ( .A(n2179), .B(n2176), .S(ADD_RD1[2]), .Z(n2180) );
  MUX2_X1 U1197 ( .A(n2180), .B(n2173), .S(ADD_RD1[0]), .Z(n2181) );
  MUX2_X1 U1198 ( .A(\REGISTERS[13][4] ), .B(\REGISTERS[29][4] ), .S(
        ADD_RD1[4]), .Z(n2182) );
  MUX2_X1 U1199 ( .A(\REGISTERS[5][4] ), .B(\REGISTERS[21][4] ), .S(ADD_RD1[4]), .Z(n2183) );
  MUX2_X1 U1200 ( .A(n2183), .B(n2182), .S(ADD_RD1[3]), .Z(n2184) );
  MUX2_X1 U1201 ( .A(\REGISTERS[9][4] ), .B(\REGISTERS[25][4] ), .S(ADD_RD1[4]), .Z(n2185) );
  MUX2_X1 U1202 ( .A(\REGISTERS[1][4] ), .B(\REGISTERS[17][4] ), .S(ADD_RD1[4]), .Z(n2186) );
  MUX2_X1 U1203 ( .A(n2186), .B(n2185), .S(ADD_RD1[3]), .Z(n2187) );
  MUX2_X1 U1204 ( .A(n2187), .B(n2184), .S(ADD_RD1[2]), .Z(n2188) );
  MUX2_X1 U1205 ( .A(\REGISTERS[12][4] ), .B(\REGISTERS[28][4] ), .S(
        ADD_RD1[4]), .Z(n2189) );
  MUX2_X1 U1206 ( .A(\REGISTERS[4][4] ), .B(\REGISTERS[20][4] ), .S(ADD_RD1[4]), .Z(n2190) );
  MUX2_X1 U1207 ( .A(n2190), .B(n2189), .S(ADD_RD1[3]), .Z(n2191) );
  MUX2_X1 U1208 ( .A(\REGISTERS[8][4] ), .B(\REGISTERS[24][4] ), .S(ADD_RD1[4]), .Z(n2192) );
  MUX2_X1 U1209 ( .A(\REGISTERS[0][4] ), .B(\REGISTERS[16][4] ), .S(ADD_RD1[4]), .Z(n2193) );
  MUX2_X1 U1210 ( .A(n2193), .B(n2192), .S(ADD_RD1[3]), .Z(n2194) );
  MUX2_X1 U1211 ( .A(n2194), .B(n2191), .S(ADD_RD1[2]), .Z(n2195) );
  MUX2_X1 U1212 ( .A(n2195), .B(n2188), .S(ADD_RD1[0]), .Z(n2196) );
  MUX2_X1 U1213 ( .A(n2196), .B(n2181), .S(ADD_RD1[1]), .Z(N383) );
  MUX2_X1 U1214 ( .A(\REGISTERS[15][5] ), .B(\REGISTERS[31][5] ), .S(
        ADD_RD1[4]), .Z(n2197) );
  MUX2_X1 U1215 ( .A(\REGISTERS[7][5] ), .B(\REGISTERS[23][5] ), .S(ADD_RD1[4]), .Z(n2198) );
  MUX2_X1 U1216 ( .A(n2198), .B(n2197), .S(ADD_RD1[3]), .Z(n2199) );
  MUX2_X1 U1217 ( .A(\REGISTERS[11][5] ), .B(\REGISTERS[27][5] ), .S(
        ADD_RD1[4]), .Z(n2200) );
  MUX2_X1 U1218 ( .A(\REGISTERS[3][5] ), .B(\REGISTERS[19][5] ), .S(ADD_RD1[4]), .Z(n2201) );
  MUX2_X1 U1219 ( .A(n2201), .B(n2200), .S(ADD_RD1[3]), .Z(n2202) );
  MUX2_X1 U1220 ( .A(n2202), .B(n2199), .S(ADD_RD1[2]), .Z(n2203) );
  MUX2_X1 U1221 ( .A(\REGISTERS[14][5] ), .B(\REGISTERS[30][5] ), .S(
        ADD_RD1[4]), .Z(n2204) );
  MUX2_X1 U1222 ( .A(\REGISTERS[6][5] ), .B(\REGISTERS[22][5] ), .S(ADD_RD1[4]), .Z(n2205) );
  MUX2_X1 U1223 ( .A(n2205), .B(n2204), .S(ADD_RD1[3]), .Z(n2206) );
  MUX2_X1 U1224 ( .A(\REGISTERS[10][5] ), .B(\REGISTERS[26][5] ), .S(
        ADD_RD1[4]), .Z(n2207) );
  MUX2_X1 U1225 ( .A(\REGISTERS[2][5] ), .B(\REGISTERS[18][5] ), .S(ADD_RD1[4]), .Z(n2208) );
  MUX2_X1 U1226 ( .A(n2208), .B(n2207), .S(ADD_RD1[3]), .Z(n2209) );
  MUX2_X1 U1227 ( .A(n2209), .B(n2206), .S(ADD_RD1[2]), .Z(n2210) );
  MUX2_X1 U1228 ( .A(n2210), .B(n2203), .S(ADD_RD1[0]), .Z(n2211) );
  MUX2_X1 U1229 ( .A(\REGISTERS[13][5] ), .B(\REGISTERS[29][5] ), .S(
        ADD_RD1[4]), .Z(n2212) );
  MUX2_X1 U1230 ( .A(\REGISTERS[5][5] ), .B(\REGISTERS[21][5] ), .S(ADD_RD1[4]), .Z(n2213) );
  MUX2_X1 U1231 ( .A(n2213), .B(n2212), .S(ADD_RD1[3]), .Z(n2214) );
  MUX2_X1 U1232 ( .A(\REGISTERS[9][5] ), .B(\REGISTERS[25][5] ), .S(ADD_RD1[4]), .Z(n2215) );
  MUX2_X1 U1233 ( .A(\REGISTERS[1][5] ), .B(\REGISTERS[17][5] ), .S(ADD_RD1[4]), .Z(n2216) );
  MUX2_X1 U1234 ( .A(n2216), .B(n2215), .S(ADD_RD1[3]), .Z(n2217) );
  MUX2_X1 U1235 ( .A(n2217), .B(n2214), .S(ADD_RD1[2]), .Z(n2218) );
  MUX2_X1 U1236 ( .A(\REGISTERS[12][5] ), .B(\REGISTERS[28][5] ), .S(
        ADD_RD1[4]), .Z(n2219) );
  MUX2_X1 U1237 ( .A(\REGISTERS[4][5] ), .B(\REGISTERS[20][5] ), .S(ADD_RD1[4]), .Z(n2220) );
  MUX2_X1 U1238 ( .A(n2220), .B(n2219), .S(ADD_RD1[3]), .Z(n2221) );
  MUX2_X1 U1239 ( .A(\REGISTERS[8][5] ), .B(\REGISTERS[24][5] ), .S(ADD_RD1[4]), .Z(n2222) );
  MUX2_X1 U1240 ( .A(\REGISTERS[0][5] ), .B(\REGISTERS[16][5] ), .S(ADD_RD1[4]), .Z(n2223) );
  MUX2_X1 U1241 ( .A(n2223), .B(n2222), .S(ADD_RD1[3]), .Z(n2224) );
  MUX2_X1 U1242 ( .A(n2224), .B(n2221), .S(ADD_RD1[2]), .Z(n2225) );
  MUX2_X1 U1243 ( .A(n2225), .B(n2218), .S(ADD_RD1[0]), .Z(n2226) );
  MUX2_X1 U1244 ( .A(n2226), .B(n2211), .S(ADD_RD1[1]), .Z(N384) );
  MUX2_X1 U1245 ( .A(\REGISTERS[15][6] ), .B(\REGISTERS[31][6] ), .S(
        ADD_RD1[4]), .Z(n2227) );
  MUX2_X1 U1246 ( .A(\REGISTERS[7][6] ), .B(\REGISTERS[23][6] ), .S(ADD_RD1[4]), .Z(n2228) );
  MUX2_X1 U1247 ( .A(n2228), .B(n2227), .S(ADD_RD1[3]), .Z(n2229) );
  MUX2_X1 U1248 ( .A(\REGISTERS[11][6] ), .B(\REGISTERS[27][6] ), .S(
        ADD_RD1[4]), .Z(n2230) );
  MUX2_X1 U1249 ( .A(\REGISTERS[3][6] ), .B(\REGISTERS[19][6] ), .S(ADD_RD1[4]), .Z(n2231) );
  MUX2_X1 U1250 ( .A(n2231), .B(n2230), .S(ADD_RD1[3]), .Z(n2232) );
  MUX2_X1 U1251 ( .A(n2232), .B(n2229), .S(ADD_RD1[2]), .Z(n2233) );
  MUX2_X1 U1252 ( .A(\REGISTERS[14][6] ), .B(\REGISTERS[30][6] ), .S(
        ADD_RD1[4]), .Z(n2234) );
  MUX2_X1 U1253 ( .A(\REGISTERS[6][6] ), .B(\REGISTERS[22][6] ), .S(ADD_RD1[4]), .Z(n2235) );
  MUX2_X1 U1254 ( .A(n2235), .B(n2234), .S(ADD_RD1[3]), .Z(n2236) );
  MUX2_X1 U1255 ( .A(\REGISTERS[10][6] ), .B(\REGISTERS[26][6] ), .S(
        ADD_RD1[4]), .Z(n2237) );
  MUX2_X1 U1256 ( .A(\REGISTERS[2][6] ), .B(\REGISTERS[18][6] ), .S(ADD_RD1[4]), .Z(n2238) );
  MUX2_X1 U1257 ( .A(n2238), .B(n2237), .S(ADD_RD1[3]), .Z(n2239) );
  MUX2_X1 U1258 ( .A(n2239), .B(n2236), .S(ADD_RD1[2]), .Z(n2240) );
  MUX2_X1 U1259 ( .A(n2240), .B(n2233), .S(ADD_RD1[0]), .Z(n2241) );
  MUX2_X1 U1260 ( .A(\REGISTERS[13][6] ), .B(\REGISTERS[29][6] ), .S(
        ADD_RD1[4]), .Z(n2242) );
  MUX2_X1 U1261 ( .A(\REGISTERS[5][6] ), .B(\REGISTERS[21][6] ), .S(ADD_RD1[4]), .Z(n2243) );
  MUX2_X1 U1262 ( .A(n2243), .B(n2242), .S(ADD_RD1[3]), .Z(n2244) );
  MUX2_X1 U1263 ( .A(\REGISTERS[9][6] ), .B(\REGISTERS[25][6] ), .S(ADD_RD1[4]), .Z(n2245) );
  MUX2_X1 U1264 ( .A(\REGISTERS[1][6] ), .B(\REGISTERS[17][6] ), .S(ADD_RD1[4]), .Z(n2246) );
  MUX2_X1 U1265 ( .A(n2246), .B(n2245), .S(ADD_RD1[3]), .Z(n2247) );
  MUX2_X1 U1266 ( .A(n2247), .B(n2244), .S(ADD_RD1[2]), .Z(n2248) );
  MUX2_X1 U1267 ( .A(\REGISTERS[12][6] ), .B(\REGISTERS[28][6] ), .S(
        ADD_RD1[4]), .Z(n2249) );
  MUX2_X1 U1268 ( .A(\REGISTERS[4][6] ), .B(\REGISTERS[20][6] ), .S(ADD_RD1[4]), .Z(n2250) );
  MUX2_X1 U1269 ( .A(n2250), .B(n2249), .S(ADD_RD1[3]), .Z(n2251) );
  MUX2_X1 U1270 ( .A(\REGISTERS[8][6] ), .B(\REGISTERS[24][6] ), .S(ADD_RD1[4]), .Z(n2252) );
  MUX2_X1 U1271 ( .A(\REGISTERS[0][6] ), .B(\REGISTERS[16][6] ), .S(ADD_RD1[4]), .Z(n2253) );
  MUX2_X1 U1272 ( .A(n2253), .B(n2252), .S(ADD_RD1[3]), .Z(n2254) );
  MUX2_X1 U1273 ( .A(n2254), .B(n2251), .S(ADD_RD1[2]), .Z(n2255) );
  MUX2_X1 U1274 ( .A(n2255), .B(n2248), .S(ADD_RD1[0]), .Z(n2256) );
  MUX2_X1 U1275 ( .A(n2256), .B(n2241), .S(ADD_RD1[1]), .Z(N385) );
  MUX2_X1 U1276 ( .A(\REGISTERS[15][7] ), .B(\REGISTERS[31][7] ), .S(
        ADD_RD1[4]), .Z(n2257) );
  MUX2_X1 U1277 ( .A(\REGISTERS[7][7] ), .B(\REGISTERS[23][7] ), .S(ADD_RD1[4]), .Z(n2258) );
  MUX2_X1 U1278 ( .A(n2258), .B(n2257), .S(ADD_RD1[3]), .Z(n2259) );
  MUX2_X1 U1279 ( .A(\REGISTERS[11][7] ), .B(\REGISTERS[27][7] ), .S(
        ADD_RD1[4]), .Z(n2260) );
  MUX2_X1 U1280 ( .A(\REGISTERS[3][7] ), .B(\REGISTERS[19][7] ), .S(ADD_RD1[4]), .Z(n2261) );
  MUX2_X1 U1281 ( .A(n2261), .B(n2260), .S(ADD_RD1[3]), .Z(n2262) );
  MUX2_X1 U1282 ( .A(n2262), .B(n2259), .S(ADD_RD1[2]), .Z(n2263) );
  MUX2_X1 U1283 ( .A(\REGISTERS[14][7] ), .B(\REGISTERS[30][7] ), .S(
        ADD_RD1[4]), .Z(n2264) );
  MUX2_X1 U1284 ( .A(\REGISTERS[6][7] ), .B(\REGISTERS[22][7] ), .S(ADD_RD1[4]), .Z(n2265) );
  MUX2_X1 U1285 ( .A(n2265), .B(n2264), .S(ADD_RD1[3]), .Z(n2266) );
  MUX2_X1 U1286 ( .A(\REGISTERS[10][7] ), .B(\REGISTERS[26][7] ), .S(
        ADD_RD1[4]), .Z(n2267) );
  MUX2_X1 U1287 ( .A(\REGISTERS[2][7] ), .B(\REGISTERS[18][7] ), .S(ADD_RD1[4]), .Z(n2268) );
  MUX2_X1 U1288 ( .A(n2268), .B(n2267), .S(ADD_RD1[3]), .Z(n2269) );
  MUX2_X1 U1289 ( .A(n2269), .B(n2266), .S(ADD_RD1[2]), .Z(n2270) );
  MUX2_X1 U1290 ( .A(n2270), .B(n2263), .S(ADD_RD1[0]), .Z(n2271) );
  MUX2_X1 U1291 ( .A(\REGISTERS[13][7] ), .B(\REGISTERS[29][7] ), .S(
        ADD_RD1[4]), .Z(n2272) );
  MUX2_X1 U1292 ( .A(\REGISTERS[5][7] ), .B(\REGISTERS[21][7] ), .S(ADD_RD1[4]), .Z(n2273) );
  MUX2_X1 U1293 ( .A(n2273), .B(n2272), .S(ADD_RD1[3]), .Z(n2274) );
  MUX2_X1 U1294 ( .A(\REGISTERS[9][7] ), .B(\REGISTERS[25][7] ), .S(ADD_RD1[4]), .Z(n2275) );
  MUX2_X1 U1295 ( .A(\REGISTERS[1][7] ), .B(\REGISTERS[17][7] ), .S(ADD_RD1[4]), .Z(n2276) );
  MUX2_X1 U1296 ( .A(n2276), .B(n2275), .S(ADD_RD1[3]), .Z(n2277) );
  MUX2_X1 U1297 ( .A(n2277), .B(n2274), .S(ADD_RD1[2]), .Z(n2278) );
  MUX2_X1 U1298 ( .A(\REGISTERS[12][7] ), .B(\REGISTERS[28][7] ), .S(
        ADD_RD1[4]), .Z(n2279) );
  MUX2_X1 U1299 ( .A(\REGISTERS[4][7] ), .B(\REGISTERS[20][7] ), .S(ADD_RD1[4]), .Z(n2280) );
  MUX2_X1 U1300 ( .A(n2280), .B(n2279), .S(ADD_RD1[3]), .Z(n2281) );
  MUX2_X1 U1301 ( .A(\REGISTERS[8][7] ), .B(\REGISTERS[24][7] ), .S(ADD_RD1[4]), .Z(n2282) );
  MUX2_X1 U1302 ( .A(\REGISTERS[0][7] ), .B(\REGISTERS[16][7] ), .S(ADD_RD1[4]), .Z(n2283) );
  MUX2_X1 U1303 ( .A(n2283), .B(n2282), .S(ADD_RD1[3]), .Z(n2284) );
  MUX2_X1 U1304 ( .A(n2284), .B(n2281), .S(ADD_RD1[2]), .Z(n2285) );
  MUX2_X1 U1305 ( .A(n2285), .B(n2278), .S(ADD_RD1[0]), .Z(n2286) );
  MUX2_X1 U1306 ( .A(n2286), .B(n2271), .S(ADD_RD1[1]), .Z(N386) );
  MUX2_X1 U1307 ( .A(\REGISTERS[15][8] ), .B(\REGISTERS[31][8] ), .S(
        ADD_RD1[4]), .Z(n2287) );
  MUX2_X1 U1308 ( .A(\REGISTERS[7][8] ), .B(\REGISTERS[23][8] ), .S(ADD_RD1[4]), .Z(n2288) );
  MUX2_X1 U1309 ( .A(n2288), .B(n2287), .S(ADD_RD1[3]), .Z(n2289) );
  MUX2_X1 U1310 ( .A(\REGISTERS[11][8] ), .B(\REGISTERS[27][8] ), .S(
        ADD_RD1[4]), .Z(n2290) );
  MUX2_X1 U1311 ( .A(\REGISTERS[3][8] ), .B(\REGISTERS[19][8] ), .S(ADD_RD1[4]), .Z(n2291) );
  MUX2_X1 U1312 ( .A(n2291), .B(n2290), .S(ADD_RD1[3]), .Z(n2292) );
  MUX2_X1 U1313 ( .A(n2292), .B(n2289), .S(ADD_RD1[2]), .Z(n2293) );
  MUX2_X1 U1314 ( .A(\REGISTERS[14][8] ), .B(\REGISTERS[30][8] ), .S(
        ADD_RD1[4]), .Z(n2294) );
  MUX2_X1 U1315 ( .A(\REGISTERS[6][8] ), .B(\REGISTERS[22][8] ), .S(ADD_RD1[4]), .Z(n2295) );
  MUX2_X1 U1316 ( .A(n2295), .B(n2294), .S(ADD_RD1[3]), .Z(n2296) );
  MUX2_X1 U1317 ( .A(\REGISTERS[10][8] ), .B(\REGISTERS[26][8] ), .S(
        ADD_RD1[4]), .Z(n2297) );
  MUX2_X1 U1318 ( .A(\REGISTERS[2][8] ), .B(\REGISTERS[18][8] ), .S(ADD_RD1[4]), .Z(n2298) );
  MUX2_X1 U1319 ( .A(n2298), .B(n2297), .S(ADD_RD1[3]), .Z(n2299) );
  MUX2_X1 U1320 ( .A(n2299), .B(n2296), .S(ADD_RD1[2]), .Z(n2300) );
  MUX2_X1 U1321 ( .A(n2300), .B(n2293), .S(ADD_RD1[0]), .Z(n2301) );
  MUX2_X1 U1322 ( .A(\REGISTERS[13][8] ), .B(\REGISTERS[29][8] ), .S(
        ADD_RD1[4]), .Z(n2302) );
  MUX2_X1 U1323 ( .A(\REGISTERS[5][8] ), .B(\REGISTERS[21][8] ), .S(ADD_RD1[4]), .Z(n2303) );
  MUX2_X1 U1324 ( .A(n2303), .B(n2302), .S(ADD_RD1[3]), .Z(n2304) );
  MUX2_X1 U1325 ( .A(\REGISTERS[9][8] ), .B(\REGISTERS[25][8] ), .S(ADD_RD1[4]), .Z(n2305) );
  MUX2_X1 U1326 ( .A(\REGISTERS[1][8] ), .B(\REGISTERS[17][8] ), .S(ADD_RD1[4]), .Z(n2306) );
  MUX2_X1 U1327 ( .A(n2306), .B(n2305), .S(ADD_RD1[3]), .Z(n2307) );
  MUX2_X1 U1328 ( .A(n2307), .B(n2304), .S(ADD_RD1[2]), .Z(n2308) );
  MUX2_X1 U1329 ( .A(\REGISTERS[12][8] ), .B(\REGISTERS[28][8] ), .S(
        ADD_RD1[4]), .Z(n2309) );
  MUX2_X1 U1330 ( .A(\REGISTERS[4][8] ), .B(\REGISTERS[20][8] ), .S(ADD_RD1[4]), .Z(n2310) );
  MUX2_X1 U1331 ( .A(n2310), .B(n2309), .S(ADD_RD1[3]), .Z(n2311) );
  MUX2_X1 U1332 ( .A(\REGISTERS[8][8] ), .B(\REGISTERS[24][8] ), .S(ADD_RD1[4]), .Z(n2312) );
  MUX2_X1 U1333 ( .A(\REGISTERS[0][8] ), .B(\REGISTERS[16][8] ), .S(ADD_RD1[4]), .Z(n2313) );
  MUX2_X1 U1334 ( .A(n2313), .B(n2312), .S(ADD_RD1[3]), .Z(n2314) );
  MUX2_X1 U1335 ( .A(n2314), .B(n2311), .S(ADD_RD1[2]), .Z(n2315) );
  MUX2_X1 U1336 ( .A(n2315), .B(n2308), .S(ADD_RD1[0]), .Z(n2316) );
  MUX2_X1 U1337 ( .A(n2316), .B(n2301), .S(ADD_RD1[1]), .Z(N387) );
  MUX2_X1 U1338 ( .A(\REGISTERS[15][9] ), .B(\REGISTERS[31][9] ), .S(
        ADD_RD1[4]), .Z(n2317) );
  MUX2_X1 U1339 ( .A(\REGISTERS[7][9] ), .B(\REGISTERS[23][9] ), .S(ADD_RD1[4]), .Z(n2318) );
  MUX2_X1 U1340 ( .A(n2318), .B(n2317), .S(ADD_RD1[3]), .Z(n2319) );
  MUX2_X1 U1341 ( .A(\REGISTERS[11][9] ), .B(\REGISTERS[27][9] ), .S(
        ADD_RD1[4]), .Z(n2320) );
  MUX2_X1 U1342 ( .A(\REGISTERS[3][9] ), .B(\REGISTERS[19][9] ), .S(ADD_RD1[4]), .Z(n2321) );
  MUX2_X1 U1343 ( .A(n2321), .B(n2320), .S(ADD_RD1[3]), .Z(n2322) );
  MUX2_X1 U1344 ( .A(n2322), .B(n2319), .S(ADD_RD1[2]), .Z(n2323) );
  MUX2_X1 U1345 ( .A(\REGISTERS[14][9] ), .B(\REGISTERS[30][9] ), .S(
        ADD_RD1[4]), .Z(n2324) );
  MUX2_X1 U1346 ( .A(\REGISTERS[6][9] ), .B(\REGISTERS[22][9] ), .S(ADD_RD1[4]), .Z(n2325) );
  MUX2_X1 U1347 ( .A(n2325), .B(n2324), .S(ADD_RD1[3]), .Z(n2326) );
  MUX2_X1 U1348 ( .A(\REGISTERS[10][9] ), .B(\REGISTERS[26][9] ), .S(
        ADD_RD1[4]), .Z(n2327) );
  MUX2_X1 U1349 ( .A(\REGISTERS[2][9] ), .B(\REGISTERS[18][9] ), .S(ADD_RD1[4]), .Z(n2328) );
  MUX2_X1 U1350 ( .A(n2328), .B(n2327), .S(ADD_RD1[3]), .Z(n2329) );
  MUX2_X1 U1351 ( .A(n2329), .B(n2326), .S(ADD_RD1[2]), .Z(n2330) );
  MUX2_X1 U1352 ( .A(n2330), .B(n2323), .S(ADD_RD1[0]), .Z(n2331) );
  MUX2_X1 U1353 ( .A(\REGISTERS[13][9] ), .B(\REGISTERS[29][9] ), .S(
        ADD_RD1[4]), .Z(n2332) );
  MUX2_X1 U1354 ( .A(\REGISTERS[5][9] ), .B(\REGISTERS[21][9] ), .S(ADD_RD1[4]), .Z(n2333) );
  MUX2_X1 U1355 ( .A(n2333), .B(n2332), .S(ADD_RD1[3]), .Z(n2334) );
  MUX2_X1 U1356 ( .A(\REGISTERS[9][9] ), .B(\REGISTERS[25][9] ), .S(ADD_RD1[4]), .Z(n2335) );
  MUX2_X1 U1357 ( .A(\REGISTERS[1][9] ), .B(\REGISTERS[17][9] ), .S(ADD_RD1[4]), .Z(n2336) );
  MUX2_X1 U1358 ( .A(n2336), .B(n2335), .S(ADD_RD1[3]), .Z(n2337) );
  MUX2_X1 U1359 ( .A(n2337), .B(n2334), .S(ADD_RD1[2]), .Z(n2338) );
  MUX2_X1 U1360 ( .A(\REGISTERS[12][9] ), .B(\REGISTERS[28][9] ), .S(
        ADD_RD1[4]), .Z(n2339) );
  MUX2_X1 U1361 ( .A(\REGISTERS[4][9] ), .B(\REGISTERS[20][9] ), .S(ADD_RD1[4]), .Z(n2340) );
  MUX2_X1 U1362 ( .A(n2340), .B(n2339), .S(ADD_RD1[3]), .Z(n2341) );
  MUX2_X1 U1363 ( .A(\REGISTERS[8][9] ), .B(\REGISTERS[24][9] ), .S(ADD_RD1[4]), .Z(n2342) );
  MUX2_X1 U1364 ( .A(\REGISTERS[0][9] ), .B(\REGISTERS[16][9] ), .S(ADD_RD1[4]), .Z(n2343) );
  MUX2_X1 U1365 ( .A(n2343), .B(n2342), .S(ADD_RD1[3]), .Z(n2344) );
  MUX2_X1 U1366 ( .A(n2344), .B(n2341), .S(ADD_RD1[2]), .Z(n2345) );
  MUX2_X1 U1367 ( .A(n2345), .B(n2338), .S(ADD_RD1[0]), .Z(n2346) );
  MUX2_X1 U1368 ( .A(n2346), .B(n2331), .S(ADD_RD1[1]), .Z(N388) );
  MUX2_X1 U1369 ( .A(\REGISTERS[15][10] ), .B(\REGISTERS[31][10] ), .S(
        ADD_RD1[4]), .Z(n2347) );
  MUX2_X1 U1370 ( .A(\REGISTERS[7][10] ), .B(\REGISTERS[23][10] ), .S(
        ADD_RD1[4]), .Z(n2348) );
  MUX2_X1 U1371 ( .A(n2348), .B(n2347), .S(ADD_RD1[3]), .Z(n2349) );
  MUX2_X1 U1372 ( .A(\REGISTERS[11][10] ), .B(\REGISTERS[27][10] ), .S(
        ADD_RD1[4]), .Z(n2350) );
  MUX2_X1 U1373 ( .A(\REGISTERS[3][10] ), .B(\REGISTERS[19][10] ), .S(
        ADD_RD1[4]), .Z(n2351) );
  MUX2_X1 U1374 ( .A(n2351), .B(n2350), .S(ADD_RD1[3]), .Z(n2352) );
  MUX2_X1 U1375 ( .A(n2352), .B(n2349), .S(ADD_RD1[2]), .Z(n2353) );
  MUX2_X1 U1376 ( .A(\REGISTERS[14][10] ), .B(\REGISTERS[30][10] ), .S(
        ADD_RD1[4]), .Z(n2354) );
  MUX2_X1 U1377 ( .A(\REGISTERS[6][10] ), .B(\REGISTERS[22][10] ), .S(
        ADD_RD1[4]), .Z(n2355) );
  MUX2_X1 U1378 ( .A(n2355), .B(n2354), .S(ADD_RD1[3]), .Z(n2356) );
  MUX2_X1 U1379 ( .A(\REGISTERS[10][10] ), .B(\REGISTERS[26][10] ), .S(
        ADD_RD1[4]), .Z(n2357) );
  MUX2_X1 U1380 ( .A(\REGISTERS[2][10] ), .B(\REGISTERS[18][10] ), .S(
        ADD_RD1[4]), .Z(n2358) );
  MUX2_X1 U1381 ( .A(n2358), .B(n2357), .S(ADD_RD1[3]), .Z(n2359) );
  MUX2_X1 U1382 ( .A(n2359), .B(n2356), .S(ADD_RD1[2]), .Z(n2360) );
  MUX2_X1 U1383 ( .A(n2360), .B(n2353), .S(ADD_RD1[0]), .Z(n2361) );
  MUX2_X1 U1384 ( .A(\REGISTERS[13][10] ), .B(\REGISTERS[29][10] ), .S(
        ADD_RD1[4]), .Z(n2362) );
  MUX2_X1 U1385 ( .A(\REGISTERS[5][10] ), .B(\REGISTERS[21][10] ), .S(
        ADD_RD1[4]), .Z(n2363) );
  MUX2_X1 U1386 ( .A(n2363), .B(n2362), .S(ADD_RD1[3]), .Z(n2364) );
  MUX2_X1 U1387 ( .A(\REGISTERS[9][10] ), .B(\REGISTERS[25][10] ), .S(
        ADD_RD1[4]), .Z(n2365) );
  MUX2_X1 U1388 ( .A(\REGISTERS[1][10] ), .B(\REGISTERS[17][10] ), .S(
        ADD_RD1[4]), .Z(n2366) );
  MUX2_X1 U1389 ( .A(n2366), .B(n2365), .S(ADD_RD1[3]), .Z(n2367) );
  MUX2_X1 U1390 ( .A(n2367), .B(n2364), .S(ADD_RD1[2]), .Z(n2368) );
  MUX2_X1 U1391 ( .A(\REGISTERS[12][10] ), .B(\REGISTERS[28][10] ), .S(
        ADD_RD1[4]), .Z(n2369) );
  MUX2_X1 U1392 ( .A(\REGISTERS[4][10] ), .B(\REGISTERS[20][10] ), .S(
        ADD_RD1[4]), .Z(n2370) );
  MUX2_X1 U1393 ( .A(n2370), .B(n2369), .S(ADD_RD1[3]), .Z(n2371) );
  MUX2_X1 U1394 ( .A(\REGISTERS[8][10] ), .B(\REGISTERS[24][10] ), .S(
        ADD_RD1[4]), .Z(n2372) );
  MUX2_X1 U1395 ( .A(\REGISTERS[0][10] ), .B(\REGISTERS[16][10] ), .S(
        ADD_RD1[4]), .Z(n2373) );
  MUX2_X1 U1396 ( .A(n2373), .B(n2372), .S(ADD_RD1[3]), .Z(n2374) );
  MUX2_X1 U1397 ( .A(n2374), .B(n2371), .S(ADD_RD1[2]), .Z(n2375) );
  MUX2_X1 U1398 ( .A(n2375), .B(n2368), .S(ADD_RD1[0]), .Z(n2376) );
  MUX2_X1 U1399 ( .A(n2376), .B(n2361), .S(ADD_RD1[1]), .Z(N389) );
  MUX2_X1 U1400 ( .A(\REGISTERS[15][11] ), .B(\REGISTERS[31][11] ), .S(
        ADD_RD1[4]), .Z(n2377) );
  MUX2_X1 U1401 ( .A(\REGISTERS[7][11] ), .B(\REGISTERS[23][11] ), .S(
        ADD_RD1[4]), .Z(n2378) );
  MUX2_X1 U1402 ( .A(n2378), .B(n2377), .S(ADD_RD1[3]), .Z(n2379) );
  MUX2_X1 U1403 ( .A(\REGISTERS[11][11] ), .B(\REGISTERS[27][11] ), .S(
        ADD_RD1[4]), .Z(n2380) );
  MUX2_X1 U1404 ( .A(\REGISTERS[3][11] ), .B(\REGISTERS[19][11] ), .S(
        ADD_RD1[4]), .Z(n2381) );
  MUX2_X1 U1405 ( .A(n2381), .B(n2380), .S(ADD_RD1[3]), .Z(n2382) );
  MUX2_X1 U1406 ( .A(n2382), .B(n2379), .S(ADD_RD1[2]), .Z(n2383) );
  MUX2_X1 U1407 ( .A(\REGISTERS[14][11] ), .B(\REGISTERS[30][11] ), .S(
        ADD_RD1[4]), .Z(n2384) );
  MUX2_X1 U1408 ( .A(\REGISTERS[6][11] ), .B(\REGISTERS[22][11] ), .S(
        ADD_RD1[4]), .Z(n2385) );
  MUX2_X1 U1409 ( .A(n2385), .B(n2384), .S(ADD_RD1[3]), .Z(n2386) );
  MUX2_X1 U1410 ( .A(\REGISTERS[10][11] ), .B(\REGISTERS[26][11] ), .S(
        ADD_RD1[4]), .Z(n2387) );
  MUX2_X1 U1411 ( .A(\REGISTERS[2][11] ), .B(\REGISTERS[18][11] ), .S(
        ADD_RD1[4]), .Z(n2388) );
  MUX2_X1 U1412 ( .A(n2388), .B(n2387), .S(ADD_RD1[3]), .Z(n2389) );
  MUX2_X1 U1413 ( .A(n2389), .B(n2386), .S(ADD_RD1[2]), .Z(n2390) );
  MUX2_X1 U1414 ( .A(n2390), .B(n2383), .S(ADD_RD1[0]), .Z(n2391) );
  MUX2_X1 U1415 ( .A(\REGISTERS[13][11] ), .B(\REGISTERS[29][11] ), .S(
        ADD_RD1[4]), .Z(n2392) );
  MUX2_X1 U1416 ( .A(\REGISTERS[5][11] ), .B(\REGISTERS[21][11] ), .S(
        ADD_RD1[4]), .Z(n2393) );
  MUX2_X1 U1417 ( .A(n2393), .B(n2392), .S(ADD_RD1[3]), .Z(n2394) );
  MUX2_X1 U1418 ( .A(\REGISTERS[9][11] ), .B(\REGISTERS[25][11] ), .S(
        ADD_RD1[4]), .Z(n2395) );
  MUX2_X1 U1419 ( .A(\REGISTERS[1][11] ), .B(\REGISTERS[17][11] ), .S(
        ADD_RD1[4]), .Z(n2396) );
  MUX2_X1 U1420 ( .A(n2396), .B(n2395), .S(ADD_RD1[3]), .Z(n2397) );
  MUX2_X1 U1421 ( .A(n2397), .B(n2394), .S(ADD_RD1[2]), .Z(n2398) );
  MUX2_X1 U1422 ( .A(\REGISTERS[12][11] ), .B(\REGISTERS[28][11] ), .S(
        ADD_RD1[4]), .Z(n2399) );
  MUX2_X1 U1423 ( .A(\REGISTERS[4][11] ), .B(\REGISTERS[20][11] ), .S(
        ADD_RD1[4]), .Z(n2400) );
  MUX2_X1 U1424 ( .A(n2400), .B(n2399), .S(ADD_RD1[3]), .Z(n2401) );
  MUX2_X1 U1425 ( .A(\REGISTERS[8][11] ), .B(\REGISTERS[24][11] ), .S(
        ADD_RD1[4]), .Z(n2402) );
  MUX2_X1 U1426 ( .A(\REGISTERS[0][11] ), .B(\REGISTERS[16][11] ), .S(
        ADD_RD1[4]), .Z(n2403) );
  MUX2_X1 U1427 ( .A(n2403), .B(n2402), .S(ADD_RD1[3]), .Z(n2404) );
  MUX2_X1 U1428 ( .A(n2404), .B(n2401), .S(ADD_RD1[2]), .Z(n2405) );
  MUX2_X1 U1429 ( .A(n2405), .B(n2398), .S(ADD_RD1[0]), .Z(n2406) );
  MUX2_X1 U1430 ( .A(n2406), .B(n2391), .S(ADD_RD1[1]), .Z(N390) );
  MUX2_X1 U1431 ( .A(\REGISTERS[15][12] ), .B(\REGISTERS[31][12] ), .S(
        ADD_RD1[4]), .Z(n2407) );
  MUX2_X1 U1432 ( .A(\REGISTERS[7][12] ), .B(\REGISTERS[23][12] ), .S(
        ADD_RD1[4]), .Z(n2408) );
  MUX2_X1 U1433 ( .A(n2408), .B(n2407), .S(ADD_RD1[3]), .Z(n2409) );
  MUX2_X1 U1434 ( .A(\REGISTERS[11][12] ), .B(\REGISTERS[27][12] ), .S(
        ADD_RD1[4]), .Z(n2410) );
  MUX2_X1 U1435 ( .A(\REGISTERS[3][12] ), .B(\REGISTERS[19][12] ), .S(
        ADD_RD1[4]), .Z(n2411) );
  MUX2_X1 U1436 ( .A(n2411), .B(n2410), .S(ADD_RD1[3]), .Z(n2412) );
  MUX2_X1 U1437 ( .A(n2412), .B(n2409), .S(ADD_RD1[2]), .Z(n2413) );
  MUX2_X1 U1438 ( .A(\REGISTERS[14][12] ), .B(\REGISTERS[30][12] ), .S(
        ADD_RD1[4]), .Z(n2414) );
  MUX2_X1 U1439 ( .A(\REGISTERS[6][12] ), .B(\REGISTERS[22][12] ), .S(
        ADD_RD1[4]), .Z(n2415) );
  MUX2_X1 U1440 ( .A(n2415), .B(n2414), .S(ADD_RD1[3]), .Z(n2416) );
  MUX2_X1 U1441 ( .A(\REGISTERS[10][12] ), .B(\REGISTERS[26][12] ), .S(
        ADD_RD1[4]), .Z(n2417) );
  MUX2_X1 U1442 ( .A(\REGISTERS[2][12] ), .B(\REGISTERS[18][12] ), .S(
        ADD_RD1[4]), .Z(n2418) );
  MUX2_X1 U1443 ( .A(n2418), .B(n2417), .S(ADD_RD1[3]), .Z(n2419) );
  MUX2_X1 U1444 ( .A(n2419), .B(n2416), .S(ADD_RD1[2]), .Z(n2420) );
  MUX2_X1 U1445 ( .A(n2420), .B(n2413), .S(ADD_RD1[0]), .Z(n2421) );
  MUX2_X1 U1446 ( .A(\REGISTERS[13][12] ), .B(\REGISTERS[29][12] ), .S(
        ADD_RD1[4]), .Z(n2422) );
  MUX2_X1 U1447 ( .A(\REGISTERS[5][12] ), .B(\REGISTERS[21][12] ), .S(
        ADD_RD1[4]), .Z(n2423) );
  MUX2_X1 U1448 ( .A(n2423), .B(n2422), .S(ADD_RD1[3]), .Z(n2424) );
  MUX2_X1 U1449 ( .A(\REGISTERS[9][12] ), .B(\REGISTERS[25][12] ), .S(
        ADD_RD1[4]), .Z(n2425) );
  MUX2_X1 U1450 ( .A(\REGISTERS[1][12] ), .B(\REGISTERS[17][12] ), .S(
        ADD_RD1[4]), .Z(n2426) );
  MUX2_X1 U1451 ( .A(n2426), .B(n2425), .S(ADD_RD1[3]), .Z(n2427) );
  MUX2_X1 U1452 ( .A(n2427), .B(n2424), .S(ADD_RD1[2]), .Z(n2428) );
  MUX2_X1 U1453 ( .A(\REGISTERS[12][12] ), .B(\REGISTERS[28][12] ), .S(
        ADD_RD1[4]), .Z(n2429) );
  MUX2_X1 U1454 ( .A(\REGISTERS[4][12] ), .B(\REGISTERS[20][12] ), .S(
        ADD_RD1[4]), .Z(n2430) );
  MUX2_X1 U1455 ( .A(n2430), .B(n2429), .S(ADD_RD1[3]), .Z(n2431) );
  MUX2_X1 U1456 ( .A(\REGISTERS[8][12] ), .B(\REGISTERS[24][12] ), .S(
        ADD_RD1[4]), .Z(n2432) );
  MUX2_X1 U1457 ( .A(\REGISTERS[0][12] ), .B(\REGISTERS[16][12] ), .S(
        ADD_RD1[4]), .Z(n2433) );
  MUX2_X1 U1458 ( .A(n2433), .B(n2432), .S(ADD_RD1[3]), .Z(n2434) );
  MUX2_X1 U1459 ( .A(n2434), .B(n2431), .S(ADD_RD1[2]), .Z(n2435) );
  MUX2_X1 U1460 ( .A(n2435), .B(n2428), .S(ADD_RD1[0]), .Z(n2436) );
  MUX2_X1 U1461 ( .A(n2436), .B(n2421), .S(ADD_RD1[1]), .Z(N391) );
  MUX2_X1 U1462 ( .A(\REGISTERS[15][13] ), .B(\REGISTERS[31][13] ), .S(
        ADD_RD1[4]), .Z(n2437) );
  MUX2_X1 U1463 ( .A(\REGISTERS[7][13] ), .B(\REGISTERS[23][13] ), .S(
        ADD_RD1[4]), .Z(n2438) );
  MUX2_X1 U1464 ( .A(n2438), .B(n2437), .S(ADD_RD1[3]), .Z(n2439) );
  MUX2_X1 U1465 ( .A(\REGISTERS[11][13] ), .B(\REGISTERS[27][13] ), .S(
        ADD_RD1[4]), .Z(n2440) );
  MUX2_X1 U1466 ( .A(\REGISTERS[3][13] ), .B(\REGISTERS[19][13] ), .S(
        ADD_RD1[4]), .Z(n2441) );
  MUX2_X1 U1467 ( .A(n2441), .B(n2440), .S(ADD_RD1[3]), .Z(n2442) );
  MUX2_X1 U1468 ( .A(n2442), .B(n2439), .S(ADD_RD1[2]), .Z(n2443) );
  MUX2_X1 U1469 ( .A(\REGISTERS[14][13] ), .B(\REGISTERS[30][13] ), .S(
        ADD_RD1[4]), .Z(n2444) );
  MUX2_X1 U1470 ( .A(\REGISTERS[6][13] ), .B(\REGISTERS[22][13] ), .S(
        ADD_RD1[4]), .Z(n2445) );
  MUX2_X1 U1471 ( .A(n2445), .B(n2444), .S(ADD_RD1[3]), .Z(n2446) );
  MUX2_X1 U1472 ( .A(\REGISTERS[10][13] ), .B(\REGISTERS[26][13] ), .S(
        ADD_RD1[4]), .Z(n2447) );
  MUX2_X1 U1473 ( .A(\REGISTERS[2][13] ), .B(\REGISTERS[18][13] ), .S(
        ADD_RD1[4]), .Z(n2448) );
  MUX2_X1 U1474 ( .A(n2448), .B(n2447), .S(ADD_RD1[3]), .Z(n2449) );
  MUX2_X1 U1475 ( .A(n2449), .B(n2446), .S(ADD_RD1[2]), .Z(n2450) );
  MUX2_X1 U1476 ( .A(n2450), .B(n2443), .S(ADD_RD1[0]), .Z(n2451) );
  MUX2_X1 U1477 ( .A(\REGISTERS[13][13] ), .B(\REGISTERS[29][13] ), .S(
        ADD_RD1[4]), .Z(n2452) );
  MUX2_X1 U1478 ( .A(\REGISTERS[5][13] ), .B(\REGISTERS[21][13] ), .S(
        ADD_RD1[4]), .Z(n2453) );
  MUX2_X1 U1479 ( .A(n2453), .B(n2452), .S(ADD_RD1[3]), .Z(n2454) );
  MUX2_X1 U1480 ( .A(\REGISTERS[9][13] ), .B(\REGISTERS[25][13] ), .S(
        ADD_RD1[4]), .Z(n2455) );
  MUX2_X1 U1481 ( .A(\REGISTERS[1][13] ), .B(\REGISTERS[17][13] ), .S(
        ADD_RD1[4]), .Z(n2456) );
  MUX2_X1 U1482 ( .A(n2456), .B(n2455), .S(ADD_RD1[3]), .Z(n2457) );
  MUX2_X1 U1483 ( .A(n2457), .B(n2454), .S(ADD_RD1[2]), .Z(n2458) );
  MUX2_X1 U1484 ( .A(\REGISTERS[12][13] ), .B(\REGISTERS[28][13] ), .S(
        ADD_RD1[4]), .Z(n2459) );
  MUX2_X1 U1485 ( .A(\REGISTERS[4][13] ), .B(\REGISTERS[20][13] ), .S(
        ADD_RD1[4]), .Z(n2460) );
  MUX2_X1 U1486 ( .A(n2460), .B(n2459), .S(ADD_RD1[3]), .Z(n2461) );
  MUX2_X1 U1487 ( .A(\REGISTERS[8][13] ), .B(\REGISTERS[24][13] ), .S(
        ADD_RD1[4]), .Z(n2462) );
  MUX2_X1 U1488 ( .A(\REGISTERS[0][13] ), .B(\REGISTERS[16][13] ), .S(
        ADD_RD1[4]), .Z(n2463) );
  MUX2_X1 U1489 ( .A(n2463), .B(n2462), .S(ADD_RD1[3]), .Z(n2464) );
  MUX2_X1 U1490 ( .A(n2464), .B(n2461), .S(ADD_RD1[2]), .Z(n2465) );
  MUX2_X1 U1491 ( .A(n2465), .B(n2458), .S(ADD_RD1[0]), .Z(n2466) );
  MUX2_X1 U1492 ( .A(n2466), .B(n2451), .S(ADD_RD1[1]), .Z(N392) );
  MUX2_X1 U1493 ( .A(\REGISTERS[15][14] ), .B(\REGISTERS[31][14] ), .S(
        ADD_RD1[4]), .Z(n2467) );
  MUX2_X1 U1494 ( .A(\REGISTERS[7][14] ), .B(\REGISTERS[23][14] ), .S(
        ADD_RD1[4]), .Z(n2468) );
  MUX2_X1 U1495 ( .A(n2468), .B(n2467), .S(ADD_RD1[3]), .Z(n2469) );
  MUX2_X1 U1496 ( .A(\REGISTERS[11][14] ), .B(\REGISTERS[27][14] ), .S(
        ADD_RD1[4]), .Z(n2470) );
  MUX2_X1 U1497 ( .A(\REGISTERS[3][14] ), .B(\REGISTERS[19][14] ), .S(
        ADD_RD1[4]), .Z(n2471) );
  MUX2_X1 U1498 ( .A(n2471), .B(n2470), .S(ADD_RD1[3]), .Z(n2472) );
  MUX2_X1 U1499 ( .A(n2472), .B(n2469), .S(ADD_RD1[2]), .Z(n2473) );
  MUX2_X1 U1500 ( .A(\REGISTERS[14][14] ), .B(\REGISTERS[30][14] ), .S(
        ADD_RD1[4]), .Z(n2474) );
  MUX2_X1 U1501 ( .A(\REGISTERS[6][14] ), .B(\REGISTERS[22][14] ), .S(
        ADD_RD1[4]), .Z(n2475) );
  MUX2_X1 U1502 ( .A(n2475), .B(n2474), .S(ADD_RD1[3]), .Z(n2476) );
  MUX2_X1 U1503 ( .A(\REGISTERS[10][14] ), .B(\REGISTERS[26][14] ), .S(
        ADD_RD1[4]), .Z(n2477) );
  MUX2_X1 U1504 ( .A(\REGISTERS[2][14] ), .B(\REGISTERS[18][14] ), .S(
        ADD_RD1[4]), .Z(n2478) );
  MUX2_X1 U1505 ( .A(n2478), .B(n2477), .S(ADD_RD1[3]), .Z(n2479) );
  MUX2_X1 U1506 ( .A(n2479), .B(n2476), .S(ADD_RD1[2]), .Z(n2480) );
  MUX2_X1 U1507 ( .A(n2480), .B(n2473), .S(ADD_RD1[0]), .Z(n2481) );
  MUX2_X1 U1508 ( .A(\REGISTERS[13][14] ), .B(\REGISTERS[29][14] ), .S(
        ADD_RD1[4]), .Z(n2482) );
  MUX2_X1 U1509 ( .A(\REGISTERS[5][14] ), .B(\REGISTERS[21][14] ), .S(
        ADD_RD1[4]), .Z(n2483) );
  MUX2_X1 U1510 ( .A(n2483), .B(n2482), .S(ADD_RD1[3]), .Z(n2484) );
  MUX2_X1 U1511 ( .A(\REGISTERS[9][14] ), .B(\REGISTERS[25][14] ), .S(
        ADD_RD1[4]), .Z(n2485) );
  MUX2_X1 U1512 ( .A(\REGISTERS[1][14] ), .B(\REGISTERS[17][14] ), .S(
        ADD_RD1[4]), .Z(n2486) );
  MUX2_X1 U1513 ( .A(n2486), .B(n2485), .S(ADD_RD1[3]), .Z(n2487) );
  MUX2_X1 U1514 ( .A(n2487), .B(n2484), .S(ADD_RD1[2]), .Z(n2488) );
  MUX2_X1 U1515 ( .A(\REGISTERS[12][14] ), .B(\REGISTERS[28][14] ), .S(
        ADD_RD1[4]), .Z(n2489) );
  MUX2_X1 U1516 ( .A(\REGISTERS[4][14] ), .B(\REGISTERS[20][14] ), .S(
        ADD_RD1[4]), .Z(n2490) );
  MUX2_X1 U1517 ( .A(n2490), .B(n2489), .S(ADD_RD1[3]), .Z(n2491) );
  MUX2_X1 U1518 ( .A(\REGISTERS[8][14] ), .B(\REGISTERS[24][14] ), .S(
        ADD_RD1[4]), .Z(n2492) );
  MUX2_X1 U1519 ( .A(\REGISTERS[0][14] ), .B(\REGISTERS[16][14] ), .S(
        ADD_RD1[4]), .Z(n2493) );
  MUX2_X1 U1520 ( .A(n2493), .B(n2492), .S(ADD_RD1[3]), .Z(n2494) );
  MUX2_X1 U1521 ( .A(n2494), .B(n2491), .S(ADD_RD1[2]), .Z(n2495) );
  MUX2_X1 U1522 ( .A(n2495), .B(n2488), .S(ADD_RD1[0]), .Z(n2496) );
  MUX2_X1 U1523 ( .A(n2496), .B(n2481), .S(ADD_RD1[1]), .Z(N393) );
  MUX2_X1 U1524 ( .A(\REGISTERS[15][15] ), .B(\REGISTERS[31][15] ), .S(
        ADD_RD1[4]), .Z(n2497) );
  MUX2_X1 U1525 ( .A(\REGISTERS[7][15] ), .B(\REGISTERS[23][15] ), .S(
        ADD_RD1[4]), .Z(n2498) );
  MUX2_X1 U1526 ( .A(n2498), .B(n2497), .S(ADD_RD1[3]), .Z(n2499) );
  MUX2_X1 U1527 ( .A(\REGISTERS[11][15] ), .B(\REGISTERS[27][15] ), .S(
        ADD_RD1[4]), .Z(n2500) );
  MUX2_X1 U1528 ( .A(\REGISTERS[3][15] ), .B(\REGISTERS[19][15] ), .S(
        ADD_RD1[4]), .Z(n2501) );
  MUX2_X1 U1529 ( .A(n2501), .B(n2500), .S(ADD_RD1[3]), .Z(n2502) );
  MUX2_X1 U1530 ( .A(n2502), .B(n2499), .S(ADD_RD1[2]), .Z(n2503) );
  MUX2_X1 U1531 ( .A(\REGISTERS[14][15] ), .B(\REGISTERS[30][15] ), .S(
        ADD_RD1[4]), .Z(n2504) );
  MUX2_X1 U1532 ( .A(\REGISTERS[6][15] ), .B(\REGISTERS[22][15] ), .S(
        ADD_RD1[4]), .Z(n2505) );
  MUX2_X1 U1533 ( .A(n2505), .B(n2504), .S(ADD_RD1[3]), .Z(n2506) );
  MUX2_X1 U1534 ( .A(\REGISTERS[10][15] ), .B(\REGISTERS[26][15] ), .S(
        ADD_RD1[4]), .Z(n2507) );
  MUX2_X1 U1535 ( .A(\REGISTERS[2][15] ), .B(\REGISTERS[18][15] ), .S(
        ADD_RD1[4]), .Z(n2508) );
  MUX2_X1 U1536 ( .A(n2508), .B(n2507), .S(ADD_RD1[3]), .Z(n2509) );
  MUX2_X1 U1537 ( .A(n2509), .B(n2506), .S(ADD_RD1[2]), .Z(n2510) );
  MUX2_X1 U1538 ( .A(n2510), .B(n2503), .S(ADD_RD1[0]), .Z(n2511) );
  MUX2_X1 U1539 ( .A(\REGISTERS[13][15] ), .B(\REGISTERS[29][15] ), .S(
        ADD_RD1[4]), .Z(n2512) );
  MUX2_X1 U1540 ( .A(\REGISTERS[5][15] ), .B(\REGISTERS[21][15] ), .S(
        ADD_RD1[4]), .Z(n2513) );
  MUX2_X1 U1541 ( .A(n2513), .B(n2512), .S(ADD_RD1[3]), .Z(n2514) );
  MUX2_X1 U1542 ( .A(\REGISTERS[9][15] ), .B(\REGISTERS[25][15] ), .S(
        ADD_RD1[4]), .Z(n2515) );
  MUX2_X1 U1543 ( .A(\REGISTERS[1][15] ), .B(\REGISTERS[17][15] ), .S(
        ADD_RD1[4]), .Z(n2516) );
  MUX2_X1 U1544 ( .A(n2516), .B(n2515), .S(ADD_RD1[3]), .Z(n2517) );
  MUX2_X1 U1545 ( .A(n2517), .B(n2514), .S(ADD_RD1[2]), .Z(n2518) );
  MUX2_X1 U1546 ( .A(\REGISTERS[12][15] ), .B(\REGISTERS[28][15] ), .S(
        ADD_RD1[4]), .Z(n2519) );
  MUX2_X1 U1547 ( .A(\REGISTERS[4][15] ), .B(\REGISTERS[20][15] ), .S(
        ADD_RD1[4]), .Z(n2520) );
  MUX2_X1 U1548 ( .A(n2520), .B(n2519), .S(ADD_RD1[3]), .Z(n2521) );
  MUX2_X1 U1549 ( .A(\REGISTERS[8][15] ), .B(\REGISTERS[24][15] ), .S(
        ADD_RD1[4]), .Z(n2522) );
  MUX2_X1 U1550 ( .A(\REGISTERS[0][15] ), .B(\REGISTERS[16][15] ), .S(
        ADD_RD1[4]), .Z(n2523) );
  MUX2_X1 U1551 ( .A(n2523), .B(n2522), .S(ADD_RD1[3]), .Z(n2524) );
  MUX2_X1 U1552 ( .A(n2524), .B(n2521), .S(ADD_RD1[2]), .Z(n2525) );
  MUX2_X1 U1553 ( .A(n2525), .B(n2518), .S(ADD_RD1[0]), .Z(n2526) );
  MUX2_X1 U1554 ( .A(n2526), .B(n2511), .S(ADD_RD1[1]), .Z(N394) );
  MUX2_X1 U1555 ( .A(\REGISTERS[15][16] ), .B(\REGISTERS[31][16] ), .S(
        ADD_RD1[4]), .Z(n2527) );
  MUX2_X1 U1556 ( .A(\REGISTERS[7][16] ), .B(\REGISTERS[23][16] ), .S(
        ADD_RD1[4]), .Z(n2528) );
  MUX2_X1 U1557 ( .A(n2528), .B(n2527), .S(ADD_RD1[3]), .Z(n2529) );
  MUX2_X1 U1558 ( .A(\REGISTERS[11][16] ), .B(\REGISTERS[27][16] ), .S(
        ADD_RD1[4]), .Z(n2530) );
  MUX2_X1 U1559 ( .A(\REGISTERS[3][16] ), .B(\REGISTERS[19][16] ), .S(
        ADD_RD1[4]), .Z(n2531) );
  MUX2_X1 U1560 ( .A(n2531), .B(n2530), .S(ADD_RD1[3]), .Z(n2532) );
  MUX2_X1 U1561 ( .A(n2532), .B(n2529), .S(ADD_RD1[2]), .Z(n2533) );
  MUX2_X1 U1562 ( .A(\REGISTERS[14][16] ), .B(\REGISTERS[30][16] ), .S(
        ADD_RD1[4]), .Z(n2534) );
  MUX2_X1 U1563 ( .A(\REGISTERS[6][16] ), .B(\REGISTERS[22][16] ), .S(
        ADD_RD1[4]), .Z(n2535) );
  MUX2_X1 U1564 ( .A(n2535), .B(n2534), .S(ADD_RD1[3]), .Z(n2536) );
  MUX2_X1 U1565 ( .A(\REGISTERS[10][16] ), .B(\REGISTERS[26][16] ), .S(
        ADD_RD1[4]), .Z(n2537) );
  MUX2_X1 U1566 ( .A(\REGISTERS[2][16] ), .B(\REGISTERS[18][16] ), .S(
        ADD_RD1[4]), .Z(n2538) );
  MUX2_X1 U1567 ( .A(n2538), .B(n2537), .S(ADD_RD1[3]), .Z(n2539) );
  MUX2_X1 U1568 ( .A(n2539), .B(n2536), .S(ADD_RD1[2]), .Z(n2540) );
  MUX2_X1 U1569 ( .A(n2540), .B(n2533), .S(ADD_RD1[0]), .Z(n2541) );
  MUX2_X1 U1570 ( .A(\REGISTERS[13][16] ), .B(\REGISTERS[29][16] ), .S(
        ADD_RD1[4]), .Z(n2542) );
  MUX2_X1 U1571 ( .A(\REGISTERS[5][16] ), .B(\REGISTERS[21][16] ), .S(
        ADD_RD1[4]), .Z(n2543) );
  MUX2_X1 U1572 ( .A(n2543), .B(n2542), .S(ADD_RD1[3]), .Z(n2544) );
  MUX2_X1 U1573 ( .A(\REGISTERS[9][16] ), .B(\REGISTERS[25][16] ), .S(
        ADD_RD1[4]), .Z(n2545) );
  MUX2_X1 U1574 ( .A(\REGISTERS[1][16] ), .B(\REGISTERS[17][16] ), .S(
        ADD_RD1[4]), .Z(n2546) );
  MUX2_X1 U1575 ( .A(n2546), .B(n2545), .S(ADD_RD1[3]), .Z(n2547) );
  MUX2_X1 U1576 ( .A(n2547), .B(n2544), .S(ADD_RD1[2]), .Z(n2548) );
  MUX2_X1 U1577 ( .A(\REGISTERS[12][16] ), .B(\REGISTERS[28][16] ), .S(
        ADD_RD1[4]), .Z(n2549) );
  MUX2_X1 U1578 ( .A(\REGISTERS[4][16] ), .B(\REGISTERS[20][16] ), .S(
        ADD_RD1[4]), .Z(n2550) );
  MUX2_X1 U1579 ( .A(n2550), .B(n2549), .S(ADD_RD1[3]), .Z(n2551) );
  MUX2_X1 U1580 ( .A(\REGISTERS[8][16] ), .B(\REGISTERS[24][16] ), .S(
        ADD_RD1[4]), .Z(n2552) );
  MUX2_X1 U1581 ( .A(\REGISTERS[0][16] ), .B(\REGISTERS[16][16] ), .S(
        ADD_RD1[4]), .Z(n2553) );
  MUX2_X1 U1582 ( .A(n2553), .B(n2552), .S(ADD_RD1[3]), .Z(n2554) );
  MUX2_X1 U1583 ( .A(n2554), .B(n2551), .S(ADD_RD1[2]), .Z(n2555) );
  MUX2_X1 U1584 ( .A(n2555), .B(n2548), .S(ADD_RD1[0]), .Z(n2556) );
  MUX2_X1 U1585 ( .A(n2556), .B(n2541), .S(ADD_RD1[1]), .Z(N395) );
  MUX2_X1 U1586 ( .A(\REGISTERS[15][17] ), .B(\REGISTERS[31][17] ), .S(
        ADD_RD1[4]), .Z(n2557) );
  MUX2_X1 U1587 ( .A(\REGISTERS[7][17] ), .B(\REGISTERS[23][17] ), .S(
        ADD_RD1[4]), .Z(n2558) );
  MUX2_X1 U1588 ( .A(n2558), .B(n2557), .S(ADD_RD1[3]), .Z(n2559) );
  MUX2_X1 U1589 ( .A(\REGISTERS[11][17] ), .B(\REGISTERS[27][17] ), .S(
        ADD_RD1[4]), .Z(n2560) );
  MUX2_X1 U1590 ( .A(\REGISTERS[3][17] ), .B(\REGISTERS[19][17] ), .S(
        ADD_RD1[4]), .Z(n2561) );
  MUX2_X1 U1591 ( .A(n2561), .B(n2560), .S(ADD_RD1[3]), .Z(n2562) );
  MUX2_X1 U1592 ( .A(n2562), .B(n2559), .S(ADD_RD1[2]), .Z(n2563) );
  MUX2_X1 U1593 ( .A(\REGISTERS[14][17] ), .B(\REGISTERS[30][17] ), .S(
        ADD_RD1[4]), .Z(n2564) );
  MUX2_X1 U1594 ( .A(\REGISTERS[6][17] ), .B(\REGISTERS[22][17] ), .S(
        ADD_RD1[4]), .Z(n2565) );
  MUX2_X1 U1595 ( .A(n2565), .B(n2564), .S(ADD_RD1[3]), .Z(n2566) );
  MUX2_X1 U1596 ( .A(\REGISTERS[10][17] ), .B(\REGISTERS[26][17] ), .S(
        ADD_RD1[4]), .Z(n2567) );
  MUX2_X1 U1597 ( .A(\REGISTERS[2][17] ), .B(\REGISTERS[18][17] ), .S(
        ADD_RD1[4]), .Z(n2568) );
  MUX2_X1 U1598 ( .A(n2568), .B(n2567), .S(ADD_RD1[3]), .Z(n2569) );
  MUX2_X1 U1599 ( .A(n2569), .B(n2566), .S(ADD_RD1[2]), .Z(n2570) );
  MUX2_X1 U1600 ( .A(n2570), .B(n2563), .S(ADD_RD1[0]), .Z(n2571) );
  MUX2_X1 U1601 ( .A(\REGISTERS[13][17] ), .B(\REGISTERS[29][17] ), .S(
        ADD_RD1[4]), .Z(n2572) );
  MUX2_X1 U1602 ( .A(\REGISTERS[5][17] ), .B(\REGISTERS[21][17] ), .S(
        ADD_RD1[4]), .Z(n2573) );
  MUX2_X1 U1603 ( .A(n2573), .B(n2572), .S(ADD_RD1[3]), .Z(n2574) );
  MUX2_X1 U1604 ( .A(\REGISTERS[9][17] ), .B(\REGISTERS[25][17] ), .S(
        ADD_RD1[4]), .Z(n2575) );
  MUX2_X1 U1605 ( .A(\REGISTERS[1][17] ), .B(\REGISTERS[17][17] ), .S(
        ADD_RD1[4]), .Z(n2576) );
  MUX2_X1 U1606 ( .A(n2576), .B(n2575), .S(ADD_RD1[3]), .Z(n2577) );
  MUX2_X1 U1607 ( .A(n2577), .B(n2574), .S(ADD_RD1[2]), .Z(n2578) );
  MUX2_X1 U1608 ( .A(\REGISTERS[12][17] ), .B(\REGISTERS[28][17] ), .S(
        ADD_RD1[4]), .Z(n2579) );
  MUX2_X1 U1609 ( .A(\REGISTERS[4][17] ), .B(\REGISTERS[20][17] ), .S(
        ADD_RD1[4]), .Z(n2580) );
  MUX2_X1 U1610 ( .A(n2580), .B(n2579), .S(ADD_RD1[3]), .Z(n2581) );
  MUX2_X1 U1611 ( .A(\REGISTERS[8][17] ), .B(\REGISTERS[24][17] ), .S(
        ADD_RD1[4]), .Z(n2582) );
  MUX2_X1 U1612 ( .A(\REGISTERS[0][17] ), .B(\REGISTERS[16][17] ), .S(
        ADD_RD1[4]), .Z(n2583) );
  MUX2_X1 U1613 ( .A(n2583), .B(n2582), .S(ADD_RD1[3]), .Z(n2584) );
  MUX2_X1 U1614 ( .A(n2584), .B(n2581), .S(ADD_RD1[2]), .Z(n2585) );
  MUX2_X1 U1615 ( .A(n2585), .B(n2578), .S(ADD_RD1[0]), .Z(n2586) );
  MUX2_X1 U1616 ( .A(n2586), .B(n2571), .S(ADD_RD1[1]), .Z(N396) );
  MUX2_X1 U1617 ( .A(\REGISTERS[15][18] ), .B(\REGISTERS[31][18] ), .S(
        ADD_RD1[4]), .Z(n2587) );
  MUX2_X1 U1618 ( .A(\REGISTERS[7][18] ), .B(\REGISTERS[23][18] ), .S(
        ADD_RD1[4]), .Z(n2588) );
  MUX2_X1 U1619 ( .A(n2588), .B(n2587), .S(ADD_RD1[3]), .Z(n2589) );
  MUX2_X1 U1620 ( .A(\REGISTERS[11][18] ), .B(\REGISTERS[27][18] ), .S(
        ADD_RD1[4]), .Z(n2590) );
  MUX2_X1 U1621 ( .A(\REGISTERS[3][18] ), .B(\REGISTERS[19][18] ), .S(
        ADD_RD1[4]), .Z(n2591) );
  MUX2_X1 U1622 ( .A(n2591), .B(n2590), .S(ADD_RD1[3]), .Z(n2592) );
  MUX2_X1 U1623 ( .A(n2592), .B(n2589), .S(ADD_RD1[2]), .Z(n2593) );
  MUX2_X1 U1624 ( .A(\REGISTERS[14][18] ), .B(\REGISTERS[30][18] ), .S(
        ADD_RD1[4]), .Z(n2594) );
  MUX2_X1 U1625 ( .A(\REGISTERS[6][18] ), .B(\REGISTERS[22][18] ), .S(
        ADD_RD1[4]), .Z(n2595) );
  MUX2_X1 U1626 ( .A(n2595), .B(n2594), .S(ADD_RD1[3]), .Z(n2596) );
  MUX2_X1 U1627 ( .A(\REGISTERS[10][18] ), .B(\REGISTERS[26][18] ), .S(
        ADD_RD1[4]), .Z(n2597) );
  MUX2_X1 U1628 ( .A(\REGISTERS[2][18] ), .B(\REGISTERS[18][18] ), .S(
        ADD_RD1[4]), .Z(n2598) );
  MUX2_X1 U1629 ( .A(n2598), .B(n2597), .S(ADD_RD1[3]), .Z(n2599) );
  MUX2_X1 U1630 ( .A(n2599), .B(n2596), .S(ADD_RD1[2]), .Z(n2600) );
  MUX2_X1 U1631 ( .A(n2600), .B(n2593), .S(ADD_RD1[0]), .Z(n2601) );
  MUX2_X1 U1632 ( .A(\REGISTERS[13][18] ), .B(\REGISTERS[29][18] ), .S(
        ADD_RD1[4]), .Z(n2602) );
  MUX2_X1 U1633 ( .A(\REGISTERS[5][18] ), .B(\REGISTERS[21][18] ), .S(
        ADD_RD1[4]), .Z(n2603) );
  MUX2_X1 U1634 ( .A(n2603), .B(n2602), .S(ADD_RD1[3]), .Z(n2604) );
  MUX2_X1 U1635 ( .A(\REGISTERS[9][18] ), .B(\REGISTERS[25][18] ), .S(
        ADD_RD1[4]), .Z(n2605) );
  MUX2_X1 U1636 ( .A(\REGISTERS[1][18] ), .B(\REGISTERS[17][18] ), .S(
        ADD_RD1[4]), .Z(n2606) );
  MUX2_X1 U1637 ( .A(n2606), .B(n2605), .S(ADD_RD1[3]), .Z(n2607) );
  MUX2_X1 U1638 ( .A(n2607), .B(n2604), .S(ADD_RD1[2]), .Z(n2608) );
  MUX2_X1 U1639 ( .A(\REGISTERS[12][18] ), .B(\REGISTERS[28][18] ), .S(
        ADD_RD1[4]), .Z(n2609) );
  MUX2_X1 U1640 ( .A(\REGISTERS[4][18] ), .B(\REGISTERS[20][18] ), .S(
        ADD_RD1[4]), .Z(n2610) );
  MUX2_X1 U1641 ( .A(n2610), .B(n2609), .S(ADD_RD1[3]), .Z(n2611) );
  MUX2_X1 U1642 ( .A(\REGISTERS[8][18] ), .B(\REGISTERS[24][18] ), .S(
        ADD_RD1[4]), .Z(n2612) );
  MUX2_X1 U1643 ( .A(\REGISTERS[0][18] ), .B(\REGISTERS[16][18] ), .S(
        ADD_RD1[4]), .Z(n2613) );
  MUX2_X1 U1644 ( .A(n2613), .B(n2612), .S(ADD_RD1[3]), .Z(n2614) );
  MUX2_X1 U1645 ( .A(n2614), .B(n2611), .S(ADD_RD1[2]), .Z(n2615) );
  MUX2_X1 U1646 ( .A(n2615), .B(n2608), .S(ADD_RD1[0]), .Z(n2616) );
  MUX2_X1 U1647 ( .A(n2616), .B(n2601), .S(ADD_RD1[1]), .Z(N397) );
  MUX2_X1 U1648 ( .A(\REGISTERS[15][19] ), .B(\REGISTERS[31][19] ), .S(
        ADD_RD1[4]), .Z(n2617) );
  MUX2_X1 U1649 ( .A(\REGISTERS[7][19] ), .B(\REGISTERS[23][19] ), .S(
        ADD_RD1[4]), .Z(n2618) );
  MUX2_X1 U1650 ( .A(n2618), .B(n2617), .S(ADD_RD1[3]), .Z(n2619) );
  MUX2_X1 U1651 ( .A(\REGISTERS[11][19] ), .B(\REGISTERS[27][19] ), .S(
        ADD_RD1[4]), .Z(n2620) );
  MUX2_X1 U1652 ( .A(\REGISTERS[3][19] ), .B(\REGISTERS[19][19] ), .S(
        ADD_RD1[4]), .Z(n2621) );
  MUX2_X1 U1653 ( .A(n2621), .B(n2620), .S(ADD_RD1[3]), .Z(n2622) );
  MUX2_X1 U1654 ( .A(n2622), .B(n2619), .S(ADD_RD1[2]), .Z(n2623) );
  MUX2_X1 U1655 ( .A(\REGISTERS[14][19] ), .B(\REGISTERS[30][19] ), .S(
        ADD_RD1[4]), .Z(n2624) );
  MUX2_X1 U1656 ( .A(\REGISTERS[6][19] ), .B(\REGISTERS[22][19] ), .S(
        ADD_RD1[4]), .Z(n2625) );
  MUX2_X1 U1657 ( .A(n2625), .B(n2624), .S(ADD_RD1[3]), .Z(n2626) );
  MUX2_X1 U1658 ( .A(\REGISTERS[10][19] ), .B(\REGISTERS[26][19] ), .S(
        ADD_RD1[4]), .Z(n2627) );
  MUX2_X1 U1659 ( .A(\REGISTERS[2][19] ), .B(\REGISTERS[18][19] ), .S(
        ADD_RD1[4]), .Z(n2628) );
  MUX2_X1 U1660 ( .A(n2628), .B(n2627), .S(ADD_RD1[3]), .Z(n2629) );
  MUX2_X1 U1661 ( .A(n2629), .B(n2626), .S(ADD_RD1[2]), .Z(n2630) );
  MUX2_X1 U1662 ( .A(n2630), .B(n2623), .S(ADD_RD1[0]), .Z(n2631) );
  MUX2_X1 U1663 ( .A(\REGISTERS[13][19] ), .B(\REGISTERS[29][19] ), .S(
        ADD_RD1[4]), .Z(n2632) );
  MUX2_X1 U1664 ( .A(\REGISTERS[5][19] ), .B(\REGISTERS[21][19] ), .S(
        ADD_RD1[4]), .Z(n2633) );
  MUX2_X1 U1665 ( .A(n2633), .B(n2632), .S(ADD_RD1[3]), .Z(n2634) );
  MUX2_X1 U1666 ( .A(\REGISTERS[9][19] ), .B(\REGISTERS[25][19] ), .S(
        ADD_RD1[4]), .Z(n2635) );
  MUX2_X1 U1667 ( .A(\REGISTERS[1][19] ), .B(\REGISTERS[17][19] ), .S(
        ADD_RD1[4]), .Z(n2636) );
  MUX2_X1 U1668 ( .A(n2636), .B(n2635), .S(ADD_RD1[3]), .Z(n2637) );
  MUX2_X1 U1669 ( .A(n2637), .B(n2634), .S(ADD_RD1[2]), .Z(n2638) );
  MUX2_X1 U1670 ( .A(\REGISTERS[12][19] ), .B(\REGISTERS[28][19] ), .S(
        ADD_RD1[4]), .Z(n2639) );
  MUX2_X1 U1671 ( .A(\REGISTERS[4][19] ), .B(\REGISTERS[20][19] ), .S(
        ADD_RD1[4]), .Z(n2640) );
  MUX2_X1 U1672 ( .A(n2640), .B(n2639), .S(ADD_RD1[3]), .Z(n2641) );
  MUX2_X1 U1673 ( .A(\REGISTERS[8][19] ), .B(\REGISTERS[24][19] ), .S(
        ADD_RD1[4]), .Z(n2642) );
  MUX2_X1 U1674 ( .A(\REGISTERS[0][19] ), .B(\REGISTERS[16][19] ), .S(
        ADD_RD1[4]), .Z(n2643) );
  MUX2_X1 U1675 ( .A(n2643), .B(n2642), .S(ADD_RD1[3]), .Z(n2644) );
  MUX2_X1 U1676 ( .A(n2644), .B(n2641), .S(ADD_RD1[2]), .Z(n2645) );
  MUX2_X1 U1677 ( .A(n2645), .B(n2638), .S(ADD_RD1[0]), .Z(n2646) );
  MUX2_X1 U1678 ( .A(n2646), .B(n2631), .S(ADD_RD1[1]), .Z(N398) );
  MUX2_X1 U1679 ( .A(\REGISTERS[15][20] ), .B(\REGISTERS[31][20] ), .S(
        ADD_RD1[4]), .Z(n2647) );
  MUX2_X1 U1680 ( .A(\REGISTERS[7][20] ), .B(\REGISTERS[23][20] ), .S(
        ADD_RD1[4]), .Z(n2648) );
  MUX2_X1 U1681 ( .A(n2648), .B(n2647), .S(ADD_RD1[3]), .Z(n2649) );
  MUX2_X1 U1682 ( .A(\REGISTERS[11][20] ), .B(\REGISTERS[27][20] ), .S(
        ADD_RD1[4]), .Z(n2650) );
  MUX2_X1 U1683 ( .A(\REGISTERS[3][20] ), .B(\REGISTERS[19][20] ), .S(
        ADD_RD1[4]), .Z(n2651) );
  MUX2_X1 U1684 ( .A(n2651), .B(n2650), .S(ADD_RD1[3]), .Z(n2652) );
  MUX2_X1 U1685 ( .A(n2652), .B(n2649), .S(ADD_RD1[2]), .Z(n2653) );
  MUX2_X1 U1686 ( .A(\REGISTERS[14][20] ), .B(\REGISTERS[30][20] ), .S(
        ADD_RD1[4]), .Z(n2654) );
  MUX2_X1 U1687 ( .A(\REGISTERS[6][20] ), .B(\REGISTERS[22][20] ), .S(
        ADD_RD1[4]), .Z(n2655) );
  MUX2_X1 U1688 ( .A(n2655), .B(n2654), .S(ADD_RD1[3]), .Z(n2656) );
  MUX2_X1 U1689 ( .A(\REGISTERS[10][20] ), .B(\REGISTERS[26][20] ), .S(
        ADD_RD1[4]), .Z(n2657) );
  MUX2_X1 U1690 ( .A(\REGISTERS[2][20] ), .B(\REGISTERS[18][20] ), .S(
        ADD_RD1[4]), .Z(n2658) );
  MUX2_X1 U1691 ( .A(n2658), .B(n2657), .S(ADD_RD1[3]), .Z(n2659) );
  MUX2_X1 U1692 ( .A(n2659), .B(n2656), .S(ADD_RD1[2]), .Z(n2660) );
  MUX2_X1 U1693 ( .A(n2660), .B(n2653), .S(ADD_RD1[0]), .Z(n2661) );
  MUX2_X1 U1694 ( .A(\REGISTERS[13][20] ), .B(\REGISTERS[29][20] ), .S(
        ADD_RD1[4]), .Z(n2662) );
  MUX2_X1 U1695 ( .A(\REGISTERS[5][20] ), .B(\REGISTERS[21][20] ), .S(
        ADD_RD1[4]), .Z(n2663) );
  MUX2_X1 U1696 ( .A(n2663), .B(n2662), .S(ADD_RD1[3]), .Z(n2664) );
  MUX2_X1 U1697 ( .A(\REGISTERS[9][20] ), .B(\REGISTERS[25][20] ), .S(
        ADD_RD1[4]), .Z(n2665) );
  MUX2_X1 U1698 ( .A(\REGISTERS[1][20] ), .B(\REGISTERS[17][20] ), .S(
        ADD_RD1[4]), .Z(n2666) );
  MUX2_X1 U1699 ( .A(n2666), .B(n2665), .S(ADD_RD1[3]), .Z(n2667) );
  MUX2_X1 U1700 ( .A(n2667), .B(n2664), .S(ADD_RD1[2]), .Z(n2668) );
  MUX2_X1 U1701 ( .A(\REGISTERS[12][20] ), .B(\REGISTERS[28][20] ), .S(
        ADD_RD1[4]), .Z(n2669) );
  MUX2_X1 U1702 ( .A(\REGISTERS[4][20] ), .B(\REGISTERS[20][20] ), .S(
        ADD_RD1[4]), .Z(n2670) );
  MUX2_X1 U1703 ( .A(n2670), .B(n2669), .S(ADD_RD1[3]), .Z(n2671) );
  MUX2_X1 U1704 ( .A(\REGISTERS[8][20] ), .B(\REGISTERS[24][20] ), .S(
        ADD_RD1[4]), .Z(n2672) );
  MUX2_X1 U1705 ( .A(\REGISTERS[0][20] ), .B(\REGISTERS[16][20] ), .S(
        ADD_RD1[4]), .Z(n2673) );
  MUX2_X1 U1706 ( .A(n2673), .B(n2672), .S(ADD_RD1[3]), .Z(n2674) );
  MUX2_X1 U1707 ( .A(n2674), .B(n2671), .S(ADD_RD1[2]), .Z(n2675) );
  MUX2_X1 U1708 ( .A(n2675), .B(n2668), .S(ADD_RD1[0]), .Z(n2676) );
  MUX2_X1 U1709 ( .A(n2676), .B(n2661), .S(ADD_RD1[1]), .Z(N399) );
  MUX2_X1 U1710 ( .A(\REGISTERS[15][21] ), .B(\REGISTERS[31][21] ), .S(
        ADD_RD1[4]), .Z(n2677) );
  MUX2_X1 U1711 ( .A(\REGISTERS[7][21] ), .B(\REGISTERS[23][21] ), .S(
        ADD_RD1[4]), .Z(n2678) );
  MUX2_X1 U1712 ( .A(n2678), .B(n2677), .S(ADD_RD1[3]), .Z(n2679) );
  MUX2_X1 U1713 ( .A(\REGISTERS[11][21] ), .B(\REGISTERS[27][21] ), .S(
        ADD_RD1[4]), .Z(n2680) );
  MUX2_X1 U1714 ( .A(\REGISTERS[3][21] ), .B(\REGISTERS[19][21] ), .S(
        ADD_RD1[4]), .Z(n2681) );
  MUX2_X1 U1715 ( .A(n2681), .B(n2680), .S(ADD_RD1[3]), .Z(n2682) );
  MUX2_X1 U1716 ( .A(n2682), .B(n2679), .S(ADD_RD1[2]), .Z(n2683) );
  MUX2_X1 U1717 ( .A(\REGISTERS[14][21] ), .B(\REGISTERS[30][21] ), .S(
        ADD_RD1[4]), .Z(n2684) );
  MUX2_X1 U1718 ( .A(\REGISTERS[6][21] ), .B(\REGISTERS[22][21] ), .S(
        ADD_RD1[4]), .Z(n2685) );
  MUX2_X1 U1719 ( .A(n2685), .B(n2684), .S(ADD_RD1[3]), .Z(n2686) );
  MUX2_X1 U1720 ( .A(\REGISTERS[10][21] ), .B(\REGISTERS[26][21] ), .S(
        ADD_RD1[4]), .Z(n2687) );
  MUX2_X1 U1721 ( .A(\REGISTERS[2][21] ), .B(\REGISTERS[18][21] ), .S(
        ADD_RD1[4]), .Z(n2688) );
  MUX2_X1 U1722 ( .A(n2688), .B(n2687), .S(ADD_RD1[3]), .Z(n2689) );
  MUX2_X1 U1723 ( .A(n2689), .B(n2686), .S(ADD_RD1[2]), .Z(n2690) );
  MUX2_X1 U1724 ( .A(n2690), .B(n2683), .S(ADD_RD1[0]), .Z(n2691) );
  MUX2_X1 U1725 ( .A(\REGISTERS[13][21] ), .B(\REGISTERS[29][21] ), .S(
        ADD_RD1[4]), .Z(n2692) );
  MUX2_X1 U1726 ( .A(\REGISTERS[5][21] ), .B(\REGISTERS[21][21] ), .S(
        ADD_RD1[4]), .Z(n2693) );
  MUX2_X1 U1727 ( .A(n2693), .B(n2692), .S(ADD_RD1[3]), .Z(n2694) );
  MUX2_X1 U1728 ( .A(\REGISTERS[9][21] ), .B(\REGISTERS[25][21] ), .S(
        ADD_RD1[4]), .Z(n2695) );
  MUX2_X1 U1729 ( .A(\REGISTERS[1][21] ), .B(\REGISTERS[17][21] ), .S(
        ADD_RD1[4]), .Z(n2696) );
  MUX2_X1 U1730 ( .A(n2696), .B(n2695), .S(ADD_RD1[3]), .Z(n2697) );
  MUX2_X1 U1731 ( .A(n2697), .B(n2694), .S(ADD_RD1[2]), .Z(n2698) );
  MUX2_X1 U1732 ( .A(\REGISTERS[12][21] ), .B(\REGISTERS[28][21] ), .S(
        ADD_RD1[4]), .Z(n2699) );
  MUX2_X1 U1733 ( .A(\REGISTERS[4][21] ), .B(\REGISTERS[20][21] ), .S(
        ADD_RD1[4]), .Z(n2700) );
  MUX2_X1 U1734 ( .A(n2700), .B(n2699), .S(ADD_RD1[3]), .Z(n2701) );
  MUX2_X1 U1735 ( .A(\REGISTERS[8][21] ), .B(\REGISTERS[24][21] ), .S(
        ADD_RD1[4]), .Z(n2702) );
  MUX2_X1 U1736 ( .A(\REGISTERS[0][21] ), .B(\REGISTERS[16][21] ), .S(
        ADD_RD1[4]), .Z(n2703) );
  MUX2_X1 U1737 ( .A(n2703), .B(n2702), .S(ADD_RD1[3]), .Z(n2704) );
  MUX2_X1 U1738 ( .A(n2704), .B(n2701), .S(ADD_RD1[2]), .Z(n2705) );
  MUX2_X1 U1739 ( .A(n2705), .B(n2698), .S(ADD_RD1[0]), .Z(n2706) );
  MUX2_X1 U1740 ( .A(n2706), .B(n2691), .S(ADD_RD1[1]), .Z(N400) );
  MUX2_X1 U1741 ( .A(\REGISTERS[15][22] ), .B(\REGISTERS[31][22] ), .S(
        ADD_RD1[4]), .Z(n2707) );
  MUX2_X1 U1742 ( .A(\REGISTERS[7][22] ), .B(\REGISTERS[23][22] ), .S(
        ADD_RD1[4]), .Z(n2708) );
  MUX2_X1 U1743 ( .A(n2708), .B(n2707), .S(ADD_RD1[3]), .Z(n2709) );
  MUX2_X1 U1744 ( .A(\REGISTERS[11][22] ), .B(\REGISTERS[27][22] ), .S(
        ADD_RD1[4]), .Z(n2710) );
  MUX2_X1 U1745 ( .A(\REGISTERS[3][22] ), .B(\REGISTERS[19][22] ), .S(
        ADD_RD1[4]), .Z(n2711) );
  MUX2_X1 U1746 ( .A(n2711), .B(n2710), .S(ADD_RD1[3]), .Z(n2712) );
  MUX2_X1 U1747 ( .A(n2712), .B(n2709), .S(ADD_RD1[2]), .Z(n2713) );
  MUX2_X1 U1748 ( .A(\REGISTERS[14][22] ), .B(\REGISTERS[30][22] ), .S(
        ADD_RD1[4]), .Z(n2714) );
  MUX2_X1 U1749 ( .A(\REGISTERS[6][22] ), .B(\REGISTERS[22][22] ), .S(
        ADD_RD1[4]), .Z(n2715) );
  MUX2_X1 U1750 ( .A(n2715), .B(n2714), .S(ADD_RD1[3]), .Z(n2716) );
  MUX2_X1 U1751 ( .A(\REGISTERS[10][22] ), .B(\REGISTERS[26][22] ), .S(
        ADD_RD1[4]), .Z(n2717) );
  MUX2_X1 U1752 ( .A(\REGISTERS[2][22] ), .B(\REGISTERS[18][22] ), .S(
        ADD_RD1[4]), .Z(n2718) );
  MUX2_X1 U1753 ( .A(n2718), .B(n2717), .S(ADD_RD1[3]), .Z(n2719) );
  MUX2_X1 U1754 ( .A(n2719), .B(n2716), .S(ADD_RD1[2]), .Z(n2720) );
  MUX2_X1 U1755 ( .A(n2720), .B(n2713), .S(ADD_RD1[0]), .Z(n2721) );
  MUX2_X1 U1756 ( .A(\REGISTERS[13][22] ), .B(\REGISTERS[29][22] ), .S(
        ADD_RD1[4]), .Z(n2722) );
  MUX2_X1 U1757 ( .A(\REGISTERS[5][22] ), .B(\REGISTERS[21][22] ), .S(
        ADD_RD1[4]), .Z(n2723) );
  MUX2_X1 U1758 ( .A(n2723), .B(n2722), .S(ADD_RD1[3]), .Z(n2724) );
  MUX2_X1 U1759 ( .A(\REGISTERS[9][22] ), .B(\REGISTERS[25][22] ), .S(
        ADD_RD1[4]), .Z(n2725) );
  MUX2_X1 U1760 ( .A(\REGISTERS[1][22] ), .B(\REGISTERS[17][22] ), .S(
        ADD_RD1[4]), .Z(n2726) );
  MUX2_X1 U1761 ( .A(n2726), .B(n2725), .S(ADD_RD1[3]), .Z(n2727) );
  MUX2_X1 U1762 ( .A(n2727), .B(n2724), .S(ADD_RD1[2]), .Z(n2728) );
  MUX2_X1 U1763 ( .A(\REGISTERS[12][22] ), .B(\REGISTERS[28][22] ), .S(
        ADD_RD1[4]), .Z(n2729) );
  MUX2_X1 U1764 ( .A(\REGISTERS[4][22] ), .B(\REGISTERS[20][22] ), .S(
        ADD_RD1[4]), .Z(n2730) );
  MUX2_X1 U1765 ( .A(n2730), .B(n2729), .S(ADD_RD1[3]), .Z(n2731) );
  MUX2_X1 U1766 ( .A(\REGISTERS[8][22] ), .B(\REGISTERS[24][22] ), .S(
        ADD_RD1[4]), .Z(n2732) );
  MUX2_X1 U1767 ( .A(\REGISTERS[0][22] ), .B(\REGISTERS[16][22] ), .S(
        ADD_RD1[4]), .Z(n2733) );
  MUX2_X1 U1768 ( .A(n2733), .B(n2732), .S(ADD_RD1[3]), .Z(n2734) );
  MUX2_X1 U1769 ( .A(n2734), .B(n2731), .S(ADD_RD1[2]), .Z(n2735) );
  MUX2_X1 U1770 ( .A(n2735), .B(n2728), .S(ADD_RD1[0]), .Z(n2736) );
  MUX2_X1 U1771 ( .A(n2736), .B(n2721), .S(ADD_RD1[1]), .Z(N401) );
  MUX2_X1 U1772 ( .A(\REGISTERS[15][23] ), .B(\REGISTERS[31][23] ), .S(
        ADD_RD1[4]), .Z(n2737) );
  MUX2_X1 U1773 ( .A(\REGISTERS[7][23] ), .B(\REGISTERS[23][23] ), .S(
        ADD_RD1[4]), .Z(n2738) );
  MUX2_X1 U1774 ( .A(n2738), .B(n2737), .S(ADD_RD1[3]), .Z(n2739) );
  MUX2_X1 U1775 ( .A(\REGISTERS[11][23] ), .B(\REGISTERS[27][23] ), .S(
        ADD_RD1[4]), .Z(n2740) );
  MUX2_X1 U1776 ( .A(\REGISTERS[3][23] ), .B(\REGISTERS[19][23] ), .S(
        ADD_RD1[4]), .Z(n2741) );
  MUX2_X1 U1777 ( .A(n2741), .B(n2740), .S(ADD_RD1[3]), .Z(n2742) );
  MUX2_X1 U1778 ( .A(n2742), .B(n2739), .S(ADD_RD1[2]), .Z(n2743) );
  MUX2_X1 U1779 ( .A(\REGISTERS[14][23] ), .B(\REGISTERS[30][23] ), .S(
        ADD_RD1[4]), .Z(n2744) );
  MUX2_X1 U1780 ( .A(\REGISTERS[6][23] ), .B(\REGISTERS[22][23] ), .S(
        ADD_RD1[4]), .Z(n2745) );
  MUX2_X1 U1781 ( .A(n2745), .B(n2744), .S(ADD_RD1[3]), .Z(n2746) );
  MUX2_X1 U1782 ( .A(\REGISTERS[10][23] ), .B(\REGISTERS[26][23] ), .S(
        ADD_RD1[4]), .Z(n2747) );
  MUX2_X1 U1783 ( .A(\REGISTERS[2][23] ), .B(\REGISTERS[18][23] ), .S(
        ADD_RD1[4]), .Z(n2748) );
  MUX2_X1 U1784 ( .A(n2748), .B(n2747), .S(ADD_RD1[3]), .Z(n2749) );
  MUX2_X1 U1785 ( .A(n2749), .B(n2746), .S(ADD_RD1[2]), .Z(n2750) );
  MUX2_X1 U1786 ( .A(n2750), .B(n2743), .S(ADD_RD1[0]), .Z(n2751) );
  MUX2_X1 U1787 ( .A(\REGISTERS[13][23] ), .B(\REGISTERS[29][23] ), .S(
        ADD_RD1[4]), .Z(n2752) );
  MUX2_X1 U1788 ( .A(\REGISTERS[5][23] ), .B(\REGISTERS[21][23] ), .S(
        ADD_RD1[4]), .Z(n2753) );
  MUX2_X1 U1789 ( .A(n2753), .B(n2752), .S(ADD_RD1[3]), .Z(n2754) );
  MUX2_X1 U1790 ( .A(\REGISTERS[9][23] ), .B(\REGISTERS[25][23] ), .S(
        ADD_RD1[4]), .Z(n2755) );
  MUX2_X1 U1791 ( .A(\REGISTERS[1][23] ), .B(\REGISTERS[17][23] ), .S(
        ADD_RD1[4]), .Z(n2756) );
  MUX2_X1 U1792 ( .A(n2756), .B(n2755), .S(ADD_RD1[3]), .Z(n2757) );
  MUX2_X1 U1793 ( .A(n2757), .B(n2754), .S(ADD_RD1[2]), .Z(n2758) );
  MUX2_X1 U1794 ( .A(\REGISTERS[12][23] ), .B(\REGISTERS[28][23] ), .S(
        ADD_RD1[4]), .Z(n2759) );
  MUX2_X1 U1795 ( .A(\REGISTERS[4][23] ), .B(\REGISTERS[20][23] ), .S(
        ADD_RD1[4]), .Z(n2760) );
  MUX2_X1 U1796 ( .A(n2760), .B(n2759), .S(ADD_RD1[3]), .Z(n2761) );
  MUX2_X1 U1797 ( .A(\REGISTERS[8][23] ), .B(\REGISTERS[24][23] ), .S(
        ADD_RD1[4]), .Z(n2762) );
  MUX2_X1 U1798 ( .A(\REGISTERS[0][23] ), .B(\REGISTERS[16][23] ), .S(
        ADD_RD1[4]), .Z(n2763) );
  MUX2_X1 U1799 ( .A(n2763), .B(n2762), .S(ADD_RD1[3]), .Z(n2764) );
  MUX2_X1 U1800 ( .A(n2764), .B(n2761), .S(ADD_RD1[2]), .Z(n2765) );
  MUX2_X1 U1801 ( .A(n2765), .B(n2758), .S(ADD_RD1[0]), .Z(n2766) );
  MUX2_X1 U1802 ( .A(n2766), .B(n2751), .S(ADD_RD1[1]), .Z(N402) );
  MUX2_X1 U1803 ( .A(\REGISTERS[15][24] ), .B(\REGISTERS[31][24] ), .S(
        ADD_RD1[4]), .Z(n2767) );
  MUX2_X1 U1804 ( .A(\REGISTERS[7][24] ), .B(\REGISTERS[23][24] ), .S(
        ADD_RD1[4]), .Z(n2768) );
  MUX2_X1 U1805 ( .A(n2768), .B(n2767), .S(ADD_RD1[3]), .Z(n2769) );
  MUX2_X1 U1806 ( .A(\REGISTERS[11][24] ), .B(\REGISTERS[27][24] ), .S(
        ADD_RD1[4]), .Z(n2770) );
  MUX2_X1 U1807 ( .A(\REGISTERS[3][24] ), .B(\REGISTERS[19][24] ), .S(
        ADD_RD1[4]), .Z(n2771) );
  MUX2_X1 U1808 ( .A(n2771), .B(n2770), .S(ADD_RD1[3]), .Z(n2772) );
  MUX2_X1 U1809 ( .A(n2772), .B(n2769), .S(ADD_RD1[2]), .Z(n2773) );
  MUX2_X1 U1810 ( .A(\REGISTERS[14][24] ), .B(\REGISTERS[30][24] ), .S(
        ADD_RD1[4]), .Z(n2774) );
  MUX2_X1 U1811 ( .A(\REGISTERS[6][24] ), .B(\REGISTERS[22][24] ), .S(
        ADD_RD1[4]), .Z(n2775) );
  MUX2_X1 U1812 ( .A(n2775), .B(n2774), .S(ADD_RD1[3]), .Z(n2776) );
  MUX2_X1 U1813 ( .A(\REGISTERS[10][24] ), .B(\REGISTERS[26][24] ), .S(
        ADD_RD1[4]), .Z(n2777) );
  MUX2_X1 U1814 ( .A(\REGISTERS[2][24] ), .B(\REGISTERS[18][24] ), .S(
        ADD_RD1[4]), .Z(n2778) );
  MUX2_X1 U1815 ( .A(n2778), .B(n2777), .S(ADD_RD1[3]), .Z(n2779) );
  MUX2_X1 U1816 ( .A(n2779), .B(n2776), .S(ADD_RD1[2]), .Z(n2780) );
  MUX2_X1 U1817 ( .A(n2780), .B(n2773), .S(ADD_RD1[0]), .Z(n2781) );
  MUX2_X1 U1818 ( .A(\REGISTERS[13][24] ), .B(\REGISTERS[29][24] ), .S(
        ADD_RD1[4]), .Z(n2782) );
  MUX2_X1 U1819 ( .A(\REGISTERS[5][24] ), .B(\REGISTERS[21][24] ), .S(
        ADD_RD1[4]), .Z(n2783) );
  MUX2_X1 U1820 ( .A(n2783), .B(n2782), .S(ADD_RD1[3]), .Z(n2784) );
  MUX2_X1 U1821 ( .A(\REGISTERS[9][24] ), .B(\REGISTERS[25][24] ), .S(
        ADD_RD1[4]), .Z(n2785) );
  MUX2_X1 U1822 ( .A(\REGISTERS[1][24] ), .B(\REGISTERS[17][24] ), .S(
        ADD_RD1[4]), .Z(n2786) );
  MUX2_X1 U1823 ( .A(n2786), .B(n2785), .S(ADD_RD1[3]), .Z(n2787) );
  MUX2_X1 U1824 ( .A(n2787), .B(n2784), .S(ADD_RD1[2]), .Z(n2788) );
  MUX2_X1 U1825 ( .A(\REGISTERS[12][24] ), .B(\REGISTERS[28][24] ), .S(
        ADD_RD1[4]), .Z(n2789) );
  MUX2_X1 U1826 ( .A(\REGISTERS[4][24] ), .B(\REGISTERS[20][24] ), .S(
        ADD_RD1[4]), .Z(n2790) );
  MUX2_X1 U1827 ( .A(n2790), .B(n2789), .S(ADD_RD1[3]), .Z(n2791) );
  MUX2_X1 U1828 ( .A(\REGISTERS[8][24] ), .B(\REGISTERS[24][24] ), .S(
        ADD_RD1[4]), .Z(n2792) );
  MUX2_X1 U1829 ( .A(\REGISTERS[0][24] ), .B(\REGISTERS[16][24] ), .S(
        ADD_RD1[4]), .Z(n2793) );
  MUX2_X1 U1830 ( .A(n2793), .B(n2792), .S(ADD_RD1[3]), .Z(n2794) );
  MUX2_X1 U1831 ( .A(n2794), .B(n2791), .S(ADD_RD1[2]), .Z(n2795) );
  MUX2_X1 U1832 ( .A(n2795), .B(n2788), .S(ADD_RD1[0]), .Z(n2796) );
  MUX2_X1 U1833 ( .A(n2796), .B(n2781), .S(ADD_RD1[1]), .Z(N403) );
  MUX2_X1 U1834 ( .A(\REGISTERS[15][25] ), .B(\REGISTERS[31][25] ), .S(
        ADD_RD1[4]), .Z(n2797) );
  MUX2_X1 U1835 ( .A(\REGISTERS[7][25] ), .B(\REGISTERS[23][25] ), .S(
        ADD_RD1[4]), .Z(n2798) );
  MUX2_X1 U1836 ( .A(n2798), .B(n2797), .S(ADD_RD1[3]), .Z(n2799) );
  MUX2_X1 U1837 ( .A(\REGISTERS[11][25] ), .B(\REGISTERS[27][25] ), .S(
        ADD_RD1[4]), .Z(n2800) );
  MUX2_X1 U1838 ( .A(\REGISTERS[3][25] ), .B(\REGISTERS[19][25] ), .S(
        ADD_RD1[4]), .Z(n2801) );
  MUX2_X1 U1839 ( .A(n2801), .B(n2800), .S(ADD_RD1[3]), .Z(n2802) );
  MUX2_X1 U1840 ( .A(n2802), .B(n2799), .S(ADD_RD1[2]), .Z(n2803) );
  MUX2_X1 U1841 ( .A(\REGISTERS[14][25] ), .B(\REGISTERS[30][25] ), .S(
        ADD_RD1[4]), .Z(n2804) );
  MUX2_X1 U1842 ( .A(\REGISTERS[6][25] ), .B(\REGISTERS[22][25] ), .S(
        ADD_RD1[4]), .Z(n2805) );
  MUX2_X1 U1843 ( .A(n2805), .B(n2804), .S(ADD_RD1[3]), .Z(n2806) );
  MUX2_X1 U1844 ( .A(\REGISTERS[10][25] ), .B(\REGISTERS[26][25] ), .S(
        ADD_RD1[4]), .Z(n2807) );
  MUX2_X1 U1845 ( .A(\REGISTERS[2][25] ), .B(\REGISTERS[18][25] ), .S(
        ADD_RD1[4]), .Z(n2808) );
  MUX2_X1 U1846 ( .A(n2808), .B(n2807), .S(ADD_RD1[3]), .Z(n2809) );
  MUX2_X1 U1847 ( .A(n2809), .B(n2806), .S(ADD_RD1[2]), .Z(n2810) );
  MUX2_X1 U1848 ( .A(n2810), .B(n2803), .S(ADD_RD1[0]), .Z(n2811) );
  MUX2_X1 U1849 ( .A(\REGISTERS[13][25] ), .B(\REGISTERS[29][25] ), .S(
        ADD_RD1[4]), .Z(n2812) );
  MUX2_X1 U1850 ( .A(\REGISTERS[5][25] ), .B(\REGISTERS[21][25] ), .S(
        ADD_RD1[4]), .Z(n2813) );
  MUX2_X1 U1851 ( .A(n2813), .B(n2812), .S(ADD_RD1[3]), .Z(n2814) );
  MUX2_X1 U1852 ( .A(\REGISTERS[9][25] ), .B(\REGISTERS[25][25] ), .S(
        ADD_RD1[4]), .Z(n2815) );
  MUX2_X1 U1853 ( .A(\REGISTERS[1][25] ), .B(\REGISTERS[17][25] ), .S(
        ADD_RD1[4]), .Z(n2816) );
  MUX2_X1 U1854 ( .A(n2816), .B(n2815), .S(ADD_RD1[3]), .Z(n2817) );
  MUX2_X1 U1855 ( .A(n2817), .B(n2814), .S(ADD_RD1[2]), .Z(n2818) );
  MUX2_X1 U1856 ( .A(\REGISTERS[12][25] ), .B(\REGISTERS[28][25] ), .S(
        ADD_RD1[4]), .Z(n2819) );
  MUX2_X1 U1857 ( .A(\REGISTERS[4][25] ), .B(\REGISTERS[20][25] ), .S(
        ADD_RD1[4]), .Z(n2820) );
  MUX2_X1 U1858 ( .A(n2820), .B(n2819), .S(ADD_RD1[3]), .Z(n2821) );
  MUX2_X1 U1859 ( .A(\REGISTERS[8][25] ), .B(\REGISTERS[24][25] ), .S(
        ADD_RD1[4]), .Z(n2822) );
  MUX2_X1 U1860 ( .A(\REGISTERS[0][25] ), .B(\REGISTERS[16][25] ), .S(
        ADD_RD1[4]), .Z(n2823) );
  MUX2_X1 U1861 ( .A(n2823), .B(n2822), .S(ADD_RD1[3]), .Z(n2824) );
  MUX2_X1 U1862 ( .A(n2824), .B(n2821), .S(ADD_RD1[2]), .Z(n2825) );
  MUX2_X1 U1863 ( .A(n2825), .B(n2818), .S(ADD_RD1[0]), .Z(n2826) );
  MUX2_X1 U1864 ( .A(n2826), .B(n2811), .S(ADD_RD1[1]), .Z(N404) );
  MUX2_X1 U1865 ( .A(\REGISTERS[15][26] ), .B(\REGISTERS[31][26] ), .S(
        ADD_RD1[4]), .Z(n2827) );
  MUX2_X1 U1866 ( .A(\REGISTERS[7][26] ), .B(\REGISTERS[23][26] ), .S(
        ADD_RD1[4]), .Z(n2828) );
  MUX2_X1 U1867 ( .A(n2828), .B(n2827), .S(ADD_RD1[3]), .Z(n2829) );
  MUX2_X1 U1868 ( .A(\REGISTERS[11][26] ), .B(\REGISTERS[27][26] ), .S(
        ADD_RD1[4]), .Z(n2830) );
  MUX2_X1 U1869 ( .A(\REGISTERS[3][26] ), .B(\REGISTERS[19][26] ), .S(
        ADD_RD1[4]), .Z(n2831) );
  MUX2_X1 U1870 ( .A(n2831), .B(n2830), .S(ADD_RD1[3]), .Z(n2832) );
  MUX2_X1 U1871 ( .A(n2832), .B(n2829), .S(ADD_RD1[2]), .Z(n2833) );
  MUX2_X1 U1872 ( .A(\REGISTERS[14][26] ), .B(\REGISTERS[30][26] ), .S(
        ADD_RD1[4]), .Z(n2834) );
  MUX2_X1 U1873 ( .A(\REGISTERS[6][26] ), .B(\REGISTERS[22][26] ), .S(
        ADD_RD1[4]), .Z(n2835) );
  MUX2_X1 U1874 ( .A(n2835), .B(n2834), .S(ADD_RD1[3]), .Z(n2836) );
  MUX2_X1 U1875 ( .A(\REGISTERS[10][26] ), .B(\REGISTERS[26][26] ), .S(
        ADD_RD1[4]), .Z(n2837) );
  MUX2_X1 U1876 ( .A(\REGISTERS[2][26] ), .B(\REGISTERS[18][26] ), .S(
        ADD_RD1[4]), .Z(n2838) );
  MUX2_X1 U1877 ( .A(n2838), .B(n2837), .S(ADD_RD1[3]), .Z(n2839) );
  MUX2_X1 U1878 ( .A(n2839), .B(n2836), .S(ADD_RD1[2]), .Z(n2840) );
  MUX2_X1 U1879 ( .A(n2840), .B(n2833), .S(ADD_RD1[0]), .Z(n2841) );
  MUX2_X1 U1880 ( .A(\REGISTERS[13][26] ), .B(\REGISTERS[29][26] ), .S(
        ADD_RD1[4]), .Z(n2842) );
  MUX2_X1 U1881 ( .A(\REGISTERS[5][26] ), .B(\REGISTERS[21][26] ), .S(
        ADD_RD1[4]), .Z(n2843) );
  MUX2_X1 U1882 ( .A(n2843), .B(n2842), .S(ADD_RD1[3]), .Z(n2844) );
  MUX2_X1 U1883 ( .A(\REGISTERS[9][26] ), .B(\REGISTERS[25][26] ), .S(
        ADD_RD1[4]), .Z(n2845) );
  MUX2_X1 U1884 ( .A(\REGISTERS[1][26] ), .B(\REGISTERS[17][26] ), .S(
        ADD_RD1[4]), .Z(n2846) );
  MUX2_X1 U1885 ( .A(n2846), .B(n2845), .S(ADD_RD1[3]), .Z(n2847) );
  MUX2_X1 U1886 ( .A(n2847), .B(n2844), .S(ADD_RD1[2]), .Z(n2848) );
  MUX2_X1 U1887 ( .A(\REGISTERS[12][26] ), .B(\REGISTERS[28][26] ), .S(
        ADD_RD1[4]), .Z(n2849) );
  MUX2_X1 U1888 ( .A(\REGISTERS[4][26] ), .B(\REGISTERS[20][26] ), .S(
        ADD_RD1[4]), .Z(n2850) );
  MUX2_X1 U1889 ( .A(n2850), .B(n2849), .S(ADD_RD1[3]), .Z(n2851) );
  MUX2_X1 U1890 ( .A(\REGISTERS[8][26] ), .B(\REGISTERS[24][26] ), .S(
        ADD_RD1[4]), .Z(n2852) );
  MUX2_X1 U1891 ( .A(\REGISTERS[0][26] ), .B(\REGISTERS[16][26] ), .S(
        ADD_RD1[4]), .Z(n2853) );
  MUX2_X1 U1892 ( .A(n2853), .B(n2852), .S(ADD_RD1[3]), .Z(n2854) );
  MUX2_X1 U1893 ( .A(n2854), .B(n2851), .S(ADD_RD1[2]), .Z(n2855) );
  MUX2_X1 U1894 ( .A(n2855), .B(n2848), .S(ADD_RD1[0]), .Z(n2856) );
  MUX2_X1 U1895 ( .A(n2856), .B(n2841), .S(ADD_RD1[1]), .Z(N405) );
  MUX2_X1 U1896 ( .A(\REGISTERS[15][27] ), .B(\REGISTERS[31][27] ), .S(
        ADD_RD1[4]), .Z(n2857) );
  MUX2_X1 U1897 ( .A(\REGISTERS[7][27] ), .B(\REGISTERS[23][27] ), .S(
        ADD_RD1[4]), .Z(n2858) );
  MUX2_X1 U1898 ( .A(n2858), .B(n2857), .S(ADD_RD1[3]), .Z(n2859) );
  MUX2_X1 U1899 ( .A(\REGISTERS[11][27] ), .B(\REGISTERS[27][27] ), .S(
        ADD_RD1[4]), .Z(n2860) );
  MUX2_X1 U1900 ( .A(\REGISTERS[3][27] ), .B(\REGISTERS[19][27] ), .S(
        ADD_RD1[4]), .Z(n2861) );
  MUX2_X1 U1901 ( .A(n2861), .B(n2860), .S(ADD_RD1[3]), .Z(n2862) );
  MUX2_X1 U1902 ( .A(n2862), .B(n2859), .S(ADD_RD1[2]), .Z(n2863) );
  MUX2_X1 U1903 ( .A(\REGISTERS[14][27] ), .B(\REGISTERS[30][27] ), .S(
        ADD_RD1[4]), .Z(n2864) );
  MUX2_X1 U1904 ( .A(\REGISTERS[6][27] ), .B(\REGISTERS[22][27] ), .S(
        ADD_RD1[4]), .Z(n2865) );
  MUX2_X1 U1905 ( .A(n2865), .B(n2864), .S(ADD_RD1[3]), .Z(n2866) );
  MUX2_X1 U1906 ( .A(\REGISTERS[10][27] ), .B(\REGISTERS[26][27] ), .S(
        ADD_RD1[4]), .Z(n2867) );
  MUX2_X1 U1907 ( .A(\REGISTERS[2][27] ), .B(\REGISTERS[18][27] ), .S(
        ADD_RD1[4]), .Z(n2868) );
  MUX2_X1 U1908 ( .A(n2868), .B(n2867), .S(ADD_RD1[3]), .Z(n2869) );
  MUX2_X1 U1909 ( .A(n2869), .B(n2866), .S(ADD_RD1[2]), .Z(n2870) );
  MUX2_X1 U1910 ( .A(n2870), .B(n2863), .S(ADD_RD1[0]), .Z(n2871) );
  MUX2_X1 U1911 ( .A(\REGISTERS[13][27] ), .B(\REGISTERS[29][27] ), .S(
        ADD_RD1[4]), .Z(n2872) );
  MUX2_X1 U1912 ( .A(\REGISTERS[5][27] ), .B(\REGISTERS[21][27] ), .S(
        ADD_RD1[4]), .Z(n2873) );
  MUX2_X1 U1913 ( .A(n2873), .B(n2872), .S(ADD_RD1[3]), .Z(n2874) );
  MUX2_X1 U1914 ( .A(\REGISTERS[9][27] ), .B(\REGISTERS[25][27] ), .S(
        ADD_RD1[4]), .Z(n2875) );
  MUX2_X1 U1915 ( .A(\REGISTERS[1][27] ), .B(\REGISTERS[17][27] ), .S(
        ADD_RD1[4]), .Z(n2876) );
  MUX2_X1 U1916 ( .A(n2876), .B(n2875), .S(ADD_RD1[3]), .Z(n2877) );
  MUX2_X1 U1917 ( .A(n2877), .B(n2874), .S(ADD_RD1[2]), .Z(n2878) );
  MUX2_X1 U1918 ( .A(\REGISTERS[12][27] ), .B(\REGISTERS[28][27] ), .S(
        ADD_RD1[4]), .Z(n2879) );
  MUX2_X1 U1919 ( .A(\REGISTERS[4][27] ), .B(\REGISTERS[20][27] ), .S(
        ADD_RD1[4]), .Z(n2880) );
  MUX2_X1 U1920 ( .A(n2880), .B(n2879), .S(ADD_RD1[3]), .Z(n2881) );
  MUX2_X1 U1921 ( .A(\REGISTERS[8][27] ), .B(\REGISTERS[24][27] ), .S(
        ADD_RD1[4]), .Z(n2882) );
  MUX2_X1 U1922 ( .A(\REGISTERS[0][27] ), .B(\REGISTERS[16][27] ), .S(
        ADD_RD1[4]), .Z(n2883) );
  MUX2_X1 U1923 ( .A(n2883), .B(n2882), .S(ADD_RD1[3]), .Z(n2884) );
  MUX2_X1 U1924 ( .A(n2884), .B(n2881), .S(ADD_RD1[2]), .Z(n2885) );
  MUX2_X1 U1925 ( .A(n2885), .B(n2878), .S(ADD_RD1[0]), .Z(n2886) );
  MUX2_X1 U1926 ( .A(n2886), .B(n2871), .S(ADD_RD1[1]), .Z(N406) );
  MUX2_X1 U1927 ( .A(\REGISTERS[15][28] ), .B(\REGISTERS[31][28] ), .S(
        ADD_RD1[4]), .Z(n2887) );
  MUX2_X1 U1928 ( .A(\REGISTERS[7][28] ), .B(\REGISTERS[23][28] ), .S(
        ADD_RD1[4]), .Z(n2888) );
  MUX2_X1 U1929 ( .A(n2888), .B(n2887), .S(ADD_RD1[3]), .Z(n2889) );
  MUX2_X1 U1930 ( .A(\REGISTERS[11][28] ), .B(\REGISTERS[27][28] ), .S(
        ADD_RD1[4]), .Z(n2890) );
  MUX2_X1 U1931 ( .A(\REGISTERS[3][28] ), .B(\REGISTERS[19][28] ), .S(
        ADD_RD1[4]), .Z(n2891) );
  MUX2_X1 U1932 ( .A(n2891), .B(n2890), .S(ADD_RD1[3]), .Z(n2892) );
  MUX2_X1 U1933 ( .A(n2892), .B(n2889), .S(ADD_RD1[2]), .Z(n2893) );
  MUX2_X1 U1934 ( .A(\REGISTERS[14][28] ), .B(\REGISTERS[30][28] ), .S(
        ADD_RD1[4]), .Z(n2894) );
  MUX2_X1 U1935 ( .A(\REGISTERS[6][28] ), .B(\REGISTERS[22][28] ), .S(
        ADD_RD1[4]), .Z(n2895) );
  MUX2_X1 U1936 ( .A(n2895), .B(n2894), .S(ADD_RD1[3]), .Z(n2896) );
  MUX2_X1 U1937 ( .A(\REGISTERS[10][28] ), .B(\REGISTERS[26][28] ), .S(
        ADD_RD1[4]), .Z(n2897) );
  MUX2_X1 U1938 ( .A(\REGISTERS[2][28] ), .B(\REGISTERS[18][28] ), .S(
        ADD_RD1[4]), .Z(n2898) );
  MUX2_X1 U1939 ( .A(n2898), .B(n2897), .S(ADD_RD1[3]), .Z(n2899) );
  MUX2_X1 U1940 ( .A(n2899), .B(n2896), .S(ADD_RD1[2]), .Z(n2900) );
  MUX2_X1 U1941 ( .A(n2900), .B(n2893), .S(ADD_RD1[0]), .Z(n2901) );
  MUX2_X1 U1942 ( .A(\REGISTERS[13][28] ), .B(\REGISTERS[29][28] ), .S(
        ADD_RD1[4]), .Z(n2902) );
  MUX2_X1 U1943 ( .A(\REGISTERS[5][28] ), .B(\REGISTERS[21][28] ), .S(
        ADD_RD1[4]), .Z(n2903) );
  MUX2_X1 U1944 ( .A(n2903), .B(n2902), .S(ADD_RD1[3]), .Z(n2904) );
  MUX2_X1 U1945 ( .A(\REGISTERS[9][28] ), .B(\REGISTERS[25][28] ), .S(
        ADD_RD1[4]), .Z(n2905) );
  MUX2_X1 U1946 ( .A(\REGISTERS[1][28] ), .B(\REGISTERS[17][28] ), .S(
        ADD_RD1[4]), .Z(n2906) );
  MUX2_X1 U1947 ( .A(n2906), .B(n2905), .S(ADD_RD1[3]), .Z(n2907) );
  MUX2_X1 U1948 ( .A(n2907), .B(n2904), .S(ADD_RD1[2]), .Z(n2908) );
  MUX2_X1 U1949 ( .A(\REGISTERS[12][28] ), .B(\REGISTERS[28][28] ), .S(
        ADD_RD1[4]), .Z(n2909) );
  MUX2_X1 U1950 ( .A(\REGISTERS[4][28] ), .B(\REGISTERS[20][28] ), .S(
        ADD_RD1[4]), .Z(n2910) );
  MUX2_X1 U1951 ( .A(n2910), .B(n2909), .S(ADD_RD1[3]), .Z(n2911) );
  MUX2_X1 U1952 ( .A(\REGISTERS[8][28] ), .B(\REGISTERS[24][28] ), .S(
        ADD_RD1[4]), .Z(n2912) );
  MUX2_X1 U1953 ( .A(\REGISTERS[0][28] ), .B(\REGISTERS[16][28] ), .S(
        ADD_RD1[4]), .Z(n2913) );
  MUX2_X1 U1954 ( .A(n2913), .B(n2912), .S(ADD_RD1[3]), .Z(n2914) );
  MUX2_X1 U1955 ( .A(n2914), .B(n2911), .S(ADD_RD1[2]), .Z(n2915) );
  MUX2_X1 U1956 ( .A(n2915), .B(n2908), .S(ADD_RD1[0]), .Z(n2916) );
  MUX2_X1 U1957 ( .A(n2916), .B(n2901), .S(ADD_RD1[1]), .Z(N407) );
  MUX2_X1 U1958 ( .A(\REGISTERS[15][29] ), .B(\REGISTERS[31][29] ), .S(
        ADD_RD1[4]), .Z(n2917) );
  MUX2_X1 U1959 ( .A(\REGISTERS[7][29] ), .B(\REGISTERS[23][29] ), .S(
        ADD_RD1[4]), .Z(n2918) );
  MUX2_X1 U1960 ( .A(n2918), .B(n2917), .S(ADD_RD1[3]), .Z(n2919) );
  MUX2_X1 U1961 ( .A(\REGISTERS[11][29] ), .B(\REGISTERS[27][29] ), .S(
        ADD_RD1[4]), .Z(n2920) );
  MUX2_X1 U1962 ( .A(\REGISTERS[3][29] ), .B(\REGISTERS[19][29] ), .S(
        ADD_RD1[4]), .Z(n2921) );
  MUX2_X1 U1963 ( .A(n2921), .B(n2920), .S(ADD_RD1[3]), .Z(n2922) );
  MUX2_X1 U1964 ( .A(n2922), .B(n2919), .S(ADD_RD1[2]), .Z(n2923) );
  MUX2_X1 U1965 ( .A(\REGISTERS[14][29] ), .B(\REGISTERS[30][29] ), .S(
        ADD_RD1[4]), .Z(n2924) );
  MUX2_X1 U1966 ( .A(\REGISTERS[6][29] ), .B(\REGISTERS[22][29] ), .S(
        ADD_RD1[4]), .Z(n2925) );
  MUX2_X1 U1967 ( .A(n2925), .B(n2924), .S(ADD_RD1[3]), .Z(n2926) );
  MUX2_X1 U1968 ( .A(\REGISTERS[10][29] ), .B(\REGISTERS[26][29] ), .S(
        ADD_RD1[4]), .Z(n2927) );
  MUX2_X1 U1969 ( .A(\REGISTERS[2][29] ), .B(\REGISTERS[18][29] ), .S(
        ADD_RD1[4]), .Z(n2928) );
  MUX2_X1 U1970 ( .A(n2928), .B(n2927), .S(ADD_RD1[3]), .Z(n2929) );
  MUX2_X1 U1971 ( .A(n2929), .B(n2926), .S(ADD_RD1[2]), .Z(n2930) );
  MUX2_X1 U1972 ( .A(n2930), .B(n2923), .S(ADD_RD1[0]), .Z(n2931) );
  MUX2_X1 U1973 ( .A(\REGISTERS[13][29] ), .B(\REGISTERS[29][29] ), .S(
        ADD_RD1[4]), .Z(n2932) );
  MUX2_X1 U1974 ( .A(\REGISTERS[5][29] ), .B(\REGISTERS[21][29] ), .S(
        ADD_RD1[4]), .Z(n2933) );
  MUX2_X1 U1975 ( .A(n2933), .B(n2932), .S(ADD_RD1[3]), .Z(n2934) );
  MUX2_X1 U1976 ( .A(\REGISTERS[9][29] ), .B(\REGISTERS[25][29] ), .S(
        ADD_RD1[4]), .Z(n2935) );
  MUX2_X1 U1977 ( .A(\REGISTERS[1][29] ), .B(\REGISTERS[17][29] ), .S(
        ADD_RD1[4]), .Z(n2936) );
  MUX2_X1 U1978 ( .A(n2936), .B(n2935), .S(ADD_RD1[3]), .Z(n2937) );
  MUX2_X1 U1979 ( .A(n2937), .B(n2934), .S(ADD_RD1[2]), .Z(n2938) );
  MUX2_X1 U1980 ( .A(\REGISTERS[12][29] ), .B(\REGISTERS[28][29] ), .S(
        ADD_RD1[4]), .Z(n2939) );
  MUX2_X1 U1981 ( .A(\REGISTERS[4][29] ), .B(\REGISTERS[20][29] ), .S(
        ADD_RD1[4]), .Z(n2940) );
  MUX2_X1 U1982 ( .A(n2940), .B(n2939), .S(ADD_RD1[3]), .Z(n2941) );
  MUX2_X1 U1983 ( .A(\REGISTERS[8][29] ), .B(\REGISTERS[24][29] ), .S(
        ADD_RD1[4]), .Z(n2942) );
  MUX2_X1 U1984 ( .A(\REGISTERS[0][29] ), .B(\REGISTERS[16][29] ), .S(
        ADD_RD1[4]), .Z(n2943) );
  MUX2_X1 U1985 ( .A(n2943), .B(n2942), .S(ADD_RD1[3]), .Z(n2944) );
  MUX2_X1 U1986 ( .A(n2944), .B(n2941), .S(ADD_RD1[2]), .Z(n2945) );
  MUX2_X1 U1987 ( .A(n2945), .B(n2938), .S(ADD_RD1[0]), .Z(n2946) );
  MUX2_X1 U1988 ( .A(n2946), .B(n2931), .S(ADD_RD1[1]), .Z(N408) );
  MUX2_X1 U1989 ( .A(\REGISTERS[15][30] ), .B(\REGISTERS[31][30] ), .S(
        ADD_RD1[4]), .Z(n2947) );
  MUX2_X1 U1990 ( .A(\REGISTERS[7][30] ), .B(\REGISTERS[23][30] ), .S(
        ADD_RD1[4]), .Z(n2948) );
  MUX2_X1 U1991 ( .A(n2948), .B(n2947), .S(ADD_RD1[3]), .Z(n2949) );
  MUX2_X1 U1992 ( .A(\REGISTERS[11][30] ), .B(\REGISTERS[27][30] ), .S(
        ADD_RD1[4]), .Z(n2950) );
  MUX2_X1 U1993 ( .A(\REGISTERS[3][30] ), .B(\REGISTERS[19][30] ), .S(
        ADD_RD1[4]), .Z(n2951) );
  MUX2_X1 U1994 ( .A(n2951), .B(n2950), .S(ADD_RD1[3]), .Z(n2952) );
  MUX2_X1 U1995 ( .A(n2952), .B(n2949), .S(ADD_RD1[2]), .Z(n2953) );
  MUX2_X1 U1996 ( .A(\REGISTERS[14][30] ), .B(\REGISTERS[30][30] ), .S(
        ADD_RD1[4]), .Z(n2954) );
  MUX2_X1 U1997 ( .A(\REGISTERS[6][30] ), .B(\REGISTERS[22][30] ), .S(
        ADD_RD1[4]), .Z(n2955) );
  MUX2_X1 U1998 ( .A(n2955), .B(n2954), .S(ADD_RD1[3]), .Z(n2956) );
  MUX2_X1 U1999 ( .A(\REGISTERS[10][30] ), .B(\REGISTERS[26][30] ), .S(
        ADD_RD1[4]), .Z(n2957) );
  MUX2_X1 U2000 ( .A(\REGISTERS[2][30] ), .B(\REGISTERS[18][30] ), .S(
        ADD_RD1[4]), .Z(n2958) );
  MUX2_X1 U2001 ( .A(n2958), .B(n2957), .S(ADD_RD1[3]), .Z(n2959) );
  MUX2_X1 U2002 ( .A(n2959), .B(n2956), .S(ADD_RD1[2]), .Z(n2960) );
  MUX2_X1 U2003 ( .A(n2960), .B(n2953), .S(ADD_RD1[0]), .Z(n2961) );
  MUX2_X1 U2004 ( .A(\REGISTERS[13][30] ), .B(\REGISTERS[29][30] ), .S(
        ADD_RD1[4]), .Z(n2962) );
  MUX2_X1 U2005 ( .A(\REGISTERS[5][30] ), .B(\REGISTERS[21][30] ), .S(
        ADD_RD1[4]), .Z(n2963) );
  MUX2_X1 U2006 ( .A(n2963), .B(n2962), .S(ADD_RD1[3]), .Z(n2964) );
  MUX2_X1 U2007 ( .A(\REGISTERS[9][30] ), .B(\REGISTERS[25][30] ), .S(
        ADD_RD1[4]), .Z(n2965) );
  MUX2_X1 U2008 ( .A(\REGISTERS[1][30] ), .B(\REGISTERS[17][30] ), .S(
        ADD_RD1[4]), .Z(n2966) );
  MUX2_X1 U2009 ( .A(n2966), .B(n2965), .S(ADD_RD1[3]), .Z(n2967) );
  MUX2_X1 U2010 ( .A(n2967), .B(n2964), .S(ADD_RD1[2]), .Z(n2968) );
  MUX2_X1 U2011 ( .A(\REGISTERS[12][30] ), .B(\REGISTERS[28][30] ), .S(
        ADD_RD1[4]), .Z(n2969) );
  MUX2_X1 U2012 ( .A(\REGISTERS[4][30] ), .B(\REGISTERS[20][30] ), .S(
        ADD_RD1[4]), .Z(n2970) );
  MUX2_X1 U2013 ( .A(n2970), .B(n2969), .S(ADD_RD1[3]), .Z(n2971) );
  MUX2_X1 U2014 ( .A(\REGISTERS[8][30] ), .B(\REGISTERS[24][30] ), .S(
        ADD_RD1[4]), .Z(n2972) );
  MUX2_X1 U2015 ( .A(\REGISTERS[0][30] ), .B(\REGISTERS[16][30] ), .S(
        ADD_RD1[4]), .Z(n2973) );
  MUX2_X1 U2016 ( .A(n2973), .B(n2972), .S(ADD_RD1[3]), .Z(n2974) );
  MUX2_X1 U2017 ( .A(n2974), .B(n2971), .S(ADD_RD1[2]), .Z(n2975) );
  MUX2_X1 U2018 ( .A(n2975), .B(n2968), .S(ADD_RD1[0]), .Z(n2976) );
  MUX2_X1 U2019 ( .A(n2976), .B(n2961), .S(ADD_RD1[1]), .Z(N409) );
  MUX2_X1 U2020 ( .A(\REGISTERS[15][31] ), .B(\REGISTERS[31][31] ), .S(
        ADD_RD1[4]), .Z(n2977) );
  MUX2_X1 U2021 ( .A(\REGISTERS[7][31] ), .B(\REGISTERS[23][31] ), .S(
        ADD_RD1[4]), .Z(n2978) );
  MUX2_X1 U2022 ( .A(n2978), .B(n2977), .S(ADD_RD1[3]), .Z(n2979) );
  MUX2_X1 U2023 ( .A(\REGISTERS[11][31] ), .B(\REGISTERS[27][31] ), .S(
        ADD_RD1[4]), .Z(n2980) );
  MUX2_X1 U2024 ( .A(\REGISTERS[3][31] ), .B(\REGISTERS[19][31] ), .S(
        ADD_RD1[4]), .Z(n2981) );
  MUX2_X1 U2025 ( .A(n2981), .B(n2980), .S(ADD_RD1[3]), .Z(n2982) );
  MUX2_X1 U2026 ( .A(n2982), .B(n2979), .S(ADD_RD1[2]), .Z(n2983) );
  MUX2_X1 U2027 ( .A(\REGISTERS[14][31] ), .B(\REGISTERS[30][31] ), .S(
        ADD_RD1[4]), .Z(n2984) );
  MUX2_X1 U2028 ( .A(\REGISTERS[6][31] ), .B(\REGISTERS[22][31] ), .S(
        ADD_RD1[4]), .Z(n2985) );
  MUX2_X1 U2029 ( .A(n2985), .B(n2984), .S(ADD_RD1[3]), .Z(n2986) );
  MUX2_X1 U2030 ( .A(\REGISTERS[10][31] ), .B(\REGISTERS[26][31] ), .S(
        ADD_RD1[4]), .Z(n2987) );
  MUX2_X1 U2031 ( .A(\REGISTERS[2][31] ), .B(\REGISTERS[18][31] ), .S(
        ADD_RD1[4]), .Z(n2988) );
  MUX2_X1 U2032 ( .A(n2988), .B(n2987), .S(ADD_RD1[3]), .Z(n2989) );
  MUX2_X1 U2033 ( .A(n2989), .B(n2986), .S(ADD_RD1[2]), .Z(n2990) );
  MUX2_X1 U2034 ( .A(n2990), .B(n2983), .S(ADD_RD1[0]), .Z(n2991) );
  MUX2_X1 U2035 ( .A(\REGISTERS[13][31] ), .B(\REGISTERS[29][31] ), .S(
        ADD_RD1[4]), .Z(n2992) );
  MUX2_X1 U2036 ( .A(\REGISTERS[5][31] ), .B(\REGISTERS[21][31] ), .S(
        ADD_RD1[4]), .Z(n2993) );
  MUX2_X1 U2037 ( .A(n2993), .B(n2992), .S(ADD_RD1[3]), .Z(n2994) );
  MUX2_X1 U2038 ( .A(\REGISTERS[9][31] ), .B(\REGISTERS[25][31] ), .S(
        ADD_RD1[4]), .Z(n2995) );
  MUX2_X1 U2039 ( .A(\REGISTERS[1][31] ), .B(\REGISTERS[17][31] ), .S(
        ADD_RD1[4]), .Z(n2996) );
  MUX2_X1 U2040 ( .A(n2996), .B(n2995), .S(ADD_RD1[3]), .Z(n2997) );
  MUX2_X1 U2041 ( .A(n2997), .B(n2994), .S(ADD_RD1[2]), .Z(n2998) );
  MUX2_X1 U2042 ( .A(\REGISTERS[12][31] ), .B(\REGISTERS[28][31] ), .S(
        ADD_RD1[4]), .Z(n2999) );
  MUX2_X1 U2043 ( .A(\REGISTERS[4][31] ), .B(\REGISTERS[20][31] ), .S(
        ADD_RD1[4]), .Z(n3000) );
  MUX2_X1 U2044 ( .A(n3000), .B(n2999), .S(ADD_RD1[3]), .Z(n3001) );
  MUX2_X1 U2045 ( .A(\REGISTERS[8][31] ), .B(\REGISTERS[24][31] ), .S(
        ADD_RD1[4]), .Z(n3002) );
  MUX2_X1 U2046 ( .A(\REGISTERS[0][31] ), .B(\REGISTERS[16][31] ), .S(
        ADD_RD1[4]), .Z(n3003) );
  MUX2_X1 U2047 ( .A(n3003), .B(n3002), .S(ADD_RD1[3]), .Z(n3004) );
  MUX2_X1 U2048 ( .A(n3004), .B(n3001), .S(ADD_RD1[2]), .Z(n3005) );
  MUX2_X1 U2049 ( .A(n3005), .B(n2998), .S(ADD_RD1[0]), .Z(n3006) );
  MUX2_X1 U2050 ( .A(n3006), .B(n2991), .S(ADD_RD1[1]), .Z(N410) );
  MUX2_X1 U2051 ( .A(\REGISTERS[0][31] ), .B(n3007), .S(n3008), .Z(n2163) );
  MUX2_X1 U2052 ( .A(\REGISTERS[0][30] ), .B(n3009), .S(n3008), .Z(n2162) );
  MUX2_X1 U2053 ( .A(\REGISTERS[0][29] ), .B(n3010), .S(n3008), .Z(n2161) );
  MUX2_X1 U2054 ( .A(\REGISTERS[0][28] ), .B(n3011), .S(n3008), .Z(n2160) );
  MUX2_X1 U2055 ( .A(\REGISTERS[0][27] ), .B(n3012), .S(n3008), .Z(n2159) );
  MUX2_X1 U2056 ( .A(\REGISTERS[0][26] ), .B(n3013), .S(n3008), .Z(n2158) );
  MUX2_X1 U2057 ( .A(\REGISTERS[0][25] ), .B(n3014), .S(n3008), .Z(n2157) );
  MUX2_X1 U2058 ( .A(\REGISTERS[0][24] ), .B(n3015), .S(n3008), .Z(n2156) );
  MUX2_X1 U2059 ( .A(\REGISTERS[0][23] ), .B(n3016), .S(n3008), .Z(n2155) );
  MUX2_X1 U2060 ( .A(\REGISTERS[0][22] ), .B(n3017), .S(n3008), .Z(n2154) );
  MUX2_X1 U2061 ( .A(\REGISTERS[0][21] ), .B(n3018), .S(n3008), .Z(n2153) );
  MUX2_X1 U2062 ( .A(\REGISTERS[0][20] ), .B(n3019), .S(n3008), .Z(n2152) );
  MUX2_X1 U2063 ( .A(\REGISTERS[0][19] ), .B(n3020), .S(n3008), .Z(n2151) );
  MUX2_X1 U2064 ( .A(\REGISTERS[0][18] ), .B(n3021), .S(n3008), .Z(n2150) );
  MUX2_X1 U2065 ( .A(\REGISTERS[0][17] ), .B(n3022), .S(n3008), .Z(n2149) );
  MUX2_X1 U2066 ( .A(\REGISTERS[0][16] ), .B(n3023), .S(n3008), .Z(n2148) );
  MUX2_X1 U2067 ( .A(\REGISTERS[0][15] ), .B(n3024), .S(n3008), .Z(n2147) );
  MUX2_X1 U2068 ( .A(\REGISTERS[0][14] ), .B(n3025), .S(n3008), .Z(n2146) );
  MUX2_X1 U2069 ( .A(\REGISTERS[0][13] ), .B(n3026), .S(n3008), .Z(n2145) );
  MUX2_X1 U2070 ( .A(\REGISTERS[0][12] ), .B(n3027), .S(n3008), .Z(n2144) );
  MUX2_X1 U2071 ( .A(\REGISTERS[0][11] ), .B(n3028), .S(n3008), .Z(n2143) );
  MUX2_X1 U2072 ( .A(\REGISTERS[0][10] ), .B(n3029), .S(n3008), .Z(n2142) );
  MUX2_X1 U2073 ( .A(\REGISTERS[0][9] ), .B(n3030), .S(n3008), .Z(n2141) );
  MUX2_X1 U2074 ( .A(\REGISTERS[0][8] ), .B(n3031), .S(n3008), .Z(n2140) );
  MUX2_X1 U2075 ( .A(\REGISTERS[0][7] ), .B(n3032), .S(n3008), .Z(n2139) );
  MUX2_X1 U2076 ( .A(\REGISTERS[0][6] ), .B(n3033), .S(n3008), .Z(n2138) );
  MUX2_X1 U2077 ( .A(\REGISTERS[0][5] ), .B(n3034), .S(n3008), .Z(n2137) );
  MUX2_X1 U2078 ( .A(\REGISTERS[0][4] ), .B(n3035), .S(n3008), .Z(n2136) );
  MUX2_X1 U2079 ( .A(\REGISTERS[0][3] ), .B(n3036), .S(n3008), .Z(n2135) );
  MUX2_X1 U2080 ( .A(\REGISTERS[0][2] ), .B(n3037), .S(n3008), .Z(n2134) );
  MUX2_X1 U2081 ( .A(\REGISTERS[0][1] ), .B(n3038), .S(n3008), .Z(n2133) );
  MUX2_X1 U2082 ( .A(\REGISTERS[0][0] ), .B(n3039), .S(n3008), .Z(n2132) );
  MUX2_X1 U2083 ( .A(\REGISTERS[1][31] ), .B(n3007), .S(n60), .Z(n2131) );
  MUX2_X1 U2084 ( .A(\REGISTERS[1][30] ), .B(n3009), .S(n60), .Z(n2130) );
  MUX2_X1 U2085 ( .A(\REGISTERS[1][29] ), .B(n3010), .S(n60), .Z(n2129) );
  MUX2_X1 U2086 ( .A(\REGISTERS[1][28] ), .B(n3011), .S(n60), .Z(n2128) );
  MUX2_X1 U2087 ( .A(\REGISTERS[1][27] ), .B(n3012), .S(n60), .Z(n2127) );
  MUX2_X1 U2088 ( .A(\REGISTERS[1][26] ), .B(n3013), .S(n60), .Z(n2126) );
  MUX2_X1 U2089 ( .A(\REGISTERS[1][25] ), .B(n3014), .S(n60), .Z(n2125) );
  MUX2_X1 U2090 ( .A(\REGISTERS[1][24] ), .B(n3015), .S(n60), .Z(n2124) );
  MUX2_X1 U2091 ( .A(\REGISTERS[1][23] ), .B(n3016), .S(n60), .Z(n2123) );
  MUX2_X1 U2092 ( .A(\REGISTERS[1][22] ), .B(n3017), .S(n60), .Z(n2122) );
  MUX2_X1 U2093 ( .A(\REGISTERS[1][21] ), .B(n3018), .S(n60), .Z(n2121) );
  MUX2_X1 U2094 ( .A(\REGISTERS[1][20] ), .B(n3019), .S(n60), .Z(n2120) );
  MUX2_X1 U2095 ( .A(\REGISTERS[1][19] ), .B(n3020), .S(n60), .Z(n2119) );
  MUX2_X1 U2096 ( .A(\REGISTERS[1][18] ), .B(n3021), .S(n60), .Z(n2118) );
  MUX2_X1 U2097 ( .A(\REGISTERS[1][17] ), .B(n3022), .S(n60), .Z(n2117) );
  MUX2_X1 U2098 ( .A(\REGISTERS[1][16] ), .B(n3023), .S(n60), .Z(n2116) );
  MUX2_X1 U2099 ( .A(\REGISTERS[1][15] ), .B(n3024), .S(n60), .Z(n2115) );
  MUX2_X1 U2100 ( .A(\REGISTERS[1][14] ), .B(n3025), .S(n60), .Z(n2114) );
  MUX2_X1 U2101 ( .A(\REGISTERS[1][13] ), .B(n3026), .S(n60), .Z(n2113) );
  MUX2_X1 U2102 ( .A(\REGISTERS[1][12] ), .B(n3027), .S(n60), .Z(n2112) );
  MUX2_X1 U2103 ( .A(\REGISTERS[1][11] ), .B(n3028), .S(n60), .Z(n2111) );
  MUX2_X1 U2104 ( .A(\REGISTERS[1][10] ), .B(n3029), .S(n60), .Z(n2110) );
  MUX2_X1 U2105 ( .A(\REGISTERS[1][9] ), .B(n3030), .S(n60), .Z(n2109) );
  MUX2_X1 U2106 ( .A(\REGISTERS[1][8] ), .B(n3031), .S(n60), .Z(n2108) );
  MUX2_X1 U2107 ( .A(\REGISTERS[1][7] ), .B(n3032), .S(n60), .Z(n2107) );
  MUX2_X1 U2108 ( .A(\REGISTERS[1][6] ), .B(n3033), .S(n60), .Z(n2106) );
  MUX2_X1 U2109 ( .A(\REGISTERS[1][5] ), .B(n3034), .S(n60), .Z(n2105) );
  MUX2_X1 U2110 ( .A(\REGISTERS[1][4] ), .B(n3035), .S(n60), .Z(n2104) );
  MUX2_X1 U2111 ( .A(\REGISTERS[1][3] ), .B(n3036), .S(n60), .Z(n2103) );
  MUX2_X1 U2112 ( .A(\REGISTERS[1][2] ), .B(n3037), .S(n60), .Z(n2102) );
  MUX2_X1 U2113 ( .A(\REGISTERS[1][1] ), .B(n3038), .S(n60), .Z(n2101) );
  MUX2_X1 U2114 ( .A(\REGISTERS[1][0] ), .B(n3039), .S(n60), .Z(n2100) );
  OAI21_X1 U2115 ( .B1(n3040), .B2(n3044), .A(n3042), .ZN(n3043) );
  MUX2_X1 U2116 ( .A(\REGISTERS[2][31] ), .B(n3007), .S(n62), .Z(n2099) );
  MUX2_X1 U2117 ( .A(\REGISTERS[2][30] ), .B(n3009), .S(n62), .Z(n2098) );
  MUX2_X1 U2118 ( .A(\REGISTERS[2][29] ), .B(n3010), .S(n62), .Z(n2097) );
  MUX2_X1 U2119 ( .A(\REGISTERS[2][28] ), .B(n3011), .S(n62), .Z(n2096) );
  MUX2_X1 U2120 ( .A(\REGISTERS[2][27] ), .B(n3012), .S(n62), .Z(n2095) );
  MUX2_X1 U2121 ( .A(\REGISTERS[2][26] ), .B(n3013), .S(n62), .Z(n2094) );
  MUX2_X1 U2122 ( .A(\REGISTERS[2][25] ), .B(n3014), .S(n62), .Z(n2093) );
  MUX2_X1 U2123 ( .A(\REGISTERS[2][24] ), .B(n3015), .S(n62), .Z(n2092) );
  MUX2_X1 U2124 ( .A(\REGISTERS[2][23] ), .B(n3016), .S(n62), .Z(n2091) );
  MUX2_X1 U2125 ( .A(\REGISTERS[2][22] ), .B(n3017), .S(n62), .Z(n2090) );
  MUX2_X1 U2126 ( .A(\REGISTERS[2][21] ), .B(n3018), .S(n62), .Z(n2089) );
  MUX2_X1 U2127 ( .A(\REGISTERS[2][20] ), .B(n3019), .S(n62), .Z(n2088) );
  MUX2_X1 U2128 ( .A(\REGISTERS[2][19] ), .B(n3020), .S(n62), .Z(n2087) );
  MUX2_X1 U2129 ( .A(\REGISTERS[2][18] ), .B(n3021), .S(n62), .Z(n2086) );
  MUX2_X1 U2130 ( .A(\REGISTERS[2][17] ), .B(n3022), .S(n62), .Z(n2085) );
  MUX2_X1 U2131 ( .A(\REGISTERS[2][16] ), .B(n3023), .S(n62), .Z(n2084) );
  MUX2_X1 U2132 ( .A(\REGISTERS[2][15] ), .B(n3024), .S(n62), .Z(n2083) );
  MUX2_X1 U2133 ( .A(\REGISTERS[2][14] ), .B(n3025), .S(n62), .Z(n2082) );
  MUX2_X1 U2134 ( .A(\REGISTERS[2][13] ), .B(n3026), .S(n62), .Z(n2081) );
  MUX2_X1 U2135 ( .A(\REGISTERS[2][12] ), .B(n3027), .S(n62), .Z(n2080) );
  MUX2_X1 U2136 ( .A(\REGISTERS[2][11] ), .B(n3028), .S(n62), .Z(n2079) );
  MUX2_X1 U2137 ( .A(\REGISTERS[2][10] ), .B(n3029), .S(n62), .Z(n2078) );
  MUX2_X1 U2138 ( .A(\REGISTERS[2][9] ), .B(n3030), .S(n62), .Z(n2077) );
  MUX2_X1 U2139 ( .A(\REGISTERS[2][8] ), .B(n3031), .S(n62), .Z(n2076) );
  MUX2_X1 U2140 ( .A(\REGISTERS[2][7] ), .B(n3032), .S(n62), .Z(n2075) );
  MUX2_X1 U2141 ( .A(\REGISTERS[2][6] ), .B(n3033), .S(n62), .Z(n2074) );
  MUX2_X1 U2142 ( .A(\REGISTERS[2][5] ), .B(n3034), .S(n62), .Z(n2073) );
  MUX2_X1 U2143 ( .A(\REGISTERS[2][4] ), .B(n3035), .S(n62), .Z(n2072) );
  MUX2_X1 U2144 ( .A(\REGISTERS[2][3] ), .B(n3036), .S(n62), .Z(n2071) );
  MUX2_X1 U2145 ( .A(\REGISTERS[2][2] ), .B(n3037), .S(n62), .Z(n2070) );
  MUX2_X1 U2146 ( .A(\REGISTERS[2][1] ), .B(n3038), .S(n62), .Z(n2069) );
  MUX2_X1 U2147 ( .A(\REGISTERS[2][0] ), .B(n3039), .S(n62), .Z(n2068) );
  OAI21_X1 U2148 ( .B1(n3040), .B2(n3046), .A(n3042), .ZN(n3045) );
  MUX2_X1 U2149 ( .A(\REGISTERS[3][31] ), .B(n3007), .S(n56), .Z(n2067) );
  MUX2_X1 U2150 ( .A(\REGISTERS[3][30] ), .B(n3009), .S(n56), .Z(n2066) );
  MUX2_X1 U2151 ( .A(\REGISTERS[3][29] ), .B(n3010), .S(n56), .Z(n2065) );
  MUX2_X1 U2152 ( .A(\REGISTERS[3][28] ), .B(n3011), .S(n56), .Z(n2064) );
  MUX2_X1 U2153 ( .A(\REGISTERS[3][27] ), .B(n3012), .S(n56), .Z(n2063) );
  MUX2_X1 U2154 ( .A(\REGISTERS[3][26] ), .B(n3013), .S(n56), .Z(n2062) );
  MUX2_X1 U2155 ( .A(\REGISTERS[3][25] ), .B(n3014), .S(n56), .Z(n2061) );
  MUX2_X1 U2156 ( .A(\REGISTERS[3][24] ), .B(n3015), .S(n56), .Z(n2060) );
  MUX2_X1 U2157 ( .A(\REGISTERS[3][23] ), .B(n3016), .S(n56), .Z(n2059) );
  MUX2_X1 U2158 ( .A(\REGISTERS[3][22] ), .B(n3017), .S(n56), .Z(n2058) );
  MUX2_X1 U2159 ( .A(\REGISTERS[3][21] ), .B(n3018), .S(n56), .Z(n2057) );
  MUX2_X1 U2160 ( .A(\REGISTERS[3][20] ), .B(n3019), .S(n56), .Z(n2056) );
  MUX2_X1 U2161 ( .A(\REGISTERS[3][19] ), .B(n3020), .S(n56), .Z(n2055) );
  MUX2_X1 U2162 ( .A(\REGISTERS[3][18] ), .B(n3021), .S(n56), .Z(n2054) );
  MUX2_X1 U2163 ( .A(\REGISTERS[3][17] ), .B(n3022), .S(n56), .Z(n2053) );
  MUX2_X1 U2164 ( .A(\REGISTERS[3][16] ), .B(n3023), .S(n56), .Z(n2052) );
  MUX2_X1 U2165 ( .A(\REGISTERS[3][15] ), .B(n3024), .S(n56), .Z(n2051) );
  MUX2_X1 U2166 ( .A(\REGISTERS[3][14] ), .B(n3025), .S(n56), .Z(n2050) );
  MUX2_X1 U2167 ( .A(\REGISTERS[3][13] ), .B(n3026), .S(n56), .Z(n2049) );
  MUX2_X1 U2168 ( .A(\REGISTERS[3][12] ), .B(n3027), .S(n56), .Z(n2048) );
  MUX2_X1 U2169 ( .A(\REGISTERS[3][11] ), .B(n3028), .S(n56), .Z(n2047) );
  MUX2_X1 U2170 ( .A(\REGISTERS[3][10] ), .B(n3029), .S(n56), .Z(n2046) );
  MUX2_X1 U2171 ( .A(\REGISTERS[3][9] ), .B(n3030), .S(n56), .Z(n2045) );
  MUX2_X1 U2172 ( .A(\REGISTERS[3][8] ), .B(n3031), .S(n56), .Z(n2044) );
  MUX2_X1 U2173 ( .A(\REGISTERS[3][7] ), .B(n3032), .S(n56), .Z(n2043) );
  MUX2_X1 U2174 ( .A(\REGISTERS[3][6] ), .B(n3033), .S(n56), .Z(n2042) );
  MUX2_X1 U2175 ( .A(\REGISTERS[3][5] ), .B(n3034), .S(n56), .Z(n2041) );
  MUX2_X1 U2176 ( .A(\REGISTERS[3][4] ), .B(n3035), .S(n56), .Z(n2040) );
  MUX2_X1 U2177 ( .A(\REGISTERS[3][3] ), .B(n3036), .S(n56), .Z(n2039) );
  MUX2_X1 U2178 ( .A(\REGISTERS[3][2] ), .B(n3037), .S(n56), .Z(n2038) );
  MUX2_X1 U2179 ( .A(\REGISTERS[3][1] ), .B(n3038), .S(n56), .Z(n2037) );
  MUX2_X1 U2180 ( .A(\REGISTERS[3][0] ), .B(n3039), .S(n56), .Z(n2036) );
  OAI21_X1 U2181 ( .B1(n3040), .B2(n3048), .A(n3042), .ZN(n3047) );
  MUX2_X1 U2182 ( .A(\REGISTERS[4][31] ), .B(n3007), .S(n58), .Z(n2035) );
  MUX2_X1 U2183 ( .A(\REGISTERS[4][30] ), .B(n3009), .S(n58), .Z(n2034) );
  MUX2_X1 U2184 ( .A(\REGISTERS[4][29] ), .B(n3010), .S(n58), .Z(n2033) );
  MUX2_X1 U2185 ( .A(\REGISTERS[4][28] ), .B(n3011), .S(n58), .Z(n2032) );
  MUX2_X1 U2186 ( .A(\REGISTERS[4][27] ), .B(n3012), .S(n58), .Z(n2031) );
  MUX2_X1 U2187 ( .A(\REGISTERS[4][26] ), .B(n3013), .S(n58), .Z(n2030) );
  MUX2_X1 U2188 ( .A(\REGISTERS[4][25] ), .B(n3014), .S(n58), .Z(n2029) );
  MUX2_X1 U2189 ( .A(\REGISTERS[4][24] ), .B(n3015), .S(n58), .Z(n2028) );
  MUX2_X1 U2190 ( .A(\REGISTERS[4][23] ), .B(n3016), .S(n58), .Z(n2027) );
  MUX2_X1 U2191 ( .A(\REGISTERS[4][22] ), .B(n3017), .S(n58), .Z(n2026) );
  MUX2_X1 U2192 ( .A(\REGISTERS[4][21] ), .B(n3018), .S(n58), .Z(n2025) );
  MUX2_X1 U2193 ( .A(\REGISTERS[4][20] ), .B(n3019), .S(n58), .Z(n2024) );
  MUX2_X1 U2194 ( .A(\REGISTERS[4][19] ), .B(n3020), .S(n58), .Z(n2023) );
  MUX2_X1 U2195 ( .A(\REGISTERS[4][18] ), .B(n3021), .S(n58), .Z(n2022) );
  MUX2_X1 U2196 ( .A(\REGISTERS[4][17] ), .B(n3022), .S(n58), .Z(n2021) );
  MUX2_X1 U2197 ( .A(\REGISTERS[4][16] ), .B(n3023), .S(n58), .Z(n2020) );
  MUX2_X1 U2198 ( .A(\REGISTERS[4][15] ), .B(n3024), .S(n58), .Z(n2019) );
  MUX2_X1 U2199 ( .A(\REGISTERS[4][14] ), .B(n3025), .S(n58), .Z(n2018) );
  MUX2_X1 U2200 ( .A(\REGISTERS[4][13] ), .B(n3026), .S(n58), .Z(n2017) );
  MUX2_X1 U2201 ( .A(\REGISTERS[4][12] ), .B(n3027), .S(n58), .Z(n2016) );
  MUX2_X1 U2202 ( .A(\REGISTERS[4][11] ), .B(n3028), .S(n58), .Z(n2015) );
  MUX2_X1 U2203 ( .A(\REGISTERS[4][10] ), .B(n3029), .S(n58), .Z(n2014) );
  MUX2_X1 U2204 ( .A(\REGISTERS[4][9] ), .B(n3030), .S(n58), .Z(n2013) );
  MUX2_X1 U2205 ( .A(\REGISTERS[4][8] ), .B(n3031), .S(n58), .Z(n2012) );
  MUX2_X1 U2206 ( .A(\REGISTERS[4][7] ), .B(n3032), .S(n58), .Z(n2011) );
  MUX2_X1 U2207 ( .A(\REGISTERS[4][6] ), .B(n3033), .S(n58), .Z(n2010) );
  MUX2_X1 U2208 ( .A(\REGISTERS[4][5] ), .B(n3034), .S(n58), .Z(n2009) );
  MUX2_X1 U2209 ( .A(\REGISTERS[4][4] ), .B(n3035), .S(n58), .Z(n2008) );
  MUX2_X1 U2210 ( .A(\REGISTERS[4][3] ), .B(n3036), .S(n58), .Z(n2007) );
  MUX2_X1 U2211 ( .A(\REGISTERS[4][2] ), .B(n3037), .S(n58), .Z(n2006) );
  MUX2_X1 U2212 ( .A(\REGISTERS[4][1] ), .B(n3038), .S(n58), .Z(n2005) );
  MUX2_X1 U2213 ( .A(\REGISTERS[4][0] ), .B(n3039), .S(n58), .Z(n2004) );
  OAI21_X1 U2214 ( .B1(n3040), .B2(n3050), .A(n3042), .ZN(n3049) );
  MUX2_X1 U2215 ( .A(\REGISTERS[5][31] ), .B(n3007), .S(n52), .Z(n2003) );
  MUX2_X1 U2216 ( .A(\REGISTERS[5][30] ), .B(n3009), .S(n52), .Z(n2002) );
  MUX2_X1 U2217 ( .A(\REGISTERS[5][29] ), .B(n3010), .S(n52), .Z(n2001) );
  MUX2_X1 U2218 ( .A(\REGISTERS[5][28] ), .B(n3011), .S(n52), .Z(n2000) );
  MUX2_X1 U2219 ( .A(\REGISTERS[5][27] ), .B(n3012), .S(n52), .Z(n1999) );
  MUX2_X1 U2220 ( .A(\REGISTERS[5][26] ), .B(n3013), .S(n52), .Z(n1998) );
  MUX2_X1 U2221 ( .A(\REGISTERS[5][25] ), .B(n3014), .S(n52), .Z(n1997) );
  MUX2_X1 U2222 ( .A(\REGISTERS[5][24] ), .B(n3015), .S(n52), .Z(n1996) );
  MUX2_X1 U2223 ( .A(\REGISTERS[5][23] ), .B(n3016), .S(n52), .Z(n1995) );
  MUX2_X1 U2224 ( .A(\REGISTERS[5][22] ), .B(n3017), .S(n52), .Z(n1994) );
  MUX2_X1 U2225 ( .A(\REGISTERS[5][21] ), .B(n3018), .S(n52), .Z(n1993) );
  MUX2_X1 U2226 ( .A(\REGISTERS[5][20] ), .B(n3019), .S(n52), .Z(n1992) );
  MUX2_X1 U2227 ( .A(\REGISTERS[5][19] ), .B(n3020), .S(n52), .Z(n1991) );
  MUX2_X1 U2228 ( .A(\REGISTERS[5][18] ), .B(n3021), .S(n52), .Z(n1990) );
  MUX2_X1 U2229 ( .A(\REGISTERS[5][17] ), .B(n3022), .S(n52), .Z(n1989) );
  MUX2_X1 U2230 ( .A(\REGISTERS[5][16] ), .B(n3023), .S(n52), .Z(n1988) );
  MUX2_X1 U2231 ( .A(\REGISTERS[5][15] ), .B(n3024), .S(n52), .Z(n1987) );
  MUX2_X1 U2232 ( .A(\REGISTERS[5][14] ), .B(n3025), .S(n52), .Z(n1986) );
  MUX2_X1 U2233 ( .A(\REGISTERS[5][13] ), .B(n3026), .S(n52), .Z(n1985) );
  MUX2_X1 U2234 ( .A(\REGISTERS[5][12] ), .B(n3027), .S(n52), .Z(n1984) );
  MUX2_X1 U2235 ( .A(\REGISTERS[5][11] ), .B(n3028), .S(n52), .Z(n1983) );
  MUX2_X1 U2236 ( .A(\REGISTERS[5][10] ), .B(n3029), .S(n52), .Z(n1982) );
  MUX2_X1 U2237 ( .A(\REGISTERS[5][9] ), .B(n3030), .S(n52), .Z(n1981) );
  MUX2_X1 U2238 ( .A(\REGISTERS[5][8] ), .B(n3031), .S(n52), .Z(n1980) );
  MUX2_X1 U2239 ( .A(\REGISTERS[5][7] ), .B(n3032), .S(n52), .Z(n1979) );
  MUX2_X1 U2240 ( .A(\REGISTERS[5][6] ), .B(n3033), .S(n52), .Z(n1978) );
  MUX2_X1 U2241 ( .A(\REGISTERS[5][5] ), .B(n3034), .S(n52), .Z(n1977) );
  MUX2_X1 U2242 ( .A(\REGISTERS[5][4] ), .B(n3035), .S(n52), .Z(n1976) );
  MUX2_X1 U2243 ( .A(\REGISTERS[5][3] ), .B(n3036), .S(n52), .Z(n1975) );
  MUX2_X1 U2244 ( .A(\REGISTERS[5][2] ), .B(n3037), .S(n52), .Z(n1974) );
  MUX2_X1 U2245 ( .A(\REGISTERS[5][1] ), .B(n3038), .S(n52), .Z(n1973) );
  MUX2_X1 U2246 ( .A(\REGISTERS[5][0] ), .B(n3039), .S(n52), .Z(n1972) );
  OAI21_X1 U2247 ( .B1(n3040), .B2(n3052), .A(n3042), .ZN(n3051) );
  MUX2_X1 U2248 ( .A(\REGISTERS[6][31] ), .B(n3007), .S(n54), .Z(n1971) );
  MUX2_X1 U2249 ( .A(\REGISTERS[6][30] ), .B(n3009), .S(n54), .Z(n1970) );
  MUX2_X1 U2250 ( .A(\REGISTERS[6][29] ), .B(n3010), .S(n54), .Z(n1969) );
  MUX2_X1 U2251 ( .A(\REGISTERS[6][28] ), .B(n3011), .S(n54), .Z(n1968) );
  MUX2_X1 U2252 ( .A(\REGISTERS[6][27] ), .B(n3012), .S(n54), .Z(n1967) );
  MUX2_X1 U2253 ( .A(\REGISTERS[6][26] ), .B(n3013), .S(n54), .Z(n1966) );
  MUX2_X1 U2254 ( .A(\REGISTERS[6][25] ), .B(n3014), .S(n54), .Z(n1965) );
  MUX2_X1 U2255 ( .A(\REGISTERS[6][24] ), .B(n3015), .S(n54), .Z(n1964) );
  MUX2_X1 U2256 ( .A(\REGISTERS[6][23] ), .B(n3016), .S(n54), .Z(n1963) );
  MUX2_X1 U2257 ( .A(\REGISTERS[6][22] ), .B(n3017), .S(n54), .Z(n1962) );
  MUX2_X1 U2258 ( .A(\REGISTERS[6][21] ), .B(n3018), .S(n54), .Z(n1961) );
  MUX2_X1 U2259 ( .A(\REGISTERS[6][20] ), .B(n3019), .S(n54), .Z(n1960) );
  MUX2_X1 U2260 ( .A(\REGISTERS[6][19] ), .B(n3020), .S(n54), .Z(n1959) );
  MUX2_X1 U2261 ( .A(\REGISTERS[6][18] ), .B(n3021), .S(n54), .Z(n1958) );
  MUX2_X1 U2262 ( .A(\REGISTERS[6][17] ), .B(n3022), .S(n54), .Z(n1957) );
  MUX2_X1 U2263 ( .A(\REGISTERS[6][16] ), .B(n3023), .S(n54), .Z(n1956) );
  MUX2_X1 U2264 ( .A(\REGISTERS[6][15] ), .B(n3024), .S(n54), .Z(n1955) );
  MUX2_X1 U2265 ( .A(\REGISTERS[6][14] ), .B(n3025), .S(n54), .Z(n1954) );
  MUX2_X1 U2266 ( .A(\REGISTERS[6][13] ), .B(n3026), .S(n54), .Z(n1953) );
  MUX2_X1 U2267 ( .A(\REGISTERS[6][12] ), .B(n3027), .S(n54), .Z(n1952) );
  MUX2_X1 U2268 ( .A(\REGISTERS[6][11] ), .B(n3028), .S(n54), .Z(n1951) );
  MUX2_X1 U2269 ( .A(\REGISTERS[6][10] ), .B(n3029), .S(n54), .Z(n1950) );
  MUX2_X1 U2270 ( .A(\REGISTERS[6][9] ), .B(n3030), .S(n54), .Z(n1949) );
  MUX2_X1 U2271 ( .A(\REGISTERS[6][8] ), .B(n3031), .S(n54), .Z(n1948) );
  MUX2_X1 U2272 ( .A(\REGISTERS[6][7] ), .B(n3032), .S(n54), .Z(n1947) );
  MUX2_X1 U2273 ( .A(\REGISTERS[6][6] ), .B(n3033), .S(n54), .Z(n1946) );
  MUX2_X1 U2274 ( .A(\REGISTERS[6][5] ), .B(n3034), .S(n54), .Z(n1945) );
  MUX2_X1 U2275 ( .A(\REGISTERS[6][4] ), .B(n3035), .S(n54), .Z(n1944) );
  MUX2_X1 U2276 ( .A(\REGISTERS[6][3] ), .B(n3036), .S(n54), .Z(n1943) );
  MUX2_X1 U2277 ( .A(\REGISTERS[6][2] ), .B(n3037), .S(n54), .Z(n1942) );
  MUX2_X1 U2278 ( .A(\REGISTERS[6][1] ), .B(n3038), .S(n54), .Z(n1941) );
  MUX2_X1 U2279 ( .A(\REGISTERS[6][0] ), .B(n3039), .S(n54), .Z(n1940) );
  OAI21_X1 U2280 ( .B1(n3040), .B2(n3054), .A(n3042), .ZN(n3053) );
  MUX2_X1 U2281 ( .A(\REGISTERS[7][31] ), .B(n3007), .S(n48), .Z(n1939) );
  MUX2_X1 U2282 ( .A(\REGISTERS[7][30] ), .B(n3009), .S(n48), .Z(n1938) );
  MUX2_X1 U2283 ( .A(\REGISTERS[7][29] ), .B(n3010), .S(n48), .Z(n1937) );
  MUX2_X1 U2284 ( .A(\REGISTERS[7][28] ), .B(n3011), .S(n48), .Z(n1936) );
  MUX2_X1 U2285 ( .A(\REGISTERS[7][27] ), .B(n3012), .S(n48), .Z(n1935) );
  MUX2_X1 U2286 ( .A(\REGISTERS[7][26] ), .B(n3013), .S(n48), .Z(n1934) );
  MUX2_X1 U2287 ( .A(\REGISTERS[7][25] ), .B(n3014), .S(n48), .Z(n1933) );
  MUX2_X1 U2288 ( .A(\REGISTERS[7][24] ), .B(n3015), .S(n48), .Z(n1932) );
  MUX2_X1 U2289 ( .A(\REGISTERS[7][23] ), .B(n3016), .S(n48), .Z(n1931) );
  MUX2_X1 U2290 ( .A(\REGISTERS[7][22] ), .B(n3017), .S(n48), .Z(n1930) );
  MUX2_X1 U2291 ( .A(\REGISTERS[7][21] ), .B(n3018), .S(n48), .Z(n1929) );
  MUX2_X1 U2292 ( .A(\REGISTERS[7][20] ), .B(n3019), .S(n48), .Z(n1928) );
  MUX2_X1 U2293 ( .A(\REGISTERS[7][19] ), .B(n3020), .S(n48), .Z(n1927) );
  MUX2_X1 U2294 ( .A(\REGISTERS[7][18] ), .B(n3021), .S(n48), .Z(n1926) );
  MUX2_X1 U2295 ( .A(\REGISTERS[7][17] ), .B(n3022), .S(n48), .Z(n1925) );
  MUX2_X1 U2296 ( .A(\REGISTERS[7][16] ), .B(n3023), .S(n48), .Z(n1924) );
  MUX2_X1 U2297 ( .A(\REGISTERS[7][15] ), .B(n3024), .S(n48), .Z(n1923) );
  MUX2_X1 U2298 ( .A(\REGISTERS[7][14] ), .B(n3025), .S(n48), .Z(n1922) );
  MUX2_X1 U2299 ( .A(\REGISTERS[7][13] ), .B(n3026), .S(n48), .Z(n1921) );
  MUX2_X1 U2300 ( .A(\REGISTERS[7][12] ), .B(n3027), .S(n48), .Z(n1920) );
  MUX2_X1 U2301 ( .A(\REGISTERS[7][11] ), .B(n3028), .S(n48), .Z(n1919) );
  MUX2_X1 U2302 ( .A(\REGISTERS[7][10] ), .B(n3029), .S(n48), .Z(n1918) );
  MUX2_X1 U2303 ( .A(\REGISTERS[7][9] ), .B(n3030), .S(n48), .Z(n1917) );
  MUX2_X1 U2304 ( .A(\REGISTERS[7][8] ), .B(n3031), .S(n48), .Z(n1916) );
  MUX2_X1 U2305 ( .A(\REGISTERS[7][7] ), .B(n3032), .S(n48), .Z(n1915) );
  MUX2_X1 U2306 ( .A(\REGISTERS[7][6] ), .B(n3033), .S(n48), .Z(n1914) );
  MUX2_X1 U2307 ( .A(\REGISTERS[7][5] ), .B(n3034), .S(n48), .Z(n1913) );
  MUX2_X1 U2308 ( .A(\REGISTERS[7][4] ), .B(n3035), .S(n48), .Z(n1912) );
  MUX2_X1 U2309 ( .A(\REGISTERS[7][3] ), .B(n3036), .S(n48), .Z(n1911) );
  MUX2_X1 U2310 ( .A(\REGISTERS[7][2] ), .B(n3037), .S(n48), .Z(n1910) );
  MUX2_X1 U2311 ( .A(\REGISTERS[7][1] ), .B(n3038), .S(n48), .Z(n1909) );
  MUX2_X1 U2312 ( .A(\REGISTERS[7][0] ), .B(n3039), .S(n48), .Z(n1908) );
  OAI21_X1 U2313 ( .B1(n3040), .B2(n3056), .A(n3042), .ZN(n3055) );
  NAND3_X1 U2314 ( .A1(n3057), .A2(n3058), .A3(n3059), .ZN(n3040) );
  MUX2_X1 U2315 ( .A(\REGISTERS[8][31] ), .B(n3007), .S(n50), .Z(n1907) );
  MUX2_X1 U2316 ( .A(\REGISTERS[8][30] ), .B(n3009), .S(n50), .Z(n1906) );
  MUX2_X1 U2317 ( .A(\REGISTERS[8][29] ), .B(n3010), .S(n50), .Z(n1905) );
  MUX2_X1 U2318 ( .A(\REGISTERS[8][28] ), .B(n3011), .S(n50), .Z(n1904) );
  MUX2_X1 U2319 ( .A(\REGISTERS[8][27] ), .B(n3012), .S(n50), .Z(n1903) );
  MUX2_X1 U2320 ( .A(\REGISTERS[8][26] ), .B(n3013), .S(n50), .Z(n1902) );
  MUX2_X1 U2321 ( .A(\REGISTERS[8][25] ), .B(n3014), .S(n50), .Z(n1901) );
  MUX2_X1 U2322 ( .A(\REGISTERS[8][24] ), .B(n3015), .S(n50), .Z(n1900) );
  MUX2_X1 U2323 ( .A(\REGISTERS[8][23] ), .B(n3016), .S(n50), .Z(n1899) );
  MUX2_X1 U2324 ( .A(\REGISTERS[8][22] ), .B(n3017), .S(n50), .Z(n1898) );
  MUX2_X1 U2325 ( .A(\REGISTERS[8][21] ), .B(n3018), .S(n50), .Z(n1897) );
  MUX2_X1 U2326 ( .A(\REGISTERS[8][20] ), .B(n3019), .S(n50), .Z(n1896) );
  MUX2_X1 U2327 ( .A(\REGISTERS[8][19] ), .B(n3020), .S(n50), .Z(n1895) );
  MUX2_X1 U2328 ( .A(\REGISTERS[8][18] ), .B(n3021), .S(n50), .Z(n1894) );
  MUX2_X1 U2329 ( .A(\REGISTERS[8][17] ), .B(n3022), .S(n50), .Z(n1893) );
  MUX2_X1 U2330 ( .A(\REGISTERS[8][16] ), .B(n3023), .S(n50), .Z(n1892) );
  MUX2_X1 U2331 ( .A(\REGISTERS[8][15] ), .B(n3024), .S(n50), .Z(n1891) );
  MUX2_X1 U2332 ( .A(\REGISTERS[8][14] ), .B(n3025), .S(n50), .Z(n1890) );
  MUX2_X1 U2333 ( .A(\REGISTERS[8][13] ), .B(n3026), .S(n50), .Z(n1889) );
  MUX2_X1 U2334 ( .A(\REGISTERS[8][12] ), .B(n3027), .S(n50), .Z(n1888) );
  MUX2_X1 U2335 ( .A(\REGISTERS[8][11] ), .B(n3028), .S(n50), .Z(n1887) );
  MUX2_X1 U2336 ( .A(\REGISTERS[8][10] ), .B(n3029), .S(n50), .Z(n1886) );
  MUX2_X1 U2337 ( .A(\REGISTERS[8][9] ), .B(n3030), .S(n50), .Z(n1885) );
  MUX2_X1 U2338 ( .A(\REGISTERS[8][8] ), .B(n3031), .S(n50), .Z(n1884) );
  MUX2_X1 U2339 ( .A(\REGISTERS[8][7] ), .B(n3032), .S(n50), .Z(n1883) );
  MUX2_X1 U2340 ( .A(\REGISTERS[8][6] ), .B(n3033), .S(n50), .Z(n1882) );
  MUX2_X1 U2341 ( .A(\REGISTERS[8][5] ), .B(n3034), .S(n50), .Z(n1881) );
  MUX2_X1 U2342 ( .A(\REGISTERS[8][4] ), .B(n3035), .S(n50), .Z(n1880) );
  MUX2_X1 U2343 ( .A(\REGISTERS[8][3] ), .B(n3036), .S(n50), .Z(n1879) );
  MUX2_X1 U2344 ( .A(\REGISTERS[8][2] ), .B(n3037), .S(n50), .Z(n1878) );
  MUX2_X1 U2345 ( .A(\REGISTERS[8][1] ), .B(n3038), .S(n50), .Z(n1877) );
  MUX2_X1 U2346 ( .A(\REGISTERS[8][0] ), .B(n3039), .S(n50), .Z(n1876) );
  OAI21_X1 U2347 ( .B1(n3041), .B2(n3061), .A(n3042), .ZN(n3060) );
  MUX2_X1 U2348 ( .A(\REGISTERS[9][31] ), .B(n3007), .S(n44), .Z(n1875) );
  MUX2_X1 U2349 ( .A(\REGISTERS[9][30] ), .B(n3009), .S(n44), .Z(n1874) );
  MUX2_X1 U2350 ( .A(\REGISTERS[9][29] ), .B(n3010), .S(n44), .Z(n1873) );
  MUX2_X1 U2351 ( .A(\REGISTERS[9][28] ), .B(n3011), .S(n44), .Z(n1872) );
  MUX2_X1 U2352 ( .A(\REGISTERS[9][27] ), .B(n3012), .S(n44), .Z(n1871) );
  MUX2_X1 U2353 ( .A(\REGISTERS[9][26] ), .B(n3013), .S(n44), .Z(n1870) );
  MUX2_X1 U2354 ( .A(\REGISTERS[9][25] ), .B(n3014), .S(n44), .Z(n1869) );
  MUX2_X1 U2355 ( .A(\REGISTERS[9][24] ), .B(n3015), .S(n44), .Z(n1868) );
  MUX2_X1 U2356 ( .A(\REGISTERS[9][23] ), .B(n3016), .S(n44), .Z(n1867) );
  MUX2_X1 U2357 ( .A(\REGISTERS[9][22] ), .B(n3017), .S(n44), .Z(n1866) );
  MUX2_X1 U2358 ( .A(\REGISTERS[9][21] ), .B(n3018), .S(n44), .Z(n1865) );
  MUX2_X1 U2359 ( .A(\REGISTERS[9][20] ), .B(n3019), .S(n44), .Z(n1864) );
  MUX2_X1 U2360 ( .A(\REGISTERS[9][19] ), .B(n3020), .S(n44), .Z(n1863) );
  MUX2_X1 U2361 ( .A(\REGISTERS[9][18] ), .B(n3021), .S(n44), .Z(n1862) );
  MUX2_X1 U2362 ( .A(\REGISTERS[9][17] ), .B(n3022), .S(n44), .Z(n1861) );
  MUX2_X1 U2363 ( .A(\REGISTERS[9][16] ), .B(n3023), .S(n44), .Z(n1860) );
  MUX2_X1 U2364 ( .A(\REGISTERS[9][15] ), .B(n3024), .S(n44), .Z(n1859) );
  MUX2_X1 U2365 ( .A(\REGISTERS[9][14] ), .B(n3025), .S(n44), .Z(n1858) );
  MUX2_X1 U2366 ( .A(\REGISTERS[9][13] ), .B(n3026), .S(n44), .Z(n1857) );
  MUX2_X1 U2367 ( .A(\REGISTERS[9][12] ), .B(n3027), .S(n44), .Z(n1856) );
  MUX2_X1 U2368 ( .A(\REGISTERS[9][11] ), .B(n3028), .S(n44), .Z(n1855) );
  MUX2_X1 U2369 ( .A(\REGISTERS[9][10] ), .B(n3029), .S(n44), .Z(n1854) );
  MUX2_X1 U2370 ( .A(\REGISTERS[9][9] ), .B(n3030), .S(n44), .Z(n1853) );
  MUX2_X1 U2371 ( .A(\REGISTERS[9][8] ), .B(n3031), .S(n44), .Z(n1852) );
  MUX2_X1 U2372 ( .A(\REGISTERS[9][7] ), .B(n3032), .S(n44), .Z(n1851) );
  MUX2_X1 U2373 ( .A(\REGISTERS[9][6] ), .B(n3033), .S(n44), .Z(n1850) );
  MUX2_X1 U2374 ( .A(\REGISTERS[9][5] ), .B(n3034), .S(n44), .Z(n1849) );
  MUX2_X1 U2375 ( .A(\REGISTERS[9][4] ), .B(n3035), .S(n44), .Z(n1848) );
  MUX2_X1 U2376 ( .A(\REGISTERS[9][3] ), .B(n3036), .S(n44), .Z(n1847) );
  MUX2_X1 U2377 ( .A(\REGISTERS[9][2] ), .B(n3037), .S(n44), .Z(n1846) );
  MUX2_X1 U2378 ( .A(\REGISTERS[9][1] ), .B(n3038), .S(n44), .Z(n1845) );
  MUX2_X1 U2379 ( .A(\REGISTERS[9][0] ), .B(n3039), .S(n44), .Z(n1844) );
  OAI21_X1 U2380 ( .B1(n3044), .B2(n3061), .A(n3042), .ZN(n3062) );
  MUX2_X1 U2381 ( .A(\REGISTERS[10][31] ), .B(n3007), .S(n46), .Z(n1843) );
  MUX2_X1 U2382 ( .A(\REGISTERS[10][30] ), .B(n3009), .S(n46), .Z(n1842) );
  MUX2_X1 U2383 ( .A(\REGISTERS[10][29] ), .B(n3010), .S(n46), .Z(n1841) );
  MUX2_X1 U2384 ( .A(\REGISTERS[10][28] ), .B(n3011), .S(n46), .Z(n1840) );
  MUX2_X1 U2385 ( .A(\REGISTERS[10][27] ), .B(n3012), .S(n46), .Z(n1839) );
  MUX2_X1 U2386 ( .A(\REGISTERS[10][26] ), .B(n3013), .S(n46), .Z(n1838) );
  MUX2_X1 U2387 ( .A(\REGISTERS[10][25] ), .B(n3014), .S(n46), .Z(n1837) );
  MUX2_X1 U2388 ( .A(\REGISTERS[10][24] ), .B(n3015), .S(n46), .Z(n1836) );
  MUX2_X1 U2389 ( .A(\REGISTERS[10][23] ), .B(n3016), .S(n46), .Z(n1835) );
  MUX2_X1 U2390 ( .A(\REGISTERS[10][22] ), .B(n3017), .S(n46), .Z(n1834) );
  MUX2_X1 U2391 ( .A(\REGISTERS[10][21] ), .B(n3018), .S(n46), .Z(n1833) );
  MUX2_X1 U2392 ( .A(\REGISTERS[10][20] ), .B(n3019), .S(n46), .Z(n1832) );
  MUX2_X1 U2393 ( .A(\REGISTERS[10][19] ), .B(n3020), .S(n46), .Z(n1831) );
  MUX2_X1 U2394 ( .A(\REGISTERS[10][18] ), .B(n3021), .S(n46), .Z(n1830) );
  MUX2_X1 U2395 ( .A(\REGISTERS[10][17] ), .B(n3022), .S(n46), .Z(n1829) );
  MUX2_X1 U2396 ( .A(\REGISTERS[10][16] ), .B(n3023), .S(n46), .Z(n1828) );
  MUX2_X1 U2397 ( .A(\REGISTERS[10][15] ), .B(n3024), .S(n46), .Z(n1827) );
  MUX2_X1 U2398 ( .A(\REGISTERS[10][14] ), .B(n3025), .S(n46), .Z(n1826) );
  MUX2_X1 U2399 ( .A(\REGISTERS[10][13] ), .B(n3026), .S(n46), .Z(n1825) );
  MUX2_X1 U2400 ( .A(\REGISTERS[10][12] ), .B(n3027), .S(n46), .Z(n1824) );
  MUX2_X1 U2401 ( .A(\REGISTERS[10][11] ), .B(n3028), .S(n46), .Z(n1823) );
  MUX2_X1 U2402 ( .A(\REGISTERS[10][10] ), .B(n3029), .S(n46), .Z(n1822) );
  MUX2_X1 U2403 ( .A(\REGISTERS[10][9] ), .B(n3030), .S(n46), .Z(n1821) );
  MUX2_X1 U2404 ( .A(\REGISTERS[10][8] ), .B(n3031), .S(n46), .Z(n1820) );
  MUX2_X1 U2405 ( .A(\REGISTERS[10][7] ), .B(n3032), .S(n46), .Z(n1819) );
  MUX2_X1 U2406 ( .A(\REGISTERS[10][6] ), .B(n3033), .S(n46), .Z(n1818) );
  MUX2_X1 U2407 ( .A(\REGISTERS[10][5] ), .B(n3034), .S(n46), .Z(n1817) );
  MUX2_X1 U2408 ( .A(\REGISTERS[10][4] ), .B(n3035), .S(n46), .Z(n1816) );
  MUX2_X1 U2409 ( .A(\REGISTERS[10][3] ), .B(n3036), .S(n46), .Z(n1815) );
  MUX2_X1 U2410 ( .A(\REGISTERS[10][2] ), .B(n3037), .S(n46), .Z(n1814) );
  MUX2_X1 U2411 ( .A(\REGISTERS[10][1] ), .B(n3038), .S(n46), .Z(n1813) );
  MUX2_X1 U2412 ( .A(\REGISTERS[10][0] ), .B(n3039), .S(n46), .Z(n1812) );
  OAI21_X1 U2413 ( .B1(n3046), .B2(n3061), .A(n3042), .ZN(n3063) );
  MUX2_X1 U2414 ( .A(\REGISTERS[11][31] ), .B(n3007), .S(n40), .Z(n1811) );
  MUX2_X1 U2415 ( .A(\REGISTERS[11][30] ), .B(n3009), .S(n40), .Z(n1810) );
  MUX2_X1 U2416 ( .A(\REGISTERS[11][29] ), .B(n3010), .S(n40), .Z(n1809) );
  MUX2_X1 U2417 ( .A(\REGISTERS[11][28] ), .B(n3011), .S(n40), .Z(n1808) );
  MUX2_X1 U2418 ( .A(\REGISTERS[11][27] ), .B(n3012), .S(n40), .Z(n1807) );
  MUX2_X1 U2419 ( .A(\REGISTERS[11][26] ), .B(n3013), .S(n40), .Z(n1806) );
  MUX2_X1 U2420 ( .A(\REGISTERS[11][25] ), .B(n3014), .S(n40), .Z(n1805) );
  MUX2_X1 U2421 ( .A(\REGISTERS[11][24] ), .B(n3015), .S(n40), .Z(n1804) );
  MUX2_X1 U2422 ( .A(\REGISTERS[11][23] ), .B(n3016), .S(n40), .Z(n1803) );
  MUX2_X1 U2423 ( .A(\REGISTERS[11][22] ), .B(n3017), .S(n40), .Z(n1802) );
  MUX2_X1 U2424 ( .A(\REGISTERS[11][21] ), .B(n3018), .S(n40), .Z(n1801) );
  MUX2_X1 U2425 ( .A(\REGISTERS[11][20] ), .B(n3019), .S(n40), .Z(n1800) );
  MUX2_X1 U2426 ( .A(\REGISTERS[11][19] ), .B(n3020), .S(n40), .Z(n1799) );
  MUX2_X1 U2427 ( .A(\REGISTERS[11][18] ), .B(n3021), .S(n40), .Z(n1798) );
  MUX2_X1 U2428 ( .A(\REGISTERS[11][17] ), .B(n3022), .S(n40), .Z(n1797) );
  MUX2_X1 U2429 ( .A(\REGISTERS[11][16] ), .B(n3023), .S(n40), .Z(n1796) );
  MUX2_X1 U2430 ( .A(\REGISTERS[11][15] ), .B(n3024), .S(n40), .Z(n1795) );
  MUX2_X1 U2431 ( .A(\REGISTERS[11][14] ), .B(n3025), .S(n40), .Z(n1794) );
  MUX2_X1 U2432 ( .A(\REGISTERS[11][13] ), .B(n3026), .S(n40), .Z(n1793) );
  MUX2_X1 U2433 ( .A(\REGISTERS[11][12] ), .B(n3027), .S(n40), .Z(n1792) );
  MUX2_X1 U2434 ( .A(\REGISTERS[11][11] ), .B(n3028), .S(n40), .Z(n1791) );
  MUX2_X1 U2435 ( .A(\REGISTERS[11][10] ), .B(n3029), .S(n40), .Z(n1790) );
  MUX2_X1 U2436 ( .A(\REGISTERS[11][9] ), .B(n3030), .S(n40), .Z(n1789) );
  MUX2_X1 U2437 ( .A(\REGISTERS[11][8] ), .B(n3031), .S(n40), .Z(n1788) );
  MUX2_X1 U2438 ( .A(\REGISTERS[11][7] ), .B(n3032), .S(n40), .Z(n1787) );
  MUX2_X1 U2439 ( .A(\REGISTERS[11][6] ), .B(n3033), .S(n40), .Z(n1786) );
  MUX2_X1 U2440 ( .A(\REGISTERS[11][5] ), .B(n3034), .S(n40), .Z(n1785) );
  MUX2_X1 U2441 ( .A(\REGISTERS[11][4] ), .B(n3035), .S(n40), .Z(n1784) );
  MUX2_X1 U2442 ( .A(\REGISTERS[11][3] ), .B(n3036), .S(n40), .Z(n1783) );
  MUX2_X1 U2443 ( .A(\REGISTERS[11][2] ), .B(n3037), .S(n40), .Z(n1782) );
  MUX2_X1 U2444 ( .A(\REGISTERS[11][1] ), .B(n3038), .S(n40), .Z(n1781) );
  MUX2_X1 U2445 ( .A(\REGISTERS[11][0] ), .B(n3039), .S(n40), .Z(n1780) );
  OAI21_X1 U2446 ( .B1(n3048), .B2(n3061), .A(n3042), .ZN(n3064) );
  MUX2_X1 U2447 ( .A(\REGISTERS[12][31] ), .B(n3007), .S(n42), .Z(n1779) );
  MUX2_X1 U2448 ( .A(\REGISTERS[12][30] ), .B(n3009), .S(n42), .Z(n1778) );
  MUX2_X1 U2449 ( .A(\REGISTERS[12][29] ), .B(n3010), .S(n42), .Z(n1777) );
  MUX2_X1 U2450 ( .A(\REGISTERS[12][28] ), .B(n3011), .S(n42), .Z(n1776) );
  MUX2_X1 U2451 ( .A(\REGISTERS[12][27] ), .B(n3012), .S(n42), .Z(n1775) );
  MUX2_X1 U2452 ( .A(\REGISTERS[12][26] ), .B(n3013), .S(n42), .Z(n1774) );
  MUX2_X1 U2453 ( .A(\REGISTERS[12][25] ), .B(n3014), .S(n42), .Z(n1773) );
  MUX2_X1 U2454 ( .A(\REGISTERS[12][24] ), .B(n3015), .S(n42), .Z(n1772) );
  MUX2_X1 U2455 ( .A(\REGISTERS[12][23] ), .B(n3016), .S(n42), .Z(n1771) );
  MUX2_X1 U2456 ( .A(\REGISTERS[12][22] ), .B(n3017), .S(n42), .Z(n1770) );
  MUX2_X1 U2457 ( .A(\REGISTERS[12][21] ), .B(n3018), .S(n42), .Z(n1769) );
  MUX2_X1 U2458 ( .A(\REGISTERS[12][20] ), .B(n3019), .S(n42), .Z(n1768) );
  MUX2_X1 U2459 ( .A(\REGISTERS[12][19] ), .B(n3020), .S(n42), .Z(n1767) );
  MUX2_X1 U2460 ( .A(\REGISTERS[12][18] ), .B(n3021), .S(n42), .Z(n1766) );
  MUX2_X1 U2461 ( .A(\REGISTERS[12][17] ), .B(n3022), .S(n42), .Z(n1765) );
  MUX2_X1 U2462 ( .A(\REGISTERS[12][16] ), .B(n3023), .S(n42), .Z(n1764) );
  MUX2_X1 U2463 ( .A(\REGISTERS[12][15] ), .B(n3024), .S(n42), .Z(n1763) );
  MUX2_X1 U2464 ( .A(\REGISTERS[12][14] ), .B(n3025), .S(n42), .Z(n1762) );
  MUX2_X1 U2465 ( .A(\REGISTERS[12][13] ), .B(n3026), .S(n42), .Z(n1761) );
  MUX2_X1 U2466 ( .A(\REGISTERS[12][12] ), .B(n3027), .S(n42), .Z(n1760) );
  MUX2_X1 U2467 ( .A(\REGISTERS[12][11] ), .B(n3028), .S(n42), .Z(n1759) );
  MUX2_X1 U2468 ( .A(\REGISTERS[12][10] ), .B(n3029), .S(n42), .Z(n1758) );
  MUX2_X1 U2469 ( .A(\REGISTERS[12][9] ), .B(n3030), .S(n42), .Z(n1757) );
  MUX2_X1 U2470 ( .A(\REGISTERS[12][8] ), .B(n3031), .S(n42), .Z(n1756) );
  MUX2_X1 U2471 ( .A(\REGISTERS[12][7] ), .B(n3032), .S(n42), .Z(n1755) );
  MUX2_X1 U2472 ( .A(\REGISTERS[12][6] ), .B(n3033), .S(n42), .Z(n1754) );
  MUX2_X1 U2473 ( .A(\REGISTERS[12][5] ), .B(n3034), .S(n42), .Z(n1753) );
  MUX2_X1 U2474 ( .A(\REGISTERS[12][4] ), .B(n3035), .S(n42), .Z(n1752) );
  MUX2_X1 U2475 ( .A(\REGISTERS[12][3] ), .B(n3036), .S(n42), .Z(n1751) );
  MUX2_X1 U2476 ( .A(\REGISTERS[12][2] ), .B(n3037), .S(n42), .Z(n1750) );
  MUX2_X1 U2477 ( .A(\REGISTERS[12][1] ), .B(n3038), .S(n42), .Z(n1749) );
  MUX2_X1 U2478 ( .A(\REGISTERS[12][0] ), .B(n3039), .S(n42), .Z(n1748) );
  OAI21_X1 U2479 ( .B1(n3050), .B2(n3061), .A(n3042), .ZN(n3065) );
  MUX2_X1 U2480 ( .A(\REGISTERS[13][31] ), .B(n3007), .S(n36), .Z(n1747) );
  MUX2_X1 U2481 ( .A(\REGISTERS[13][30] ), .B(n3009), .S(n36), .Z(n1746) );
  MUX2_X1 U2482 ( .A(\REGISTERS[13][29] ), .B(n3010), .S(n36), .Z(n1745) );
  MUX2_X1 U2483 ( .A(\REGISTERS[13][28] ), .B(n3011), .S(n36), .Z(n1744) );
  MUX2_X1 U2484 ( .A(\REGISTERS[13][27] ), .B(n3012), .S(n36), .Z(n1743) );
  MUX2_X1 U2485 ( .A(\REGISTERS[13][26] ), .B(n3013), .S(n36), .Z(n1742) );
  MUX2_X1 U2486 ( .A(\REGISTERS[13][25] ), .B(n3014), .S(n36), .Z(n1741) );
  MUX2_X1 U2487 ( .A(\REGISTERS[13][24] ), .B(n3015), .S(n36), .Z(n1740) );
  MUX2_X1 U2488 ( .A(\REGISTERS[13][23] ), .B(n3016), .S(n36), .Z(n1739) );
  MUX2_X1 U2489 ( .A(\REGISTERS[13][22] ), .B(n3017), .S(n36), .Z(n1738) );
  MUX2_X1 U2490 ( .A(\REGISTERS[13][21] ), .B(n3018), .S(n36), .Z(n1737) );
  MUX2_X1 U2491 ( .A(\REGISTERS[13][20] ), .B(n3019), .S(n36), .Z(n1736) );
  MUX2_X1 U2492 ( .A(\REGISTERS[13][19] ), .B(n3020), .S(n36), .Z(n1735) );
  MUX2_X1 U2493 ( .A(\REGISTERS[13][18] ), .B(n3021), .S(n36), .Z(n1734) );
  MUX2_X1 U2494 ( .A(\REGISTERS[13][17] ), .B(n3022), .S(n36), .Z(n1733) );
  MUX2_X1 U2495 ( .A(\REGISTERS[13][16] ), .B(n3023), .S(n36), .Z(n1732) );
  MUX2_X1 U2496 ( .A(\REGISTERS[13][15] ), .B(n3024), .S(n36), .Z(n1731) );
  MUX2_X1 U2497 ( .A(\REGISTERS[13][14] ), .B(n3025), .S(n36), .Z(n1730) );
  MUX2_X1 U2498 ( .A(\REGISTERS[13][13] ), .B(n3026), .S(n36), .Z(n1729) );
  MUX2_X1 U2499 ( .A(\REGISTERS[13][12] ), .B(n3027), .S(n36), .Z(n1728) );
  MUX2_X1 U2500 ( .A(\REGISTERS[13][11] ), .B(n3028), .S(n36), .Z(n1727) );
  MUX2_X1 U2501 ( .A(\REGISTERS[13][10] ), .B(n3029), .S(n36), .Z(n1726) );
  MUX2_X1 U2502 ( .A(\REGISTERS[13][9] ), .B(n3030), .S(n36), .Z(n1725) );
  MUX2_X1 U2503 ( .A(\REGISTERS[13][8] ), .B(n3031), .S(n36), .Z(n1724) );
  MUX2_X1 U2504 ( .A(\REGISTERS[13][7] ), .B(n3032), .S(n36), .Z(n1723) );
  MUX2_X1 U2505 ( .A(\REGISTERS[13][6] ), .B(n3033), .S(n36), .Z(n1722) );
  MUX2_X1 U2506 ( .A(\REGISTERS[13][5] ), .B(n3034), .S(n36), .Z(n1721) );
  MUX2_X1 U2507 ( .A(\REGISTERS[13][4] ), .B(n3035), .S(n36), .Z(n1720) );
  MUX2_X1 U2508 ( .A(\REGISTERS[13][3] ), .B(n3036), .S(n36), .Z(n1719) );
  MUX2_X1 U2509 ( .A(\REGISTERS[13][2] ), .B(n3037), .S(n36), .Z(n1718) );
  MUX2_X1 U2510 ( .A(\REGISTERS[13][1] ), .B(n3038), .S(n36), .Z(n1717) );
  MUX2_X1 U2511 ( .A(\REGISTERS[13][0] ), .B(n3039), .S(n36), .Z(n1716) );
  OAI21_X1 U2512 ( .B1(n3052), .B2(n3061), .A(n3042), .ZN(n3066) );
  MUX2_X1 U2513 ( .A(\REGISTERS[14][31] ), .B(n3007), .S(n38), .Z(n1715) );
  MUX2_X1 U2514 ( .A(\REGISTERS[14][30] ), .B(n3009), .S(n38), .Z(n1714) );
  MUX2_X1 U2515 ( .A(\REGISTERS[14][29] ), .B(n3010), .S(n38), .Z(n1713) );
  MUX2_X1 U2516 ( .A(\REGISTERS[14][28] ), .B(n3011), .S(n38), .Z(n1712) );
  MUX2_X1 U2517 ( .A(\REGISTERS[14][27] ), .B(n3012), .S(n38), .Z(n1711) );
  MUX2_X1 U2518 ( .A(\REGISTERS[14][26] ), .B(n3013), .S(n38), .Z(n1710) );
  MUX2_X1 U2519 ( .A(\REGISTERS[14][25] ), .B(n3014), .S(n38), .Z(n1709) );
  MUX2_X1 U2520 ( .A(\REGISTERS[14][24] ), .B(n3015), .S(n38), .Z(n1708) );
  MUX2_X1 U2521 ( .A(\REGISTERS[14][23] ), .B(n3016), .S(n38), .Z(n1707) );
  MUX2_X1 U2522 ( .A(\REGISTERS[14][22] ), .B(n3017), .S(n38), .Z(n1706) );
  MUX2_X1 U2523 ( .A(\REGISTERS[14][21] ), .B(n3018), .S(n38), .Z(n1705) );
  MUX2_X1 U2524 ( .A(\REGISTERS[14][20] ), .B(n3019), .S(n38), .Z(n1704) );
  MUX2_X1 U2525 ( .A(\REGISTERS[14][19] ), .B(n3020), .S(n38), .Z(n1703) );
  MUX2_X1 U2526 ( .A(\REGISTERS[14][18] ), .B(n3021), .S(n38), .Z(n1702) );
  MUX2_X1 U2527 ( .A(\REGISTERS[14][17] ), .B(n3022), .S(n38), .Z(n1701) );
  MUX2_X1 U2528 ( .A(\REGISTERS[14][16] ), .B(n3023), .S(n38), .Z(n1700) );
  MUX2_X1 U2529 ( .A(\REGISTERS[14][15] ), .B(n3024), .S(n38), .Z(n1699) );
  MUX2_X1 U2530 ( .A(\REGISTERS[14][14] ), .B(n3025), .S(n38), .Z(n1698) );
  MUX2_X1 U2531 ( .A(\REGISTERS[14][13] ), .B(n3026), .S(n38), .Z(n1697) );
  MUX2_X1 U2532 ( .A(\REGISTERS[14][12] ), .B(n3027), .S(n38), .Z(n1696) );
  MUX2_X1 U2533 ( .A(\REGISTERS[14][11] ), .B(n3028), .S(n38), .Z(n1695) );
  MUX2_X1 U2534 ( .A(\REGISTERS[14][10] ), .B(n3029), .S(n38), .Z(n1694) );
  MUX2_X1 U2535 ( .A(\REGISTERS[14][9] ), .B(n3030), .S(n38), .Z(n1693) );
  MUX2_X1 U2536 ( .A(\REGISTERS[14][8] ), .B(n3031), .S(n38), .Z(n1692) );
  MUX2_X1 U2537 ( .A(\REGISTERS[14][7] ), .B(n3032), .S(n38), .Z(n1691) );
  MUX2_X1 U2538 ( .A(\REGISTERS[14][6] ), .B(n3033), .S(n38), .Z(n1690) );
  MUX2_X1 U2539 ( .A(\REGISTERS[14][5] ), .B(n3034), .S(n38), .Z(n1689) );
  MUX2_X1 U2540 ( .A(\REGISTERS[14][4] ), .B(n3035), .S(n38), .Z(n1688) );
  MUX2_X1 U2541 ( .A(\REGISTERS[14][3] ), .B(n3036), .S(n38), .Z(n1687) );
  MUX2_X1 U2542 ( .A(\REGISTERS[14][2] ), .B(n3037), .S(n38), .Z(n1686) );
  MUX2_X1 U2543 ( .A(\REGISTERS[14][1] ), .B(n3038), .S(n38), .Z(n1685) );
  MUX2_X1 U2544 ( .A(\REGISTERS[14][0] ), .B(n3039), .S(n38), .Z(n1684) );
  OAI21_X1 U2545 ( .B1(n3054), .B2(n3061), .A(n3042), .ZN(n3067) );
  MUX2_X1 U2546 ( .A(\REGISTERS[15][31] ), .B(n3007), .S(n32), .Z(n1683) );
  MUX2_X1 U2547 ( .A(\REGISTERS[15][30] ), .B(n3009), .S(n32), .Z(n1682) );
  MUX2_X1 U2548 ( .A(\REGISTERS[15][29] ), .B(n3010), .S(n32), .Z(n1681) );
  MUX2_X1 U2549 ( .A(\REGISTERS[15][28] ), .B(n3011), .S(n32), .Z(n1680) );
  MUX2_X1 U2550 ( .A(\REGISTERS[15][27] ), .B(n3012), .S(n32), .Z(n1679) );
  MUX2_X1 U2551 ( .A(\REGISTERS[15][26] ), .B(n3013), .S(n32), .Z(n1678) );
  MUX2_X1 U2552 ( .A(\REGISTERS[15][25] ), .B(n3014), .S(n32), .Z(n1677) );
  MUX2_X1 U2553 ( .A(\REGISTERS[15][24] ), .B(n3015), .S(n32), .Z(n1676) );
  MUX2_X1 U2554 ( .A(\REGISTERS[15][23] ), .B(n3016), .S(n32), .Z(n1675) );
  MUX2_X1 U2555 ( .A(\REGISTERS[15][22] ), .B(n3017), .S(n32), .Z(n1674) );
  MUX2_X1 U2556 ( .A(\REGISTERS[15][21] ), .B(n3018), .S(n32), .Z(n1673) );
  MUX2_X1 U2557 ( .A(\REGISTERS[15][20] ), .B(n3019), .S(n32), .Z(n1672) );
  MUX2_X1 U2558 ( .A(\REGISTERS[15][19] ), .B(n3020), .S(n32), .Z(n1671) );
  MUX2_X1 U2559 ( .A(\REGISTERS[15][18] ), .B(n3021), .S(n32), .Z(n1670) );
  MUX2_X1 U2560 ( .A(\REGISTERS[15][17] ), .B(n3022), .S(n32), .Z(n1669) );
  MUX2_X1 U2561 ( .A(\REGISTERS[15][16] ), .B(n3023), .S(n32), .Z(n1668) );
  MUX2_X1 U2562 ( .A(\REGISTERS[15][15] ), .B(n3024), .S(n32), .Z(n1667) );
  MUX2_X1 U2563 ( .A(\REGISTERS[15][14] ), .B(n3025), .S(n32), .Z(n1666) );
  MUX2_X1 U2564 ( .A(\REGISTERS[15][13] ), .B(n3026), .S(n32), .Z(n1665) );
  MUX2_X1 U2565 ( .A(\REGISTERS[15][12] ), .B(n3027), .S(n32), .Z(n1664) );
  MUX2_X1 U2566 ( .A(\REGISTERS[15][11] ), .B(n3028), .S(n32), .Z(n1663) );
  MUX2_X1 U2567 ( .A(\REGISTERS[15][10] ), .B(n3029), .S(n32), .Z(n1662) );
  MUX2_X1 U2568 ( .A(\REGISTERS[15][9] ), .B(n3030), .S(n32), .Z(n1661) );
  MUX2_X1 U2569 ( .A(\REGISTERS[15][8] ), .B(n3031), .S(n32), .Z(n1660) );
  MUX2_X1 U2570 ( .A(\REGISTERS[15][7] ), .B(n3032), .S(n32), .Z(n1659) );
  MUX2_X1 U2571 ( .A(\REGISTERS[15][6] ), .B(n3033), .S(n32), .Z(n1658) );
  MUX2_X1 U2572 ( .A(\REGISTERS[15][5] ), .B(n3034), .S(n32), .Z(n1657) );
  MUX2_X1 U2573 ( .A(\REGISTERS[15][4] ), .B(n3035), .S(n32), .Z(n1656) );
  MUX2_X1 U2574 ( .A(\REGISTERS[15][3] ), .B(n3036), .S(n32), .Z(n1655) );
  MUX2_X1 U2575 ( .A(\REGISTERS[15][2] ), .B(n3037), .S(n32), .Z(n1654) );
  MUX2_X1 U2576 ( .A(\REGISTERS[15][1] ), .B(n3038), .S(n32), .Z(n1653) );
  MUX2_X1 U2577 ( .A(\REGISTERS[15][0] ), .B(n3039), .S(n32), .Z(n1652) );
  OAI21_X1 U2578 ( .B1(n3056), .B2(n3061), .A(n3042), .ZN(n3068) );
  NAND3_X1 U2579 ( .A1(n3059), .A2(n3058), .A3(ADD_WR[3]), .ZN(n3061) );
  INV_X1 U2580 ( .A(ADD_WR[4]), .ZN(n3058) );
  MUX2_X1 U2581 ( .A(\REGISTERS[16][31] ), .B(n3007), .S(n34), .Z(n1651) );
  MUX2_X1 U2582 ( .A(\REGISTERS[16][30] ), .B(n3009), .S(n34), .Z(n1650) );
  MUX2_X1 U2583 ( .A(\REGISTERS[16][29] ), .B(n3010), .S(n34), .Z(n1649) );
  MUX2_X1 U2584 ( .A(\REGISTERS[16][28] ), .B(n3011), .S(n34), .Z(n1648) );
  MUX2_X1 U2585 ( .A(\REGISTERS[16][27] ), .B(n3012), .S(n34), .Z(n1647) );
  MUX2_X1 U2586 ( .A(\REGISTERS[16][26] ), .B(n3013), .S(n34), .Z(n1646) );
  MUX2_X1 U2587 ( .A(\REGISTERS[16][25] ), .B(n3014), .S(n34), .Z(n1645) );
  MUX2_X1 U2588 ( .A(\REGISTERS[16][24] ), .B(n3015), .S(n34), .Z(n1644) );
  MUX2_X1 U2589 ( .A(\REGISTERS[16][23] ), .B(n3016), .S(n34), .Z(n1643) );
  MUX2_X1 U2590 ( .A(\REGISTERS[16][22] ), .B(n3017), .S(n34), .Z(n1642) );
  MUX2_X1 U2591 ( .A(\REGISTERS[16][21] ), .B(n3018), .S(n34), .Z(n1641) );
  MUX2_X1 U2592 ( .A(\REGISTERS[16][20] ), .B(n3019), .S(n34), .Z(n1640) );
  MUX2_X1 U2593 ( .A(\REGISTERS[16][19] ), .B(n3020), .S(n34), .Z(n1639) );
  MUX2_X1 U2594 ( .A(\REGISTERS[16][18] ), .B(n3021), .S(n34), .Z(n1638) );
  MUX2_X1 U2595 ( .A(\REGISTERS[16][17] ), .B(n3022), .S(n34), .Z(n1637) );
  MUX2_X1 U2596 ( .A(\REGISTERS[16][16] ), .B(n3023), .S(n34), .Z(n1636) );
  MUX2_X1 U2597 ( .A(\REGISTERS[16][15] ), .B(n3024), .S(n34), .Z(n1635) );
  MUX2_X1 U2598 ( .A(\REGISTERS[16][14] ), .B(n3025), .S(n34), .Z(n1634) );
  MUX2_X1 U2599 ( .A(\REGISTERS[16][13] ), .B(n3026), .S(n34), .Z(n1633) );
  MUX2_X1 U2600 ( .A(\REGISTERS[16][12] ), .B(n3027), .S(n34), .Z(n1632) );
  MUX2_X1 U2601 ( .A(\REGISTERS[16][11] ), .B(n3028), .S(n34), .Z(n1631) );
  MUX2_X1 U2602 ( .A(\REGISTERS[16][10] ), .B(n3029), .S(n34), .Z(n1630) );
  MUX2_X1 U2603 ( .A(\REGISTERS[16][9] ), .B(n3030), .S(n34), .Z(n1629) );
  MUX2_X1 U2604 ( .A(\REGISTERS[16][8] ), .B(n3031), .S(n34), .Z(n1628) );
  MUX2_X1 U2605 ( .A(\REGISTERS[16][7] ), .B(n3032), .S(n34), .Z(n1627) );
  MUX2_X1 U2606 ( .A(\REGISTERS[16][6] ), .B(n3033), .S(n34), .Z(n1626) );
  MUX2_X1 U2607 ( .A(\REGISTERS[16][5] ), .B(n3034), .S(n34), .Z(n1625) );
  MUX2_X1 U2608 ( .A(\REGISTERS[16][4] ), .B(n3035), .S(n34), .Z(n1624) );
  MUX2_X1 U2609 ( .A(\REGISTERS[16][3] ), .B(n3036), .S(n34), .Z(n1623) );
  MUX2_X1 U2610 ( .A(\REGISTERS[16][2] ), .B(n3037), .S(n34), .Z(n1622) );
  MUX2_X1 U2611 ( .A(\REGISTERS[16][1] ), .B(n3038), .S(n34), .Z(n1621) );
  MUX2_X1 U2612 ( .A(\REGISTERS[16][0] ), .B(n3039), .S(n34), .Z(n1620) );
  OAI21_X1 U2613 ( .B1(n3041), .B2(n3070), .A(n3042), .ZN(n3069) );
  MUX2_X1 U2614 ( .A(\REGISTERS[17][31] ), .B(n3007), .S(n28), .Z(n1619) );
  MUX2_X1 U2615 ( .A(\REGISTERS[17][30] ), .B(n3009), .S(n28), .Z(n1618) );
  MUX2_X1 U2616 ( .A(\REGISTERS[17][29] ), .B(n3010), .S(n28), .Z(n1617) );
  MUX2_X1 U2617 ( .A(\REGISTERS[17][28] ), .B(n3011), .S(n28), .Z(n1616) );
  MUX2_X1 U2618 ( .A(\REGISTERS[17][27] ), .B(n3012), .S(n28), .Z(n1615) );
  MUX2_X1 U2619 ( .A(\REGISTERS[17][26] ), .B(n3013), .S(n28), .Z(n1614) );
  MUX2_X1 U2620 ( .A(\REGISTERS[17][25] ), .B(n3014), .S(n28), .Z(n1613) );
  MUX2_X1 U2621 ( .A(\REGISTERS[17][24] ), .B(n3015), .S(n28), .Z(n1612) );
  MUX2_X1 U2622 ( .A(\REGISTERS[17][23] ), .B(n3016), .S(n28), .Z(n1611) );
  MUX2_X1 U2623 ( .A(\REGISTERS[17][22] ), .B(n3017), .S(n28), .Z(n1610) );
  MUX2_X1 U2624 ( .A(\REGISTERS[17][21] ), .B(n3018), .S(n28), .Z(n1609) );
  MUX2_X1 U2625 ( .A(\REGISTERS[17][20] ), .B(n3019), .S(n28), .Z(n1608) );
  MUX2_X1 U2626 ( .A(\REGISTERS[17][19] ), .B(n3020), .S(n28), .Z(n1607) );
  MUX2_X1 U2627 ( .A(\REGISTERS[17][18] ), .B(n3021), .S(n28), .Z(n1606) );
  MUX2_X1 U2628 ( .A(\REGISTERS[17][17] ), .B(n3022), .S(n28), .Z(n1605) );
  MUX2_X1 U2629 ( .A(\REGISTERS[17][16] ), .B(n3023), .S(n28), .Z(n1604) );
  MUX2_X1 U2630 ( .A(\REGISTERS[17][15] ), .B(n3024), .S(n28), .Z(n1603) );
  MUX2_X1 U2631 ( .A(\REGISTERS[17][14] ), .B(n3025), .S(n28), .Z(n1602) );
  MUX2_X1 U2632 ( .A(\REGISTERS[17][13] ), .B(n3026), .S(n28), .Z(n1601) );
  MUX2_X1 U2633 ( .A(\REGISTERS[17][12] ), .B(n3027), .S(n28), .Z(n1600) );
  MUX2_X1 U2634 ( .A(\REGISTERS[17][11] ), .B(n3028), .S(n28), .Z(n1599) );
  MUX2_X1 U2635 ( .A(\REGISTERS[17][10] ), .B(n3029), .S(n28), .Z(n1598) );
  MUX2_X1 U2636 ( .A(\REGISTERS[17][9] ), .B(n3030), .S(n28), .Z(n1597) );
  MUX2_X1 U2637 ( .A(\REGISTERS[17][8] ), .B(n3031), .S(n28), .Z(n1596) );
  MUX2_X1 U2638 ( .A(\REGISTERS[17][7] ), .B(n3032), .S(n28), .Z(n1595) );
  MUX2_X1 U2639 ( .A(\REGISTERS[17][6] ), .B(n3033), .S(n28), .Z(n1594) );
  MUX2_X1 U2640 ( .A(\REGISTERS[17][5] ), .B(n3034), .S(n28), .Z(n1593) );
  MUX2_X1 U2641 ( .A(\REGISTERS[17][4] ), .B(n3035), .S(n28), .Z(n1592) );
  MUX2_X1 U2642 ( .A(\REGISTERS[17][3] ), .B(n3036), .S(n28), .Z(n1591) );
  MUX2_X1 U2643 ( .A(\REGISTERS[17][2] ), .B(n3037), .S(n28), .Z(n1590) );
  MUX2_X1 U2644 ( .A(\REGISTERS[17][1] ), .B(n3038), .S(n28), .Z(n1589) );
  MUX2_X1 U2645 ( .A(\REGISTERS[17][0] ), .B(n3039), .S(n28), .Z(n1588) );
  OAI21_X1 U2646 ( .B1(n3044), .B2(n3070), .A(n3042), .ZN(n3071) );
  MUX2_X1 U2647 ( .A(\REGISTERS[18][31] ), .B(n3007), .S(n30), .Z(n1587) );
  MUX2_X1 U2648 ( .A(\REGISTERS[18][30] ), .B(n3009), .S(n30), .Z(n1586) );
  MUX2_X1 U2649 ( .A(\REGISTERS[18][29] ), .B(n3010), .S(n30), .Z(n1585) );
  MUX2_X1 U2650 ( .A(\REGISTERS[18][28] ), .B(n3011), .S(n30), .Z(n1584) );
  MUX2_X1 U2651 ( .A(\REGISTERS[18][27] ), .B(n3012), .S(n30), .Z(n1583) );
  MUX2_X1 U2652 ( .A(\REGISTERS[18][26] ), .B(n3013), .S(n30), .Z(n1582) );
  MUX2_X1 U2653 ( .A(\REGISTERS[18][25] ), .B(n3014), .S(n30), .Z(n1581) );
  MUX2_X1 U2654 ( .A(\REGISTERS[18][24] ), .B(n3015), .S(n30), .Z(n1580) );
  MUX2_X1 U2655 ( .A(\REGISTERS[18][23] ), .B(n3016), .S(n30), .Z(n1579) );
  MUX2_X1 U2656 ( .A(\REGISTERS[18][22] ), .B(n3017), .S(n30), .Z(n1578) );
  MUX2_X1 U2657 ( .A(\REGISTERS[18][21] ), .B(n3018), .S(n30), .Z(n1577) );
  MUX2_X1 U2658 ( .A(\REGISTERS[18][20] ), .B(n3019), .S(n30), .Z(n1576) );
  MUX2_X1 U2659 ( .A(\REGISTERS[18][19] ), .B(n3020), .S(n30), .Z(n1575) );
  MUX2_X1 U2660 ( .A(\REGISTERS[18][18] ), .B(n3021), .S(n30), .Z(n1574) );
  MUX2_X1 U2661 ( .A(\REGISTERS[18][17] ), .B(n3022), .S(n30), .Z(n1573) );
  MUX2_X1 U2662 ( .A(\REGISTERS[18][16] ), .B(n3023), .S(n30), .Z(n1572) );
  MUX2_X1 U2663 ( .A(\REGISTERS[18][15] ), .B(n3024), .S(n30), .Z(n1571) );
  MUX2_X1 U2664 ( .A(\REGISTERS[18][14] ), .B(n3025), .S(n30), .Z(n1570) );
  MUX2_X1 U2665 ( .A(\REGISTERS[18][13] ), .B(n3026), .S(n30), .Z(n1569) );
  MUX2_X1 U2666 ( .A(\REGISTERS[18][12] ), .B(n3027), .S(n30), .Z(n1568) );
  MUX2_X1 U2667 ( .A(\REGISTERS[18][11] ), .B(n3028), .S(n30), .Z(n1567) );
  MUX2_X1 U2668 ( .A(\REGISTERS[18][10] ), .B(n3029), .S(n30), .Z(n1566) );
  MUX2_X1 U2669 ( .A(\REGISTERS[18][9] ), .B(n3030), .S(n30), .Z(n1565) );
  MUX2_X1 U2670 ( .A(\REGISTERS[18][8] ), .B(n3031), .S(n30), .Z(n1564) );
  MUX2_X1 U2671 ( .A(\REGISTERS[18][7] ), .B(n3032), .S(n30), .Z(n1563) );
  MUX2_X1 U2672 ( .A(\REGISTERS[18][6] ), .B(n3033), .S(n30), .Z(n1562) );
  MUX2_X1 U2673 ( .A(\REGISTERS[18][5] ), .B(n3034), .S(n30), .Z(n1561) );
  MUX2_X1 U2674 ( .A(\REGISTERS[18][4] ), .B(n3035), .S(n30), .Z(n1560) );
  MUX2_X1 U2675 ( .A(\REGISTERS[18][3] ), .B(n3036), .S(n30), .Z(n1559) );
  MUX2_X1 U2676 ( .A(\REGISTERS[18][2] ), .B(n3037), .S(n30), .Z(n1558) );
  MUX2_X1 U2677 ( .A(\REGISTERS[18][1] ), .B(n3038), .S(n30), .Z(n1557) );
  MUX2_X1 U2678 ( .A(\REGISTERS[18][0] ), .B(n3039), .S(n30), .Z(n1556) );
  OAI21_X1 U2679 ( .B1(n3046), .B2(n3070), .A(n3042), .ZN(n3072) );
  MUX2_X1 U2680 ( .A(\REGISTERS[19][31] ), .B(n3007), .S(n24), .Z(n1555) );
  MUX2_X1 U2681 ( .A(\REGISTERS[19][30] ), .B(n3009), .S(n24), .Z(n1554) );
  MUX2_X1 U2682 ( .A(\REGISTERS[19][29] ), .B(n3010), .S(n24), .Z(n1553) );
  MUX2_X1 U2683 ( .A(\REGISTERS[19][28] ), .B(n3011), .S(n24), .Z(n1552) );
  MUX2_X1 U2684 ( .A(\REGISTERS[19][27] ), .B(n3012), .S(n24), .Z(n1551) );
  MUX2_X1 U2685 ( .A(\REGISTERS[19][26] ), .B(n3013), .S(n24), .Z(n1550) );
  MUX2_X1 U2686 ( .A(\REGISTERS[19][25] ), .B(n3014), .S(n24), .Z(n1549) );
  MUX2_X1 U2687 ( .A(\REGISTERS[19][24] ), .B(n3015), .S(n24), .Z(n1548) );
  MUX2_X1 U2688 ( .A(\REGISTERS[19][23] ), .B(n3016), .S(n24), .Z(n1547) );
  MUX2_X1 U2689 ( .A(\REGISTERS[19][22] ), .B(n3017), .S(n24), .Z(n1546) );
  MUX2_X1 U2690 ( .A(\REGISTERS[19][21] ), .B(n3018), .S(n24), .Z(n1545) );
  MUX2_X1 U2691 ( .A(\REGISTERS[19][20] ), .B(n3019), .S(n24), .Z(n1544) );
  MUX2_X1 U2692 ( .A(\REGISTERS[19][19] ), .B(n3020), .S(n24), .Z(n1543) );
  MUX2_X1 U2693 ( .A(\REGISTERS[19][18] ), .B(n3021), .S(n24), .Z(n1542) );
  MUX2_X1 U2694 ( .A(\REGISTERS[19][17] ), .B(n3022), .S(n24), .Z(n1541) );
  MUX2_X1 U2695 ( .A(\REGISTERS[19][16] ), .B(n3023), .S(n24), .Z(n1540) );
  MUX2_X1 U2696 ( .A(\REGISTERS[19][15] ), .B(n3024), .S(n24), .Z(n1539) );
  MUX2_X1 U2697 ( .A(\REGISTERS[19][14] ), .B(n3025), .S(n24), .Z(n1538) );
  MUX2_X1 U2698 ( .A(\REGISTERS[19][13] ), .B(n3026), .S(n24), .Z(n1537) );
  MUX2_X1 U2699 ( .A(\REGISTERS[19][12] ), .B(n3027), .S(n24), .Z(n1536) );
  MUX2_X1 U2700 ( .A(\REGISTERS[19][11] ), .B(n3028), .S(n24), .Z(n1535) );
  MUX2_X1 U2701 ( .A(\REGISTERS[19][10] ), .B(n3029), .S(n24), .Z(n1534) );
  MUX2_X1 U2702 ( .A(\REGISTERS[19][9] ), .B(n3030), .S(n24), .Z(n1533) );
  MUX2_X1 U2703 ( .A(\REGISTERS[19][8] ), .B(n3031), .S(n24), .Z(n1532) );
  MUX2_X1 U2704 ( .A(\REGISTERS[19][7] ), .B(n3032), .S(n24), .Z(n1531) );
  MUX2_X1 U2705 ( .A(\REGISTERS[19][6] ), .B(n3033), .S(n24), .Z(n1530) );
  MUX2_X1 U2706 ( .A(\REGISTERS[19][5] ), .B(n3034), .S(n24), .Z(n1529) );
  MUX2_X1 U2707 ( .A(\REGISTERS[19][4] ), .B(n3035), .S(n24), .Z(n1528) );
  MUX2_X1 U2708 ( .A(\REGISTERS[19][3] ), .B(n3036), .S(n24), .Z(n1527) );
  MUX2_X1 U2709 ( .A(\REGISTERS[19][2] ), .B(n3037), .S(n24), .Z(n1526) );
  MUX2_X1 U2710 ( .A(\REGISTERS[19][1] ), .B(n3038), .S(n24), .Z(n1525) );
  MUX2_X1 U2711 ( .A(\REGISTERS[19][0] ), .B(n3039), .S(n24), .Z(n1524) );
  OAI21_X1 U2712 ( .B1(n3048), .B2(n3070), .A(n3042), .ZN(n3073) );
  MUX2_X1 U2713 ( .A(\REGISTERS[20][31] ), .B(n3007), .S(n26), .Z(n1523) );
  MUX2_X1 U2714 ( .A(\REGISTERS[20][30] ), .B(n3009), .S(n26), .Z(n1522) );
  MUX2_X1 U2715 ( .A(\REGISTERS[20][29] ), .B(n3010), .S(n26), .Z(n1521) );
  MUX2_X1 U2716 ( .A(\REGISTERS[20][28] ), .B(n3011), .S(n26), .Z(n1520) );
  MUX2_X1 U2717 ( .A(\REGISTERS[20][27] ), .B(n3012), .S(n26), .Z(n1519) );
  MUX2_X1 U2718 ( .A(\REGISTERS[20][26] ), .B(n3013), .S(n26), .Z(n1518) );
  MUX2_X1 U2719 ( .A(\REGISTERS[20][25] ), .B(n3014), .S(n26), .Z(n1517) );
  MUX2_X1 U2720 ( .A(\REGISTERS[20][24] ), .B(n3015), .S(n26), .Z(n1516) );
  MUX2_X1 U2721 ( .A(\REGISTERS[20][23] ), .B(n3016), .S(n26), .Z(n1515) );
  MUX2_X1 U2722 ( .A(\REGISTERS[20][22] ), .B(n3017), .S(n26), .Z(n1514) );
  MUX2_X1 U2723 ( .A(\REGISTERS[20][21] ), .B(n3018), .S(n26), .Z(n1513) );
  MUX2_X1 U2724 ( .A(\REGISTERS[20][20] ), .B(n3019), .S(n26), .Z(n1512) );
  MUX2_X1 U2725 ( .A(\REGISTERS[20][19] ), .B(n3020), .S(n26), .Z(n1511) );
  MUX2_X1 U2726 ( .A(\REGISTERS[20][18] ), .B(n3021), .S(n26), .Z(n1510) );
  MUX2_X1 U2727 ( .A(\REGISTERS[20][17] ), .B(n3022), .S(n26), .Z(n1509) );
  MUX2_X1 U2728 ( .A(\REGISTERS[20][16] ), .B(n3023), .S(n26), .Z(n1508) );
  MUX2_X1 U2729 ( .A(\REGISTERS[20][15] ), .B(n3024), .S(n26), .Z(n1507) );
  MUX2_X1 U2730 ( .A(\REGISTERS[20][14] ), .B(n3025), .S(n26), .Z(n1506) );
  MUX2_X1 U2731 ( .A(\REGISTERS[20][13] ), .B(n3026), .S(n26), .Z(n1505) );
  MUX2_X1 U2732 ( .A(\REGISTERS[20][12] ), .B(n3027), .S(n26), .Z(n1504) );
  MUX2_X1 U2733 ( .A(\REGISTERS[20][11] ), .B(n3028), .S(n26), .Z(n1503) );
  MUX2_X1 U2734 ( .A(\REGISTERS[20][10] ), .B(n3029), .S(n26), .Z(n1502) );
  MUX2_X1 U2735 ( .A(\REGISTERS[20][9] ), .B(n3030), .S(n26), .Z(n1501) );
  MUX2_X1 U2736 ( .A(\REGISTERS[20][8] ), .B(n3031), .S(n26), .Z(n1500) );
  MUX2_X1 U2737 ( .A(\REGISTERS[20][7] ), .B(n3032), .S(n26), .Z(n1499) );
  MUX2_X1 U2738 ( .A(\REGISTERS[20][6] ), .B(n3033), .S(n26), .Z(n1498) );
  MUX2_X1 U2739 ( .A(\REGISTERS[20][5] ), .B(n3034), .S(n26), .Z(n1497) );
  MUX2_X1 U2740 ( .A(\REGISTERS[20][4] ), .B(n3035), .S(n26), .Z(n1496) );
  MUX2_X1 U2741 ( .A(\REGISTERS[20][3] ), .B(n3036), .S(n26), .Z(n1495) );
  MUX2_X1 U2742 ( .A(\REGISTERS[20][2] ), .B(n3037), .S(n26), .Z(n1494) );
  MUX2_X1 U2743 ( .A(\REGISTERS[20][1] ), .B(n3038), .S(n26), .Z(n1493) );
  MUX2_X1 U2744 ( .A(\REGISTERS[20][0] ), .B(n3039), .S(n26), .Z(n1492) );
  OAI21_X1 U2745 ( .B1(n3050), .B2(n3070), .A(n3042), .ZN(n3074) );
  MUX2_X1 U2746 ( .A(\REGISTERS[21][31] ), .B(n3007), .S(n20), .Z(n1491) );
  MUX2_X1 U2747 ( .A(\REGISTERS[21][30] ), .B(n3009), .S(n20), .Z(n1490) );
  MUX2_X1 U2748 ( .A(\REGISTERS[21][29] ), .B(n3010), .S(n20), .Z(n1489) );
  MUX2_X1 U2749 ( .A(\REGISTERS[21][28] ), .B(n3011), .S(n20), .Z(n1488) );
  MUX2_X1 U2750 ( .A(\REGISTERS[21][27] ), .B(n3012), .S(n20), .Z(n1487) );
  MUX2_X1 U2751 ( .A(\REGISTERS[21][26] ), .B(n3013), .S(n20), .Z(n1486) );
  MUX2_X1 U2752 ( .A(\REGISTERS[21][25] ), .B(n3014), .S(n20), .Z(n1485) );
  MUX2_X1 U2753 ( .A(\REGISTERS[21][24] ), .B(n3015), .S(n20), .Z(n1484) );
  MUX2_X1 U2754 ( .A(\REGISTERS[21][23] ), .B(n3016), .S(n20), .Z(n1483) );
  MUX2_X1 U2755 ( .A(\REGISTERS[21][22] ), .B(n3017), .S(n20), .Z(n1482) );
  MUX2_X1 U2756 ( .A(\REGISTERS[21][21] ), .B(n3018), .S(n20), .Z(n1481) );
  MUX2_X1 U2757 ( .A(\REGISTERS[21][20] ), .B(n3019), .S(n20), .Z(n1480) );
  MUX2_X1 U2758 ( .A(\REGISTERS[21][19] ), .B(n3020), .S(n20), .Z(n1479) );
  MUX2_X1 U2759 ( .A(\REGISTERS[21][18] ), .B(n3021), .S(n20), .Z(n1478) );
  MUX2_X1 U2760 ( .A(\REGISTERS[21][17] ), .B(n3022), .S(n20), .Z(n1477) );
  MUX2_X1 U2761 ( .A(\REGISTERS[21][16] ), .B(n3023), .S(n20), .Z(n1476) );
  MUX2_X1 U2762 ( .A(\REGISTERS[21][15] ), .B(n3024), .S(n20), .Z(n1475) );
  MUX2_X1 U2763 ( .A(\REGISTERS[21][14] ), .B(n3025), .S(n20), .Z(n1474) );
  MUX2_X1 U2764 ( .A(\REGISTERS[21][13] ), .B(n3026), .S(n20), .Z(n1473) );
  MUX2_X1 U2765 ( .A(\REGISTERS[21][12] ), .B(n3027), .S(n20), .Z(n1472) );
  MUX2_X1 U2766 ( .A(\REGISTERS[21][11] ), .B(n3028), .S(n20), .Z(n1471) );
  MUX2_X1 U2767 ( .A(\REGISTERS[21][10] ), .B(n3029), .S(n20), .Z(n1470) );
  MUX2_X1 U2768 ( .A(\REGISTERS[21][9] ), .B(n3030), .S(n20), .Z(n1469) );
  MUX2_X1 U2769 ( .A(\REGISTERS[21][8] ), .B(n3031), .S(n20), .Z(n1468) );
  MUX2_X1 U2770 ( .A(\REGISTERS[21][7] ), .B(n3032), .S(n20), .Z(n1467) );
  MUX2_X1 U2771 ( .A(\REGISTERS[21][6] ), .B(n3033), .S(n20), .Z(n1466) );
  MUX2_X1 U2772 ( .A(\REGISTERS[21][5] ), .B(n3034), .S(n20), .Z(n1465) );
  MUX2_X1 U2773 ( .A(\REGISTERS[21][4] ), .B(n3035), .S(n20), .Z(n1464) );
  MUX2_X1 U2774 ( .A(\REGISTERS[21][3] ), .B(n3036), .S(n20), .Z(n1463) );
  MUX2_X1 U2775 ( .A(\REGISTERS[21][2] ), .B(n3037), .S(n20), .Z(n1462) );
  MUX2_X1 U2776 ( .A(\REGISTERS[21][1] ), .B(n3038), .S(n20), .Z(n1461) );
  MUX2_X1 U2777 ( .A(\REGISTERS[21][0] ), .B(n3039), .S(n20), .Z(n1460) );
  OAI21_X1 U2778 ( .B1(n3052), .B2(n3070), .A(n3042), .ZN(n3075) );
  MUX2_X1 U2779 ( .A(\REGISTERS[22][31] ), .B(n3007), .S(n22), .Z(n1459) );
  MUX2_X1 U2780 ( .A(\REGISTERS[22][30] ), .B(n3009), .S(n22), .Z(n1458) );
  MUX2_X1 U2781 ( .A(\REGISTERS[22][29] ), .B(n3010), .S(n22), .Z(n1457) );
  MUX2_X1 U2782 ( .A(\REGISTERS[22][28] ), .B(n3011), .S(n22), .Z(n1456) );
  MUX2_X1 U2783 ( .A(\REGISTERS[22][27] ), .B(n3012), .S(n22), .Z(n1455) );
  MUX2_X1 U2784 ( .A(\REGISTERS[22][26] ), .B(n3013), .S(n22), .Z(n1454) );
  MUX2_X1 U2785 ( .A(\REGISTERS[22][25] ), .B(n3014), .S(n22), .Z(n1453) );
  MUX2_X1 U2786 ( .A(\REGISTERS[22][24] ), .B(n3015), .S(n22), .Z(n1452) );
  MUX2_X1 U2787 ( .A(\REGISTERS[22][23] ), .B(n3016), .S(n22), .Z(n1451) );
  MUX2_X1 U2788 ( .A(\REGISTERS[22][22] ), .B(n3017), .S(n22), .Z(n1450) );
  MUX2_X1 U2789 ( .A(\REGISTERS[22][21] ), .B(n3018), .S(n22), .Z(n1449) );
  MUX2_X1 U2790 ( .A(\REGISTERS[22][20] ), .B(n3019), .S(n22), .Z(n1448) );
  MUX2_X1 U2791 ( .A(\REGISTERS[22][19] ), .B(n3020), .S(n22), .Z(n1447) );
  MUX2_X1 U2792 ( .A(\REGISTERS[22][18] ), .B(n3021), .S(n22), .Z(n1446) );
  MUX2_X1 U2793 ( .A(\REGISTERS[22][17] ), .B(n3022), .S(n22), .Z(n1445) );
  MUX2_X1 U2794 ( .A(\REGISTERS[22][16] ), .B(n3023), .S(n22), .Z(n1444) );
  MUX2_X1 U2795 ( .A(\REGISTERS[22][15] ), .B(n3024), .S(n22), .Z(n1443) );
  MUX2_X1 U2796 ( .A(\REGISTERS[22][14] ), .B(n3025), .S(n22), .Z(n1442) );
  MUX2_X1 U2797 ( .A(\REGISTERS[22][13] ), .B(n3026), .S(n22), .Z(n1441) );
  MUX2_X1 U2798 ( .A(\REGISTERS[22][12] ), .B(n3027), .S(n22), .Z(n1440) );
  MUX2_X1 U2799 ( .A(\REGISTERS[22][11] ), .B(n3028), .S(n22), .Z(n1439) );
  MUX2_X1 U2800 ( .A(\REGISTERS[22][10] ), .B(n3029), .S(n22), .Z(n1438) );
  MUX2_X1 U2801 ( .A(\REGISTERS[22][9] ), .B(n3030), .S(n22), .Z(n1437) );
  MUX2_X1 U2802 ( .A(\REGISTERS[22][8] ), .B(n3031), .S(n22), .Z(n1436) );
  MUX2_X1 U2803 ( .A(\REGISTERS[22][7] ), .B(n3032), .S(n22), .Z(n1435) );
  MUX2_X1 U2804 ( .A(\REGISTERS[22][6] ), .B(n3033), .S(n22), .Z(n1434) );
  MUX2_X1 U2805 ( .A(\REGISTERS[22][5] ), .B(n3034), .S(n22), .Z(n1433) );
  MUX2_X1 U2806 ( .A(\REGISTERS[22][4] ), .B(n3035), .S(n22), .Z(n1432) );
  MUX2_X1 U2807 ( .A(\REGISTERS[22][3] ), .B(n3036), .S(n22), .Z(n1431) );
  MUX2_X1 U2808 ( .A(\REGISTERS[22][2] ), .B(n3037), .S(n22), .Z(n1430) );
  MUX2_X1 U2809 ( .A(\REGISTERS[22][1] ), .B(n3038), .S(n22), .Z(n1429) );
  MUX2_X1 U2810 ( .A(\REGISTERS[22][0] ), .B(n3039), .S(n22), .Z(n1428) );
  OAI21_X1 U2811 ( .B1(n3054), .B2(n3070), .A(n3042), .ZN(n3076) );
  MUX2_X1 U2812 ( .A(\REGISTERS[23][31] ), .B(n3007), .S(n16), .Z(n1427) );
  MUX2_X1 U2813 ( .A(\REGISTERS[23][30] ), .B(n3009), .S(n16), .Z(n1426) );
  MUX2_X1 U2814 ( .A(\REGISTERS[23][29] ), .B(n3010), .S(n16), .Z(n1425) );
  MUX2_X1 U2815 ( .A(\REGISTERS[23][28] ), .B(n3011), .S(n16), .Z(n1424) );
  MUX2_X1 U2816 ( .A(\REGISTERS[23][27] ), .B(n3012), .S(n16), .Z(n1423) );
  MUX2_X1 U2817 ( .A(\REGISTERS[23][26] ), .B(n3013), .S(n16), .Z(n1422) );
  MUX2_X1 U2818 ( .A(\REGISTERS[23][25] ), .B(n3014), .S(n16), .Z(n1421) );
  MUX2_X1 U2819 ( .A(\REGISTERS[23][24] ), .B(n3015), .S(n16), .Z(n1420) );
  MUX2_X1 U2820 ( .A(\REGISTERS[23][23] ), .B(n3016), .S(n16), .Z(n1419) );
  MUX2_X1 U2821 ( .A(\REGISTERS[23][22] ), .B(n3017), .S(n16), .Z(n1418) );
  MUX2_X1 U2822 ( .A(\REGISTERS[23][21] ), .B(n3018), .S(n16), .Z(n1417) );
  MUX2_X1 U2823 ( .A(\REGISTERS[23][20] ), .B(n3019), .S(n16), .Z(n1416) );
  MUX2_X1 U2824 ( .A(\REGISTERS[23][19] ), .B(n3020), .S(n16), .Z(n1415) );
  MUX2_X1 U2825 ( .A(\REGISTERS[23][18] ), .B(n3021), .S(n16), .Z(n1414) );
  MUX2_X1 U2826 ( .A(\REGISTERS[23][17] ), .B(n3022), .S(n16), .Z(n1413) );
  MUX2_X1 U2827 ( .A(\REGISTERS[23][16] ), .B(n3023), .S(n16), .Z(n1412) );
  MUX2_X1 U2828 ( .A(\REGISTERS[23][15] ), .B(n3024), .S(n16), .Z(n1411) );
  MUX2_X1 U2829 ( .A(\REGISTERS[23][14] ), .B(n3025), .S(n16), .Z(n1410) );
  MUX2_X1 U2830 ( .A(\REGISTERS[23][13] ), .B(n3026), .S(n16), .Z(n1409) );
  MUX2_X1 U2831 ( .A(\REGISTERS[23][12] ), .B(n3027), .S(n16), .Z(n1408) );
  MUX2_X1 U2832 ( .A(\REGISTERS[23][11] ), .B(n3028), .S(n16), .Z(n1407) );
  MUX2_X1 U2833 ( .A(\REGISTERS[23][10] ), .B(n3029), .S(n16), .Z(n1406) );
  MUX2_X1 U2834 ( .A(\REGISTERS[23][9] ), .B(n3030), .S(n16), .Z(n1405) );
  MUX2_X1 U2835 ( .A(\REGISTERS[23][8] ), .B(n3031), .S(n16), .Z(n1404) );
  MUX2_X1 U2836 ( .A(\REGISTERS[23][7] ), .B(n3032), .S(n16), .Z(n1403) );
  MUX2_X1 U2837 ( .A(\REGISTERS[23][6] ), .B(n3033), .S(n16), .Z(n1402) );
  MUX2_X1 U2838 ( .A(\REGISTERS[23][5] ), .B(n3034), .S(n16), .Z(n1401) );
  MUX2_X1 U2839 ( .A(\REGISTERS[23][4] ), .B(n3035), .S(n16), .Z(n1400) );
  MUX2_X1 U2840 ( .A(\REGISTERS[23][3] ), .B(n3036), .S(n16), .Z(n1399) );
  MUX2_X1 U2841 ( .A(\REGISTERS[23][2] ), .B(n3037), .S(n16), .Z(n1398) );
  MUX2_X1 U2842 ( .A(\REGISTERS[23][1] ), .B(n3038), .S(n16), .Z(n1397) );
  MUX2_X1 U2843 ( .A(\REGISTERS[23][0] ), .B(n3039), .S(n16), .Z(n1396) );
  OAI21_X1 U2844 ( .B1(n3056), .B2(n3070), .A(n3042), .ZN(n3077) );
  NAND3_X1 U2845 ( .A1(n3059), .A2(n3057), .A3(ADD_WR[4]), .ZN(n3070) );
  INV_X1 U2846 ( .A(ADD_WR[3]), .ZN(n3057) );
  MUX2_X1 U2847 ( .A(\REGISTERS[24][31] ), .B(n3007), .S(n18), .Z(n1395) );
  MUX2_X1 U2848 ( .A(\REGISTERS[24][30] ), .B(n3009), .S(n18), .Z(n1394) );
  MUX2_X1 U2849 ( .A(\REGISTERS[24][29] ), .B(n3010), .S(n18), .Z(n1393) );
  MUX2_X1 U2850 ( .A(\REGISTERS[24][28] ), .B(n3011), .S(n18), .Z(n1392) );
  MUX2_X1 U2851 ( .A(\REGISTERS[24][27] ), .B(n3012), .S(n18), .Z(n1391) );
  MUX2_X1 U2852 ( .A(\REGISTERS[24][26] ), .B(n3013), .S(n18), .Z(n1390) );
  MUX2_X1 U2853 ( .A(\REGISTERS[24][25] ), .B(n3014), .S(n18), .Z(n1389) );
  MUX2_X1 U2854 ( .A(\REGISTERS[24][24] ), .B(n3015), .S(n18), .Z(n1388) );
  MUX2_X1 U2855 ( .A(\REGISTERS[24][23] ), .B(n3016), .S(n18), .Z(n1387) );
  MUX2_X1 U2856 ( .A(\REGISTERS[24][22] ), .B(n3017), .S(n18), .Z(n1386) );
  MUX2_X1 U2857 ( .A(\REGISTERS[24][21] ), .B(n3018), .S(n18), .Z(n1385) );
  MUX2_X1 U2858 ( .A(\REGISTERS[24][20] ), .B(n3019), .S(n18), .Z(n1384) );
  MUX2_X1 U2859 ( .A(\REGISTERS[24][19] ), .B(n3020), .S(n18), .Z(n1383) );
  MUX2_X1 U2860 ( .A(\REGISTERS[24][18] ), .B(n3021), .S(n18), .Z(n1382) );
  MUX2_X1 U2861 ( .A(\REGISTERS[24][17] ), .B(n3022), .S(n18), .Z(n1381) );
  MUX2_X1 U2862 ( .A(\REGISTERS[24][16] ), .B(n3023), .S(n18), .Z(n1380) );
  MUX2_X1 U2863 ( .A(\REGISTERS[24][15] ), .B(n3024), .S(n18), .Z(n1379) );
  MUX2_X1 U2864 ( .A(\REGISTERS[24][14] ), .B(n3025), .S(n18), .Z(n1378) );
  MUX2_X1 U2865 ( .A(\REGISTERS[24][13] ), .B(n3026), .S(n18), .Z(n1377) );
  MUX2_X1 U2866 ( .A(\REGISTERS[24][12] ), .B(n3027), .S(n18), .Z(n1376) );
  MUX2_X1 U2867 ( .A(\REGISTERS[24][11] ), .B(n3028), .S(n18), .Z(n1375) );
  MUX2_X1 U2868 ( .A(\REGISTERS[24][10] ), .B(n3029), .S(n18), .Z(n1374) );
  MUX2_X1 U2869 ( .A(\REGISTERS[24][9] ), .B(n3030), .S(n18), .Z(n1373) );
  MUX2_X1 U2870 ( .A(\REGISTERS[24][8] ), .B(n3031), .S(n18), .Z(n1372) );
  MUX2_X1 U2871 ( .A(\REGISTERS[24][7] ), .B(n3032), .S(n18), .Z(n1371) );
  MUX2_X1 U2872 ( .A(\REGISTERS[24][6] ), .B(n3033), .S(n18), .Z(n1370) );
  MUX2_X1 U2873 ( .A(\REGISTERS[24][5] ), .B(n3034), .S(n18), .Z(n1369) );
  MUX2_X1 U2874 ( .A(\REGISTERS[24][4] ), .B(n3035), .S(n18), .Z(n1368) );
  MUX2_X1 U2875 ( .A(\REGISTERS[24][3] ), .B(n3036), .S(n18), .Z(n1367) );
  MUX2_X1 U2876 ( .A(\REGISTERS[24][2] ), .B(n3037), .S(n18), .Z(n1366) );
  MUX2_X1 U2877 ( .A(\REGISTERS[24][1] ), .B(n3038), .S(n18), .Z(n1365) );
  MUX2_X1 U2878 ( .A(\REGISTERS[24][0] ), .B(n3039), .S(n18), .Z(n1364) );
  OAI21_X1 U2879 ( .B1(n3041), .B2(n3079), .A(n3042), .ZN(n3078) );
  NAND3_X1 U2880 ( .A1(n3080), .A2(n3081), .A3(n3082), .ZN(n3041) );
  MUX2_X1 U2881 ( .A(\REGISTERS[25][31] ), .B(n3007), .S(n2), .Z(n1363) );
  MUX2_X1 U2882 ( .A(\REGISTERS[25][30] ), .B(n3009), .S(n2), .Z(n1362) );
  MUX2_X1 U2883 ( .A(\REGISTERS[25][29] ), .B(n3010), .S(n2), .Z(n1361) );
  MUX2_X1 U2884 ( .A(\REGISTERS[25][28] ), .B(n3011), .S(n2), .Z(n1360) );
  MUX2_X1 U2885 ( .A(\REGISTERS[25][27] ), .B(n3012), .S(n2), .Z(n1359) );
  MUX2_X1 U2886 ( .A(\REGISTERS[25][26] ), .B(n3013), .S(n2), .Z(n1358) );
  MUX2_X1 U2887 ( .A(\REGISTERS[25][25] ), .B(n3014), .S(n2), .Z(n1357) );
  MUX2_X1 U2888 ( .A(\REGISTERS[25][24] ), .B(n3015), .S(n2), .Z(n1356) );
  MUX2_X1 U2889 ( .A(\REGISTERS[25][23] ), .B(n3016), .S(n2), .Z(n1355) );
  MUX2_X1 U2890 ( .A(\REGISTERS[25][22] ), .B(n3017), .S(n2), .Z(n1354) );
  MUX2_X1 U2891 ( .A(\REGISTERS[25][21] ), .B(n3018), .S(n2), .Z(n1353) );
  MUX2_X1 U2892 ( .A(\REGISTERS[25][20] ), .B(n3019), .S(n2), .Z(n1352) );
  MUX2_X1 U2893 ( .A(\REGISTERS[25][19] ), .B(n3020), .S(n2), .Z(n1351) );
  MUX2_X1 U2894 ( .A(\REGISTERS[25][18] ), .B(n3021), .S(n2), .Z(n1350) );
  MUX2_X1 U2895 ( .A(\REGISTERS[25][17] ), .B(n3022), .S(n2), .Z(n1349) );
  MUX2_X1 U2896 ( .A(\REGISTERS[25][16] ), .B(n3023), .S(n2), .Z(n1348) );
  MUX2_X1 U2897 ( .A(\REGISTERS[25][15] ), .B(n3024), .S(n2), .Z(n1347) );
  MUX2_X1 U2898 ( .A(\REGISTERS[25][14] ), .B(n3025), .S(n2), .Z(n1346) );
  MUX2_X1 U2899 ( .A(\REGISTERS[25][13] ), .B(n3026), .S(n2), .Z(n1345) );
  MUX2_X1 U2900 ( .A(\REGISTERS[25][12] ), .B(n3027), .S(n2), .Z(n1344) );
  MUX2_X1 U2901 ( .A(\REGISTERS[25][11] ), .B(n3028), .S(n2), .Z(n1343) );
  MUX2_X1 U2902 ( .A(\REGISTERS[25][10] ), .B(n3029), .S(n2), .Z(n1342) );
  MUX2_X1 U2903 ( .A(\REGISTERS[25][9] ), .B(n3030), .S(n2), .Z(n1341) );
  MUX2_X1 U2904 ( .A(\REGISTERS[25][8] ), .B(n3031), .S(n2), .Z(n1340) );
  MUX2_X1 U2905 ( .A(\REGISTERS[25][7] ), .B(n3032), .S(n2), .Z(n1339) );
  MUX2_X1 U2906 ( .A(\REGISTERS[25][6] ), .B(n3033), .S(n2), .Z(n1338) );
  MUX2_X1 U2907 ( .A(\REGISTERS[25][5] ), .B(n3034), .S(n2), .Z(n1337) );
  MUX2_X1 U2908 ( .A(\REGISTERS[25][4] ), .B(n3035), .S(n2), .Z(n1336) );
  MUX2_X1 U2909 ( .A(\REGISTERS[25][3] ), .B(n3036), .S(n2), .Z(n1335) );
  MUX2_X1 U2910 ( .A(\REGISTERS[25][2] ), .B(n3037), .S(n2), .Z(n1334) );
  MUX2_X1 U2911 ( .A(\REGISTERS[25][1] ), .B(n3038), .S(n2), .Z(n1333) );
  MUX2_X1 U2912 ( .A(\REGISTERS[25][0] ), .B(n3039), .S(n2), .Z(n1332) );
  OAI21_X1 U2913 ( .B1(n3044), .B2(n3079), .A(n3042), .ZN(n3083) );
  NAND3_X1 U2914 ( .A1(n3080), .A2(n3081), .A3(ADD_WR[0]), .ZN(n3044) );
  MUX2_X1 U2915 ( .A(\REGISTERS[26][31] ), .B(n3007), .S(n4), .Z(n1331) );
  MUX2_X1 U2916 ( .A(\REGISTERS[26][30] ), .B(n3009), .S(n4), .Z(n1330) );
  MUX2_X1 U2917 ( .A(\REGISTERS[26][29] ), .B(n3010), .S(n4), .Z(n1329) );
  MUX2_X1 U2918 ( .A(\REGISTERS[26][28] ), .B(n3011), .S(n4), .Z(n1328) );
  MUX2_X1 U2919 ( .A(\REGISTERS[26][27] ), .B(n3012), .S(n4), .Z(n1327) );
  MUX2_X1 U2920 ( .A(\REGISTERS[26][26] ), .B(n3013), .S(n4), .Z(n1326) );
  MUX2_X1 U2921 ( .A(\REGISTERS[26][25] ), .B(n3014), .S(n4), .Z(n1325) );
  MUX2_X1 U2922 ( .A(\REGISTERS[26][24] ), .B(n3015), .S(n4), .Z(n1324) );
  MUX2_X1 U2923 ( .A(\REGISTERS[26][23] ), .B(n3016), .S(n4), .Z(n1323) );
  MUX2_X1 U2924 ( .A(\REGISTERS[26][22] ), .B(n3017), .S(n4), .Z(n1322) );
  MUX2_X1 U2925 ( .A(\REGISTERS[26][21] ), .B(n3018), .S(n4), .Z(n1321) );
  MUX2_X1 U2926 ( .A(\REGISTERS[26][20] ), .B(n3019), .S(n4), .Z(n1320) );
  MUX2_X1 U2927 ( .A(\REGISTERS[26][19] ), .B(n3020), .S(n4), .Z(n1319) );
  MUX2_X1 U2928 ( .A(\REGISTERS[26][18] ), .B(n3021), .S(n4), .Z(n1318) );
  MUX2_X1 U2929 ( .A(\REGISTERS[26][17] ), .B(n3022), .S(n4), .Z(n1317) );
  MUX2_X1 U2930 ( .A(\REGISTERS[26][16] ), .B(n3023), .S(n4), .Z(n1316) );
  MUX2_X1 U2931 ( .A(\REGISTERS[26][15] ), .B(n3024), .S(n4), .Z(n1315) );
  MUX2_X1 U2932 ( .A(\REGISTERS[26][14] ), .B(n3025), .S(n4), .Z(n1314) );
  MUX2_X1 U2933 ( .A(\REGISTERS[26][13] ), .B(n3026), .S(n4), .Z(n1313) );
  MUX2_X1 U2934 ( .A(\REGISTERS[26][12] ), .B(n3027), .S(n4), .Z(n1312) );
  MUX2_X1 U2935 ( .A(\REGISTERS[26][11] ), .B(n3028), .S(n4), .Z(n1311) );
  MUX2_X1 U2936 ( .A(\REGISTERS[26][10] ), .B(n3029), .S(n4), .Z(n1310) );
  MUX2_X1 U2937 ( .A(\REGISTERS[26][9] ), .B(n3030), .S(n4), .Z(n1309) );
  MUX2_X1 U2938 ( .A(\REGISTERS[26][8] ), .B(n3031), .S(n4), .Z(n1308) );
  MUX2_X1 U2939 ( .A(\REGISTERS[26][7] ), .B(n3032), .S(n4), .Z(n1307) );
  MUX2_X1 U2940 ( .A(\REGISTERS[26][6] ), .B(n3033), .S(n4), .Z(n1306) );
  MUX2_X1 U2941 ( .A(\REGISTERS[26][5] ), .B(n3034), .S(n4), .Z(n1305) );
  MUX2_X1 U2942 ( .A(\REGISTERS[26][4] ), .B(n3035), .S(n4), .Z(n1304) );
  MUX2_X1 U2943 ( .A(\REGISTERS[26][3] ), .B(n3036), .S(n4), .Z(n1303) );
  MUX2_X1 U2944 ( .A(\REGISTERS[26][2] ), .B(n3037), .S(n4), .Z(n1302) );
  MUX2_X1 U2945 ( .A(\REGISTERS[26][1] ), .B(n3038), .S(n4), .Z(n1301) );
  MUX2_X1 U2946 ( .A(\REGISTERS[26][0] ), .B(n3039), .S(n4), .Z(n1300) );
  OAI21_X1 U2947 ( .B1(n3046), .B2(n3079), .A(n3042), .ZN(n3084) );
  NAND3_X1 U2948 ( .A1(n3082), .A2(n3081), .A3(ADD_WR[1]), .ZN(n3046) );
  MUX2_X1 U2949 ( .A(\REGISTERS[27][31] ), .B(n3007), .S(n6), .Z(n1299) );
  MUX2_X1 U2950 ( .A(\REGISTERS[27][30] ), .B(n3009), .S(n6), .Z(n1298) );
  MUX2_X1 U2951 ( .A(\REGISTERS[27][29] ), .B(n3010), .S(n6), .Z(n1297) );
  MUX2_X1 U2952 ( .A(\REGISTERS[27][28] ), .B(n3011), .S(n6), .Z(n1296) );
  MUX2_X1 U2953 ( .A(\REGISTERS[27][27] ), .B(n3012), .S(n6), .Z(n1295) );
  MUX2_X1 U2954 ( .A(\REGISTERS[27][26] ), .B(n3013), .S(n6), .Z(n1294) );
  MUX2_X1 U2955 ( .A(\REGISTERS[27][25] ), .B(n3014), .S(n6), .Z(n1293) );
  MUX2_X1 U2956 ( .A(\REGISTERS[27][24] ), .B(n3015), .S(n6), .Z(n1292) );
  MUX2_X1 U2957 ( .A(\REGISTERS[27][23] ), .B(n3016), .S(n6), .Z(n1291) );
  MUX2_X1 U2958 ( .A(\REGISTERS[27][22] ), .B(n3017), .S(n6), .Z(n1290) );
  MUX2_X1 U2959 ( .A(\REGISTERS[27][21] ), .B(n3018), .S(n6), .Z(n1289) );
  MUX2_X1 U2960 ( .A(\REGISTERS[27][20] ), .B(n3019), .S(n6), .Z(n1288) );
  MUX2_X1 U2961 ( .A(\REGISTERS[27][19] ), .B(n3020), .S(n6), .Z(n1287) );
  MUX2_X1 U2962 ( .A(\REGISTERS[27][18] ), .B(n3021), .S(n6), .Z(n1286) );
  MUX2_X1 U2963 ( .A(\REGISTERS[27][17] ), .B(n3022), .S(n6), .Z(n1285) );
  MUX2_X1 U2964 ( .A(\REGISTERS[27][16] ), .B(n3023), .S(n6), .Z(n1284) );
  MUX2_X1 U2965 ( .A(\REGISTERS[27][15] ), .B(n3024), .S(n6), .Z(n1283) );
  MUX2_X1 U2966 ( .A(\REGISTERS[27][14] ), .B(n3025), .S(n6), .Z(n1282) );
  MUX2_X1 U2967 ( .A(\REGISTERS[27][13] ), .B(n3026), .S(n6), .Z(n1281) );
  MUX2_X1 U2968 ( .A(\REGISTERS[27][12] ), .B(n3027), .S(n6), .Z(n1280) );
  MUX2_X1 U2969 ( .A(\REGISTERS[27][11] ), .B(n3028), .S(n6), .Z(n1279) );
  MUX2_X1 U2970 ( .A(\REGISTERS[27][10] ), .B(n3029), .S(n6), .Z(n1278) );
  MUX2_X1 U2971 ( .A(\REGISTERS[27][9] ), .B(n3030), .S(n6), .Z(n1277) );
  MUX2_X1 U2972 ( .A(\REGISTERS[27][8] ), .B(n3031), .S(n6), .Z(n1276) );
  MUX2_X1 U2973 ( .A(\REGISTERS[27][7] ), .B(n3032), .S(n6), .Z(n1275) );
  MUX2_X1 U2974 ( .A(\REGISTERS[27][6] ), .B(n3033), .S(n6), .Z(n1274) );
  MUX2_X1 U2975 ( .A(\REGISTERS[27][5] ), .B(n3034), .S(n6), .Z(n1273) );
  MUX2_X1 U2976 ( .A(\REGISTERS[27][4] ), .B(n3035), .S(n6), .Z(n1272) );
  MUX2_X1 U2977 ( .A(\REGISTERS[27][3] ), .B(n3036), .S(n6), .Z(n1271) );
  MUX2_X1 U2978 ( .A(\REGISTERS[27][2] ), .B(n3037), .S(n6), .Z(n1270) );
  MUX2_X1 U2979 ( .A(\REGISTERS[27][1] ), .B(n3038), .S(n6), .Z(n1269) );
  MUX2_X1 U2980 ( .A(\REGISTERS[27][0] ), .B(n3039), .S(n6), .Z(n1268) );
  OAI21_X1 U2981 ( .B1(n3048), .B2(n3079), .A(n3042), .ZN(n3085) );
  NAND3_X1 U2982 ( .A1(ADD_WR[0]), .A2(n3081), .A3(ADD_WR[1]), .ZN(n3048) );
  INV_X1 U2983 ( .A(ADD_WR[2]), .ZN(n3081) );
  MUX2_X1 U2984 ( .A(\REGISTERS[28][31] ), .B(n3007), .S(n8), .Z(n1267) );
  MUX2_X1 U2985 ( .A(\REGISTERS[28][30] ), .B(n3009), .S(n8), .Z(n1266) );
  MUX2_X1 U2986 ( .A(\REGISTERS[28][29] ), .B(n3010), .S(n8), .Z(n1265) );
  MUX2_X1 U2987 ( .A(\REGISTERS[28][28] ), .B(n3011), .S(n8), .Z(n1264) );
  MUX2_X1 U2988 ( .A(\REGISTERS[28][27] ), .B(n3012), .S(n8), .Z(n1263) );
  MUX2_X1 U2989 ( .A(\REGISTERS[28][26] ), .B(n3013), .S(n8), .Z(n1262) );
  MUX2_X1 U2990 ( .A(\REGISTERS[28][25] ), .B(n3014), .S(n8), .Z(n1261) );
  MUX2_X1 U2991 ( .A(\REGISTERS[28][24] ), .B(n3015), .S(n8), .Z(n1260) );
  MUX2_X1 U2992 ( .A(\REGISTERS[28][23] ), .B(n3016), .S(n8), .Z(n1259) );
  MUX2_X1 U2993 ( .A(\REGISTERS[28][22] ), .B(n3017), .S(n8), .Z(n1258) );
  MUX2_X1 U2994 ( .A(\REGISTERS[28][21] ), .B(n3018), .S(n8), .Z(n1257) );
  MUX2_X1 U2995 ( .A(\REGISTERS[28][20] ), .B(n3019), .S(n8), .Z(n1256) );
  MUX2_X1 U2996 ( .A(\REGISTERS[28][19] ), .B(n3020), .S(n8), .Z(n1255) );
  MUX2_X1 U2997 ( .A(\REGISTERS[28][18] ), .B(n3021), .S(n8), .Z(n1254) );
  MUX2_X1 U2998 ( .A(\REGISTERS[28][17] ), .B(n3022), .S(n8), .Z(n1253) );
  MUX2_X1 U2999 ( .A(\REGISTERS[28][16] ), .B(n3023), .S(n8), .Z(n1252) );
  MUX2_X1 U3000 ( .A(\REGISTERS[28][15] ), .B(n3024), .S(n8), .Z(n1251) );
  MUX2_X1 U3001 ( .A(\REGISTERS[28][14] ), .B(n3025), .S(n8), .Z(n1250) );
  MUX2_X1 U3002 ( .A(\REGISTERS[28][13] ), .B(n3026), .S(n8), .Z(n1249) );
  MUX2_X1 U3003 ( .A(\REGISTERS[28][12] ), .B(n3027), .S(n8), .Z(n1248) );
  MUX2_X1 U3004 ( .A(\REGISTERS[28][11] ), .B(n3028), .S(n8), .Z(n1247) );
  MUX2_X1 U3005 ( .A(\REGISTERS[28][10] ), .B(n3029), .S(n8), .Z(n1246) );
  MUX2_X1 U3006 ( .A(\REGISTERS[28][9] ), .B(n3030), .S(n8), .Z(n1245) );
  MUX2_X1 U3007 ( .A(\REGISTERS[28][8] ), .B(n3031), .S(n8), .Z(n1244) );
  MUX2_X1 U3008 ( .A(\REGISTERS[28][7] ), .B(n3032), .S(n8), .Z(n1243) );
  MUX2_X1 U3009 ( .A(\REGISTERS[28][6] ), .B(n3033), .S(n8), .Z(n1242) );
  MUX2_X1 U3010 ( .A(\REGISTERS[28][5] ), .B(n3034), .S(n8), .Z(n1241) );
  MUX2_X1 U3011 ( .A(\REGISTERS[28][4] ), .B(n3035), .S(n8), .Z(n1240) );
  MUX2_X1 U3012 ( .A(\REGISTERS[28][3] ), .B(n3036), .S(n8), .Z(n1239) );
  MUX2_X1 U3013 ( .A(\REGISTERS[28][2] ), .B(n3037), .S(n8), .Z(n1238) );
  MUX2_X1 U3014 ( .A(\REGISTERS[28][1] ), .B(n3038), .S(n8), .Z(n1237) );
  MUX2_X1 U3015 ( .A(\REGISTERS[28][0] ), .B(n3039), .S(n8), .Z(n1236) );
  OAI21_X1 U3016 ( .B1(n3050), .B2(n3079), .A(n3042), .ZN(n3086) );
  NAND3_X1 U3017 ( .A1(n3082), .A2(n3080), .A3(ADD_WR[2]), .ZN(n3050) );
  MUX2_X1 U3018 ( .A(\REGISTERS[29][31] ), .B(n3007), .S(n10), .Z(n1235) );
  MUX2_X1 U3019 ( .A(\REGISTERS[29][30] ), .B(n3009), .S(n10), .Z(n1234) );
  MUX2_X1 U3020 ( .A(\REGISTERS[29][29] ), .B(n3010), .S(n10), .Z(n1233) );
  MUX2_X1 U3021 ( .A(\REGISTERS[29][28] ), .B(n3011), .S(n10), .Z(n1232) );
  MUX2_X1 U3022 ( .A(\REGISTERS[29][27] ), .B(n3012), .S(n10), .Z(n1231) );
  MUX2_X1 U3023 ( .A(\REGISTERS[29][26] ), .B(n3013), .S(n10), .Z(n1230) );
  MUX2_X1 U3024 ( .A(\REGISTERS[29][25] ), .B(n3014), .S(n10), .Z(n1229) );
  MUX2_X1 U3025 ( .A(\REGISTERS[29][24] ), .B(n3015), .S(n10), .Z(n1228) );
  MUX2_X1 U3026 ( .A(\REGISTERS[29][23] ), .B(n3016), .S(n10), .Z(n1227) );
  MUX2_X1 U3027 ( .A(\REGISTERS[29][22] ), .B(n3017), .S(n10), .Z(n1226) );
  MUX2_X1 U3028 ( .A(\REGISTERS[29][21] ), .B(n3018), .S(n10), .Z(n1225) );
  MUX2_X1 U3029 ( .A(\REGISTERS[29][20] ), .B(n3019), .S(n10), .Z(n1224) );
  MUX2_X1 U3030 ( .A(\REGISTERS[29][19] ), .B(n3020), .S(n10), .Z(n1223) );
  MUX2_X1 U3031 ( .A(\REGISTERS[29][18] ), .B(n3021), .S(n10), .Z(n1222) );
  MUX2_X1 U3032 ( .A(\REGISTERS[29][17] ), .B(n3022), .S(n10), .Z(n1221) );
  MUX2_X1 U3033 ( .A(\REGISTERS[29][16] ), .B(n3023), .S(n10), .Z(n1220) );
  MUX2_X1 U3034 ( .A(\REGISTERS[29][15] ), .B(n3024), .S(n10), .Z(n1219) );
  MUX2_X1 U3035 ( .A(\REGISTERS[29][14] ), .B(n3025), .S(n10), .Z(n1218) );
  MUX2_X1 U3036 ( .A(\REGISTERS[29][13] ), .B(n3026), .S(n10), .Z(n1217) );
  MUX2_X1 U3037 ( .A(\REGISTERS[29][12] ), .B(n3027), .S(n10), .Z(n1216) );
  MUX2_X1 U3038 ( .A(\REGISTERS[29][11] ), .B(n3028), .S(n10), .Z(n1215) );
  MUX2_X1 U3039 ( .A(\REGISTERS[29][10] ), .B(n3029), .S(n10), .Z(n1214) );
  MUX2_X1 U3040 ( .A(\REGISTERS[29][9] ), .B(n3030), .S(n10), .Z(n1213) );
  MUX2_X1 U3041 ( .A(\REGISTERS[29][8] ), .B(n3031), .S(n10), .Z(n1212) );
  MUX2_X1 U3042 ( .A(\REGISTERS[29][7] ), .B(n3032), .S(n10), .Z(n1211) );
  MUX2_X1 U3043 ( .A(\REGISTERS[29][6] ), .B(n3033), .S(n10), .Z(n1210) );
  MUX2_X1 U3044 ( .A(\REGISTERS[29][5] ), .B(n3034), .S(n10), .Z(n1209) );
  MUX2_X1 U3045 ( .A(\REGISTERS[29][4] ), .B(n3035), .S(n10), .Z(n1208) );
  MUX2_X1 U3046 ( .A(\REGISTERS[29][3] ), .B(n3036), .S(n10), .Z(n1207) );
  MUX2_X1 U3047 ( .A(\REGISTERS[29][2] ), .B(n3037), .S(n10), .Z(n1206) );
  MUX2_X1 U3048 ( .A(\REGISTERS[29][1] ), .B(n3038), .S(n10), .Z(n1205) );
  MUX2_X1 U3049 ( .A(\REGISTERS[29][0] ), .B(n3039), .S(n10), .Z(n1204) );
  OAI21_X1 U3050 ( .B1(n3052), .B2(n3079), .A(n3042), .ZN(n3087) );
  NAND3_X1 U3051 ( .A1(ADD_WR[0]), .A2(n3080), .A3(ADD_WR[2]), .ZN(n3052) );
  INV_X1 U3052 ( .A(ADD_WR[1]), .ZN(n3080) );
  MUX2_X1 U3053 ( .A(\REGISTERS[30][31] ), .B(n3007), .S(n12), .Z(n1203) );
  MUX2_X1 U3054 ( .A(\REGISTERS[30][30] ), .B(n3009), .S(n12), .Z(n1202) );
  MUX2_X1 U3055 ( .A(\REGISTERS[30][29] ), .B(n3010), .S(n12), .Z(n1201) );
  MUX2_X1 U3056 ( .A(\REGISTERS[30][28] ), .B(n3011), .S(n12), .Z(n1200) );
  MUX2_X1 U3057 ( .A(\REGISTERS[30][27] ), .B(n3012), .S(n12), .Z(n1199) );
  MUX2_X1 U3058 ( .A(\REGISTERS[30][26] ), .B(n3013), .S(n12), .Z(n1198) );
  MUX2_X1 U3059 ( .A(\REGISTERS[30][25] ), .B(n3014), .S(n12), .Z(n1197) );
  MUX2_X1 U3060 ( .A(\REGISTERS[30][24] ), .B(n3015), .S(n12), .Z(n1196) );
  MUX2_X1 U3061 ( .A(\REGISTERS[30][23] ), .B(n3016), .S(n12), .Z(n1195) );
  MUX2_X1 U3062 ( .A(\REGISTERS[30][22] ), .B(n3017), .S(n12), .Z(n1194) );
  MUX2_X1 U3063 ( .A(\REGISTERS[30][21] ), .B(n3018), .S(n12), .Z(n1193) );
  MUX2_X1 U3064 ( .A(\REGISTERS[30][20] ), .B(n3019), .S(n12), .Z(n1192) );
  MUX2_X1 U3065 ( .A(\REGISTERS[30][19] ), .B(n3020), .S(n12), .Z(n1191) );
  MUX2_X1 U3066 ( .A(\REGISTERS[30][18] ), .B(n3021), .S(n12), .Z(n1190) );
  MUX2_X1 U3067 ( .A(\REGISTERS[30][17] ), .B(n3022), .S(n12), .Z(n1189) );
  MUX2_X1 U3068 ( .A(\REGISTERS[30][16] ), .B(n3023), .S(n12), .Z(n1188) );
  MUX2_X1 U3069 ( .A(\REGISTERS[30][15] ), .B(n3024), .S(n12), .Z(n1187) );
  MUX2_X1 U3070 ( .A(\REGISTERS[30][14] ), .B(n3025), .S(n12), .Z(n1186) );
  MUX2_X1 U3071 ( .A(\REGISTERS[30][13] ), .B(n3026), .S(n12), .Z(n1185) );
  MUX2_X1 U3072 ( .A(\REGISTERS[30][12] ), .B(n3027), .S(n12), .Z(n1184) );
  MUX2_X1 U3073 ( .A(\REGISTERS[30][11] ), .B(n3028), .S(n12), .Z(n1183) );
  MUX2_X1 U3074 ( .A(\REGISTERS[30][10] ), .B(n3029), .S(n12), .Z(n1182) );
  MUX2_X1 U3075 ( .A(\REGISTERS[30][9] ), .B(n3030), .S(n12), .Z(n1181) );
  MUX2_X1 U3076 ( .A(\REGISTERS[30][8] ), .B(n3031), .S(n12), .Z(n1180) );
  MUX2_X1 U3077 ( .A(\REGISTERS[30][7] ), .B(n3032), .S(n12), .Z(n1179) );
  MUX2_X1 U3078 ( .A(\REGISTERS[30][6] ), .B(n3033), .S(n12), .Z(n1178) );
  MUX2_X1 U3079 ( .A(\REGISTERS[30][5] ), .B(n3034), .S(n12), .Z(n1177) );
  MUX2_X1 U3080 ( .A(\REGISTERS[30][4] ), .B(n3035), .S(n12), .Z(n1176) );
  MUX2_X1 U3081 ( .A(\REGISTERS[30][3] ), .B(n3036), .S(n12), .Z(n1175) );
  MUX2_X1 U3082 ( .A(\REGISTERS[30][2] ), .B(n3037), .S(n12), .Z(n1174) );
  MUX2_X1 U3083 ( .A(\REGISTERS[30][1] ), .B(n3038), .S(n12), .Z(n1173) );
  MUX2_X1 U3084 ( .A(\REGISTERS[30][0] ), .B(n3039), .S(n12), .Z(n1172) );
  OAI21_X1 U3085 ( .B1(n3054), .B2(n3079), .A(n3042), .ZN(n3088) );
  NAND3_X1 U3086 ( .A1(ADD_WR[1]), .A2(n3082), .A3(ADD_WR[2]), .ZN(n3054) );
  INV_X1 U3087 ( .A(ADD_WR[0]), .ZN(n3082) );
  MUX2_X1 U3088 ( .A(\REGISTERS[31][31] ), .B(n3007), .S(n14), .Z(n1171) );
  AND2_X1 U3089 ( .A1(DATAIN[31]), .A2(n3042), .ZN(n3007) );
  MUX2_X1 U3090 ( .A(\REGISTERS[31][30] ), .B(n3009), .S(n14), .Z(n1170) );
  AND2_X1 U3091 ( .A1(DATAIN[30]), .A2(n3042), .ZN(n3009) );
  MUX2_X1 U3092 ( .A(\REGISTERS[31][29] ), .B(n3010), .S(n14), .Z(n1169) );
  AND2_X1 U3093 ( .A1(DATAIN[29]), .A2(n3042), .ZN(n3010) );
  MUX2_X1 U3094 ( .A(\REGISTERS[31][28] ), .B(n3011), .S(n14), .Z(n1168) );
  AND2_X1 U3095 ( .A1(DATAIN[28]), .A2(n3042), .ZN(n3011) );
  MUX2_X1 U3096 ( .A(\REGISTERS[31][27] ), .B(n3012), .S(n14), .Z(n1167) );
  AND2_X1 U3097 ( .A1(DATAIN[27]), .A2(n3042), .ZN(n3012) );
  MUX2_X1 U3098 ( .A(\REGISTERS[31][26] ), .B(n3013), .S(n14), .Z(n1166) );
  AND2_X1 U3099 ( .A1(DATAIN[26]), .A2(n3042), .ZN(n3013) );
  MUX2_X1 U3100 ( .A(\REGISTERS[31][25] ), .B(n3014), .S(n14), .Z(n1165) );
  AND2_X1 U3101 ( .A1(DATAIN[25]), .A2(n3042), .ZN(n3014) );
  MUX2_X1 U3102 ( .A(\REGISTERS[31][24] ), .B(n3015), .S(n14), .Z(n1164) );
  AND2_X1 U3103 ( .A1(DATAIN[24]), .A2(n3042), .ZN(n3015) );
  MUX2_X1 U3104 ( .A(\REGISTERS[31][23] ), .B(n3016), .S(n14), .Z(n1163) );
  AND2_X1 U3105 ( .A1(DATAIN[23]), .A2(n3042), .ZN(n3016) );
  MUX2_X1 U3106 ( .A(\REGISTERS[31][22] ), .B(n3017), .S(n14), .Z(n1162) );
  AND2_X1 U3107 ( .A1(DATAIN[22]), .A2(n3042), .ZN(n3017) );
  MUX2_X1 U3108 ( .A(\REGISTERS[31][21] ), .B(n3018), .S(n14), .Z(n1161) );
  AND2_X1 U3109 ( .A1(DATAIN[21]), .A2(n3042), .ZN(n3018) );
  MUX2_X1 U3110 ( .A(\REGISTERS[31][20] ), .B(n3019), .S(n14), .Z(n1160) );
  AND2_X1 U3111 ( .A1(DATAIN[20]), .A2(n3042), .ZN(n3019) );
  MUX2_X1 U3112 ( .A(\REGISTERS[31][19] ), .B(n3020), .S(n14), .Z(n1159) );
  AND2_X1 U3113 ( .A1(DATAIN[19]), .A2(n3042), .ZN(n3020) );
  MUX2_X1 U3114 ( .A(\REGISTERS[31][18] ), .B(n3021), .S(n14), .Z(n1158) );
  AND2_X1 U3115 ( .A1(DATAIN[18]), .A2(n3042), .ZN(n3021) );
  MUX2_X1 U3116 ( .A(\REGISTERS[31][17] ), .B(n3022), .S(n14), .Z(n1157) );
  AND2_X1 U3117 ( .A1(DATAIN[17]), .A2(n3042), .ZN(n3022) );
  MUX2_X1 U3118 ( .A(\REGISTERS[31][16] ), .B(n3023), .S(n14), .Z(n1156) );
  AND2_X1 U3119 ( .A1(DATAIN[16]), .A2(n3042), .ZN(n3023) );
  MUX2_X1 U3120 ( .A(\REGISTERS[31][15] ), .B(n3024), .S(n14), .Z(n1155) );
  AND2_X1 U3121 ( .A1(DATAIN[15]), .A2(n3042), .ZN(n3024) );
  MUX2_X1 U3122 ( .A(\REGISTERS[31][14] ), .B(n3025), .S(n14), .Z(n1154) );
  AND2_X1 U3123 ( .A1(DATAIN[14]), .A2(n3042), .ZN(n3025) );
  MUX2_X1 U3124 ( .A(\REGISTERS[31][13] ), .B(n3026), .S(n14), .Z(n1153) );
  AND2_X1 U3125 ( .A1(DATAIN[13]), .A2(n3042), .ZN(n3026) );
  MUX2_X1 U3126 ( .A(\REGISTERS[31][12] ), .B(n3027), .S(n14), .Z(n1152) );
  AND2_X1 U3127 ( .A1(DATAIN[12]), .A2(n3042), .ZN(n3027) );
  MUX2_X1 U3128 ( .A(\REGISTERS[31][11] ), .B(n3028), .S(n14), .Z(n1151) );
  AND2_X1 U3129 ( .A1(DATAIN[11]), .A2(n3042), .ZN(n3028) );
  MUX2_X1 U3130 ( .A(\REGISTERS[31][10] ), .B(n3029), .S(n14), .Z(n1150) );
  AND2_X1 U3131 ( .A1(DATAIN[10]), .A2(n3042), .ZN(n3029) );
  MUX2_X1 U3132 ( .A(\REGISTERS[31][9] ), .B(n3030), .S(n14), .Z(n1149) );
  AND2_X1 U3133 ( .A1(DATAIN[9]), .A2(n3042), .ZN(n3030) );
  MUX2_X1 U3134 ( .A(\REGISTERS[31][8] ), .B(n3031), .S(n14), .Z(n1148) );
  AND2_X1 U3135 ( .A1(DATAIN[8]), .A2(n3042), .ZN(n3031) );
  MUX2_X1 U3136 ( .A(\REGISTERS[31][7] ), .B(n3032), .S(n14), .Z(n1147) );
  AND2_X1 U3137 ( .A1(DATAIN[7]), .A2(n3042), .ZN(n3032) );
  MUX2_X1 U3138 ( .A(\REGISTERS[31][6] ), .B(n3033), .S(n14), .Z(n1146) );
  AND2_X1 U3139 ( .A1(DATAIN[6]), .A2(n3042), .ZN(n3033) );
  MUX2_X1 U3140 ( .A(\REGISTERS[31][5] ), .B(n3034), .S(n14), .Z(n1145) );
  AND2_X1 U3141 ( .A1(DATAIN[5]), .A2(n3042), .ZN(n3034) );
  MUX2_X1 U3142 ( .A(\REGISTERS[31][4] ), .B(n3035), .S(n14), .Z(n1144) );
  AND2_X1 U3143 ( .A1(DATAIN[4]), .A2(n3042), .ZN(n3035) );
  MUX2_X1 U3144 ( .A(\REGISTERS[31][3] ), .B(n3036), .S(n14), .Z(n1143) );
  AND2_X1 U3145 ( .A1(DATAIN[3]), .A2(n3042), .ZN(n3036) );
  MUX2_X1 U3146 ( .A(\REGISTERS[31][2] ), .B(n3037), .S(n14), .Z(n1142) );
  AND2_X1 U3147 ( .A1(DATAIN[2]), .A2(n3042), .ZN(n3037) );
  MUX2_X1 U3148 ( .A(\REGISTERS[31][1] ), .B(n3038), .S(n14), .Z(n1141) );
  AND2_X1 U3149 ( .A1(DATAIN[1]), .A2(n3042), .ZN(n3038) );
  MUX2_X1 U3150 ( .A(\REGISTERS[31][0] ), .B(n3039), .S(n14), .Z(n1140) );
  OAI21_X1 U3151 ( .B1(n3056), .B2(n3079), .A(n3042), .ZN(n3089) );
  NAND3_X1 U3152 ( .A1(ADD_WR[3]), .A2(n3059), .A3(ADD_WR[4]), .ZN(n3079) );
  AND2_X1 U3153 ( .A1(WR), .A2(ENABLE), .ZN(n3059) );
  NAND3_X1 U3154 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n3056)
         );
  AND2_X1 U3155 ( .A1(DATAIN[0]), .A2(n3042), .ZN(n3039) );
  AND2_X1 U3156 ( .A1(RD2), .A2(ENABLE), .ZN(N445) );
  AND2_X1 U3157 ( .A1(RD1), .A2(ENABLE), .ZN(N444) );
endmodule


module ffd_0 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n3, n1, n2, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n3) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_132 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_131 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_130 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_129 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_128 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_127 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_126 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_125 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_124 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_123 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_122 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_121 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_120 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_119 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_118 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_117 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_116 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_115 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_114 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_113 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_112 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_111 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_110 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_109 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_108 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_107 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_106 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_105 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_104 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_103 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_102 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_0 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_0 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_132 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_131 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_130 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_129 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_128 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_127 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_126 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_125 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_124 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_123 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_122 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_121 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_120 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_119 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_118 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_117 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_116 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_115 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_114 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_113 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_112 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_111 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_110 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_109 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_108 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_107 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_106 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_105 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_104 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_103 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_102 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_101 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_100 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_99 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_98 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_97 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_96 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_95 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_94 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_93 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_92 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_91 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_90 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_89 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_88 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_87 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_86 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_85 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_84 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_83 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_82 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_81 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_80 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_79 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_78 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_77 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_76 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_75 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_74 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_73 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_72 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_71 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_70 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_3 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_101 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_100 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_99 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_98 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_97 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_96 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_95 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_94 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_93 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_92 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_91 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_90 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_89 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_88 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_87 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_86 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_85 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_84 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_83 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_82 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_81 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_80 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_79 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_78 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_77 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_76 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_75 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_74 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_73 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_72 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_71 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_70 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_69 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_68 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_67 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_66 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_65 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_64 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_63 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_62 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_61 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_60 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_59 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_58 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_57 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_56 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_55 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_54 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_53 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_52 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_51 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_50 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_49 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_48 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_47 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_46 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_45 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_44 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_43 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_42 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_41 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_40 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_39 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_38 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_2 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_69 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_68 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_67 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_66 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_65 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_64 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_63 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_62 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_61 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_60 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_59 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_58 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_57 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_56 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_55 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_54 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_53 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_52 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_51 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_50 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_49 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_48 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_47 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_46 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_45 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_44 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_43 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_42 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_41 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_40 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_39 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_38 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_37 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_36 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_35 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_34 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_33 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_32 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_31 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_30 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_29 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_28 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_27 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_26 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_25 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_24 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_23 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_22 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_21 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_20 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_19 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_18 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_17 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_16 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_15 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_14 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_13 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_12 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_11 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_10 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_9 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_8 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_7 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_6 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_1 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_37 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_36 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_35 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_34 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_33 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_32 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_31 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_30 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_29 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_28 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_27 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_26 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_25 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_24 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_23 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_22 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_21 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_20 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_19 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_18 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_17 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_16 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_15 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_14 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_13 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_12 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_11 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_10 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_9 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_8 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_7 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_6 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_5 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_4 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_3 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_2 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_1 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N5 ( regIn, Clk, Reset, Enable, regOut );
  input [4:0] regIn;
  output [4:0] regOut;
  input Clk, Reset, Enable;


  ffd_5 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_4 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_3 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_2 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_1 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module MUX41_GENERIC_N32 ( SHIFTER_OUT, ADD_OUT, CMP_OUT, LOGICALS_OUT, SEL, Y
 );
  input [31:0] SHIFTER_OUT;
  input [31:0] ADD_OUT;
  input [31:0] CMP_OUT;
  input [31:0] LOGICALS_OUT;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  OR2_X1 U1 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n1) );
  OR2_X1 U2 ( .A1(n71), .A2(SEL[1]), .ZN(n2) );
  INV_X2 U3 ( .A(n2), .ZN(n3) );
  INV_X2 U4 ( .A(n1), .ZN(n4) );
  AND2_X2 U5 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n8) );
  AND2_X2 U6 ( .A1(SEL[1]), .A2(n71), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n5), .A2(n6), .ZN(Y[9]) );
  AOI22_X1 U8 ( .A1(CMP_OUT[9]), .A2(n7), .B1(LOGICALS_OUT[9]), .B2(n8), .ZN(
        n6) );
  AOI22_X1 U9 ( .A1(SHIFTER_OUT[9]), .A2(n4), .B1(ADD_OUT[9]), .B2(n3), .ZN(n5) );
  NAND2_X1 U10 ( .A1(n9), .A2(n10), .ZN(Y[8]) );
  AOI22_X1 U11 ( .A1(CMP_OUT[8]), .A2(n7), .B1(LOGICALS_OUT[8]), .B2(n8), .ZN(
        n10) );
  AOI22_X1 U12 ( .A1(SHIFTER_OUT[8]), .A2(n4), .B1(ADD_OUT[8]), .B2(n3), .ZN(
        n9) );
  NAND2_X1 U13 ( .A1(n11), .A2(n12), .ZN(Y[7]) );
  AOI22_X1 U14 ( .A1(CMP_OUT[7]), .A2(n7), .B1(LOGICALS_OUT[7]), .B2(n8), .ZN(
        n12) );
  AOI22_X1 U15 ( .A1(SHIFTER_OUT[7]), .A2(n4), .B1(ADD_OUT[7]), .B2(n3), .ZN(
        n11) );
  NAND2_X1 U16 ( .A1(n13), .A2(n14), .ZN(Y[6]) );
  AOI22_X1 U17 ( .A1(CMP_OUT[6]), .A2(n7), .B1(LOGICALS_OUT[6]), .B2(n8), .ZN(
        n14) );
  AOI22_X1 U18 ( .A1(SHIFTER_OUT[6]), .A2(n4), .B1(ADD_OUT[6]), .B2(n3), .ZN(
        n13) );
  NAND2_X1 U19 ( .A1(n15), .A2(n16), .ZN(Y[5]) );
  AOI22_X1 U20 ( .A1(CMP_OUT[5]), .A2(n7), .B1(LOGICALS_OUT[5]), .B2(n8), .ZN(
        n16) );
  AOI22_X1 U21 ( .A1(SHIFTER_OUT[5]), .A2(n4), .B1(ADD_OUT[5]), .B2(n3), .ZN(
        n15) );
  NAND2_X1 U22 ( .A1(n17), .A2(n18), .ZN(Y[4]) );
  AOI22_X1 U23 ( .A1(CMP_OUT[4]), .A2(n7), .B1(LOGICALS_OUT[4]), .B2(n8), .ZN(
        n18) );
  AOI22_X1 U24 ( .A1(SHIFTER_OUT[4]), .A2(n4), .B1(ADD_OUT[4]), .B2(n3), .ZN(
        n17) );
  NAND2_X1 U25 ( .A1(n19), .A2(n20), .ZN(Y[3]) );
  AOI22_X1 U26 ( .A1(CMP_OUT[3]), .A2(n7), .B1(LOGICALS_OUT[3]), .B2(n8), .ZN(
        n20) );
  AOI22_X1 U27 ( .A1(SHIFTER_OUT[3]), .A2(n4), .B1(ADD_OUT[3]), .B2(n3), .ZN(
        n19) );
  NAND2_X1 U28 ( .A1(n21), .A2(n22), .ZN(Y[31]) );
  AOI22_X1 U29 ( .A1(CMP_OUT[31]), .A2(n7), .B1(LOGICALS_OUT[31]), .B2(n8), 
        .ZN(n22) );
  AOI22_X1 U30 ( .A1(SHIFTER_OUT[31]), .A2(n4), .B1(ADD_OUT[31]), .B2(n3), 
        .ZN(n21) );
  NAND2_X1 U31 ( .A1(n23), .A2(n24), .ZN(Y[30]) );
  AOI22_X1 U32 ( .A1(CMP_OUT[30]), .A2(n7), .B1(LOGICALS_OUT[30]), .B2(n8), 
        .ZN(n24) );
  AOI22_X1 U33 ( .A1(SHIFTER_OUT[30]), .A2(n4), .B1(ADD_OUT[30]), .B2(n3), 
        .ZN(n23) );
  NAND2_X1 U34 ( .A1(n25), .A2(n26), .ZN(Y[2]) );
  AOI22_X1 U35 ( .A1(CMP_OUT[2]), .A2(n7), .B1(LOGICALS_OUT[2]), .B2(n8), .ZN(
        n26) );
  AOI22_X1 U36 ( .A1(SHIFTER_OUT[2]), .A2(n4), .B1(ADD_OUT[2]), .B2(n3), .ZN(
        n25) );
  NAND2_X1 U37 ( .A1(n27), .A2(n28), .ZN(Y[29]) );
  AOI22_X1 U38 ( .A1(CMP_OUT[29]), .A2(n7), .B1(LOGICALS_OUT[29]), .B2(n8), 
        .ZN(n28) );
  AOI22_X1 U39 ( .A1(SHIFTER_OUT[29]), .A2(n4), .B1(ADD_OUT[29]), .B2(n3), 
        .ZN(n27) );
  NAND2_X1 U40 ( .A1(n29), .A2(n30), .ZN(Y[28]) );
  AOI22_X1 U41 ( .A1(CMP_OUT[28]), .A2(n7), .B1(LOGICALS_OUT[28]), .B2(n8), 
        .ZN(n30) );
  AOI22_X1 U42 ( .A1(SHIFTER_OUT[28]), .A2(n4), .B1(ADD_OUT[28]), .B2(n3), 
        .ZN(n29) );
  NAND2_X1 U43 ( .A1(n31), .A2(n32), .ZN(Y[27]) );
  AOI22_X1 U44 ( .A1(CMP_OUT[27]), .A2(n7), .B1(LOGICALS_OUT[27]), .B2(n8), 
        .ZN(n32) );
  AOI22_X1 U45 ( .A1(SHIFTER_OUT[27]), .A2(n4), .B1(ADD_OUT[27]), .B2(n3), 
        .ZN(n31) );
  NAND2_X1 U46 ( .A1(n33), .A2(n34), .ZN(Y[26]) );
  AOI22_X1 U47 ( .A1(CMP_OUT[26]), .A2(n7), .B1(LOGICALS_OUT[26]), .B2(n8), 
        .ZN(n34) );
  AOI22_X1 U48 ( .A1(SHIFTER_OUT[26]), .A2(n4), .B1(ADD_OUT[26]), .B2(n3), 
        .ZN(n33) );
  NAND2_X1 U49 ( .A1(n35), .A2(n36), .ZN(Y[25]) );
  AOI22_X1 U50 ( .A1(CMP_OUT[25]), .A2(n7), .B1(LOGICALS_OUT[25]), .B2(n8), 
        .ZN(n36) );
  AOI22_X1 U51 ( .A1(SHIFTER_OUT[25]), .A2(n4), .B1(ADD_OUT[25]), .B2(n3), 
        .ZN(n35) );
  NAND2_X1 U52 ( .A1(n37), .A2(n38), .ZN(Y[24]) );
  AOI22_X1 U53 ( .A1(CMP_OUT[24]), .A2(n7), .B1(LOGICALS_OUT[24]), .B2(n8), 
        .ZN(n38) );
  AOI22_X1 U54 ( .A1(SHIFTER_OUT[24]), .A2(n4), .B1(ADD_OUT[24]), .B2(n3), 
        .ZN(n37) );
  NAND2_X1 U55 ( .A1(n39), .A2(n40), .ZN(Y[23]) );
  AOI22_X1 U56 ( .A1(CMP_OUT[23]), .A2(n7), .B1(LOGICALS_OUT[23]), .B2(n8), 
        .ZN(n40) );
  AOI22_X1 U57 ( .A1(SHIFTER_OUT[23]), .A2(n4), .B1(ADD_OUT[23]), .B2(n3), 
        .ZN(n39) );
  NAND2_X1 U58 ( .A1(n41), .A2(n42), .ZN(Y[22]) );
  AOI22_X1 U59 ( .A1(CMP_OUT[22]), .A2(n7), .B1(LOGICALS_OUT[22]), .B2(n8), 
        .ZN(n42) );
  AOI22_X1 U60 ( .A1(SHIFTER_OUT[22]), .A2(n4), .B1(ADD_OUT[22]), .B2(n3), 
        .ZN(n41) );
  NAND2_X1 U61 ( .A1(n43), .A2(n44), .ZN(Y[21]) );
  AOI22_X1 U62 ( .A1(CMP_OUT[21]), .A2(n7), .B1(LOGICALS_OUT[21]), .B2(n8), 
        .ZN(n44) );
  AOI22_X1 U63 ( .A1(SHIFTER_OUT[21]), .A2(n4), .B1(ADD_OUT[21]), .B2(n3), 
        .ZN(n43) );
  NAND2_X1 U64 ( .A1(n45), .A2(n46), .ZN(Y[20]) );
  AOI22_X1 U65 ( .A1(CMP_OUT[20]), .A2(n7), .B1(LOGICALS_OUT[20]), .B2(n8), 
        .ZN(n46) );
  AOI22_X1 U66 ( .A1(SHIFTER_OUT[20]), .A2(n4), .B1(ADD_OUT[20]), .B2(n3), 
        .ZN(n45) );
  NAND2_X1 U67 ( .A1(n47), .A2(n48), .ZN(Y[1]) );
  AOI22_X1 U68 ( .A1(CMP_OUT[1]), .A2(n7), .B1(LOGICALS_OUT[1]), .B2(n8), .ZN(
        n48) );
  AOI22_X1 U69 ( .A1(SHIFTER_OUT[1]), .A2(n4), .B1(ADD_OUT[1]), .B2(n3), .ZN(
        n47) );
  NAND2_X1 U70 ( .A1(n49), .A2(n50), .ZN(Y[19]) );
  AOI22_X1 U71 ( .A1(CMP_OUT[19]), .A2(n7), .B1(LOGICALS_OUT[19]), .B2(n8), 
        .ZN(n50) );
  AOI22_X1 U72 ( .A1(SHIFTER_OUT[19]), .A2(n4), .B1(ADD_OUT[19]), .B2(n3), 
        .ZN(n49) );
  NAND2_X1 U73 ( .A1(n51), .A2(n52), .ZN(Y[18]) );
  AOI22_X1 U74 ( .A1(CMP_OUT[18]), .A2(n7), .B1(LOGICALS_OUT[18]), .B2(n8), 
        .ZN(n52) );
  AOI22_X1 U75 ( .A1(SHIFTER_OUT[18]), .A2(n4), .B1(ADD_OUT[18]), .B2(n3), 
        .ZN(n51) );
  NAND2_X1 U76 ( .A1(n53), .A2(n54), .ZN(Y[17]) );
  AOI22_X1 U77 ( .A1(CMP_OUT[17]), .A2(n7), .B1(LOGICALS_OUT[17]), .B2(n8), 
        .ZN(n54) );
  AOI22_X1 U78 ( .A1(SHIFTER_OUT[17]), .A2(n4), .B1(ADD_OUT[17]), .B2(n3), 
        .ZN(n53) );
  NAND2_X1 U79 ( .A1(n55), .A2(n56), .ZN(Y[16]) );
  AOI22_X1 U80 ( .A1(CMP_OUT[16]), .A2(n7), .B1(LOGICALS_OUT[16]), .B2(n8), 
        .ZN(n56) );
  AOI22_X1 U81 ( .A1(SHIFTER_OUT[16]), .A2(n4), .B1(ADD_OUT[16]), .B2(n3), 
        .ZN(n55) );
  NAND2_X1 U82 ( .A1(n57), .A2(n58), .ZN(Y[15]) );
  AOI22_X1 U83 ( .A1(CMP_OUT[15]), .A2(n7), .B1(LOGICALS_OUT[15]), .B2(n8), 
        .ZN(n58) );
  AOI22_X1 U84 ( .A1(SHIFTER_OUT[15]), .A2(n4), .B1(ADD_OUT[15]), .B2(n3), 
        .ZN(n57) );
  NAND2_X1 U85 ( .A1(n59), .A2(n60), .ZN(Y[14]) );
  AOI22_X1 U86 ( .A1(CMP_OUT[14]), .A2(n7), .B1(LOGICALS_OUT[14]), .B2(n8), 
        .ZN(n60) );
  AOI22_X1 U87 ( .A1(SHIFTER_OUT[14]), .A2(n4), .B1(ADD_OUT[14]), .B2(n3), 
        .ZN(n59) );
  NAND2_X1 U88 ( .A1(n61), .A2(n62), .ZN(Y[13]) );
  AOI22_X1 U89 ( .A1(CMP_OUT[13]), .A2(n7), .B1(LOGICALS_OUT[13]), .B2(n8), 
        .ZN(n62) );
  AOI22_X1 U90 ( .A1(SHIFTER_OUT[13]), .A2(n4), .B1(ADD_OUT[13]), .B2(n3), 
        .ZN(n61) );
  NAND2_X1 U91 ( .A1(n63), .A2(n64), .ZN(Y[12]) );
  AOI22_X1 U92 ( .A1(CMP_OUT[12]), .A2(n7), .B1(LOGICALS_OUT[12]), .B2(n8), 
        .ZN(n64) );
  AOI22_X1 U93 ( .A1(SHIFTER_OUT[12]), .A2(n4), .B1(ADD_OUT[12]), .B2(n3), 
        .ZN(n63) );
  NAND2_X1 U94 ( .A1(n65), .A2(n66), .ZN(Y[11]) );
  AOI22_X1 U95 ( .A1(CMP_OUT[11]), .A2(n7), .B1(LOGICALS_OUT[11]), .B2(n8), 
        .ZN(n66) );
  AOI22_X1 U96 ( .A1(SHIFTER_OUT[11]), .A2(n4), .B1(ADD_OUT[11]), .B2(n3), 
        .ZN(n65) );
  NAND2_X1 U97 ( .A1(n67), .A2(n68), .ZN(Y[10]) );
  AOI22_X1 U98 ( .A1(CMP_OUT[10]), .A2(n7), .B1(LOGICALS_OUT[10]), .B2(n8), 
        .ZN(n68) );
  AOI22_X1 U99 ( .A1(SHIFTER_OUT[10]), .A2(n4), .B1(ADD_OUT[10]), .B2(n3), 
        .ZN(n67) );
  NAND2_X1 U100 ( .A1(n69), .A2(n70), .ZN(Y[0]) );
  AOI22_X1 U101 ( .A1(CMP_OUT[0]), .A2(n7), .B1(LOGICALS_OUT[0]), .B2(n8), 
        .ZN(n70) );
  AOI22_X1 U102 ( .A1(SHIFTER_OUT[0]), .A2(n4), .B1(ADD_OUT[0]), .B2(n3), .ZN(
        n69) );
  INV_X1 U103 ( .A(SEL[0]), .ZN(n71) );
endmodule


module IR_decoder_N32 ( IR_IN, RS1, RS2, RD, imm16, imm26 );
  input [31:0] IR_IN;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [15:0] imm16;
  output [25:0] imm26;
  wire   \IR_IN[25] , \IR_IN[24] , \IR_IN[23] , \IR_IN[22] , \IR_IN[21] ,
         \IR_IN[20] , \IR_IN[19] , \IR_IN[18] , \IR_IN[17] , \IR_IN[16] ,
         \IR_IN[15] , \IR_IN[14] , \IR_IN[13] , \IR_IN[12] , \IR_IN[11] ,
         \IR_IN[10] , \IR_IN[9] , \IR_IN[8] , \IR_IN[7] , \IR_IN[6] ,
         \IR_IN[5] , \IR_IN[4] , \IR_IN[3] , \IR_IN[2] , \IR_IN[1] ,
         \IR_IN[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9;
  assign imm26[25] = \IR_IN[25] ;
  assign RS1[4] = \IR_IN[25] ;
  assign \IR_IN[25]  = IR_IN[25];
  assign imm26[24] = \IR_IN[24] ;
  assign RS1[3] = \IR_IN[24] ;
  assign \IR_IN[24]  = IR_IN[24];
  assign imm26[23] = \IR_IN[23] ;
  assign RS1[2] = \IR_IN[23] ;
  assign \IR_IN[23]  = IR_IN[23];
  assign imm26[22] = \IR_IN[22] ;
  assign RS1[1] = \IR_IN[22] ;
  assign \IR_IN[22]  = IR_IN[22];
  assign imm26[21] = \IR_IN[21] ;
  assign RS1[0] = \IR_IN[21] ;
  assign \IR_IN[21]  = IR_IN[21];
  assign imm26[20] = \IR_IN[20] ;
  assign RS2[4] = \IR_IN[20] ;
  assign \IR_IN[20]  = IR_IN[20];
  assign imm26[19] = \IR_IN[19] ;
  assign RS2[3] = \IR_IN[19] ;
  assign \IR_IN[19]  = IR_IN[19];
  assign imm26[18] = \IR_IN[18] ;
  assign RS2[2] = \IR_IN[18] ;
  assign \IR_IN[18]  = IR_IN[18];
  assign imm26[17] = \IR_IN[17] ;
  assign RS2[1] = \IR_IN[17] ;
  assign \IR_IN[17]  = IR_IN[17];
  assign imm26[16] = \IR_IN[16] ;
  assign RS2[0] = \IR_IN[16] ;
  assign \IR_IN[16]  = IR_IN[16];
  assign imm26[15] = \IR_IN[15] ;
  assign imm16[15] = \IR_IN[15] ;
  assign \IR_IN[15]  = IR_IN[15];
  assign imm26[14] = \IR_IN[14] ;
  assign imm16[14] = \IR_IN[14] ;
  assign \IR_IN[14]  = IR_IN[14];
  assign imm26[13] = \IR_IN[13] ;
  assign imm16[13] = \IR_IN[13] ;
  assign \IR_IN[13]  = IR_IN[13];
  assign imm26[12] = \IR_IN[12] ;
  assign imm16[12] = \IR_IN[12] ;
  assign \IR_IN[12]  = IR_IN[12];
  assign imm26[11] = \IR_IN[11] ;
  assign imm16[11] = \IR_IN[11] ;
  assign \IR_IN[11]  = IR_IN[11];
  assign imm26[10] = \IR_IN[10] ;
  assign imm16[10] = \IR_IN[10] ;
  assign \IR_IN[10]  = IR_IN[10];
  assign imm26[9] = \IR_IN[9] ;
  assign imm16[9] = \IR_IN[9] ;
  assign \IR_IN[9]  = IR_IN[9];
  assign imm26[8] = \IR_IN[8] ;
  assign imm16[8] = \IR_IN[8] ;
  assign \IR_IN[8]  = IR_IN[8];
  assign imm26[7] = \IR_IN[7] ;
  assign imm16[7] = \IR_IN[7] ;
  assign \IR_IN[7]  = IR_IN[7];
  assign imm26[6] = \IR_IN[6] ;
  assign imm16[6] = \IR_IN[6] ;
  assign \IR_IN[6]  = IR_IN[6];
  assign imm26[5] = \IR_IN[5] ;
  assign imm16[5] = \IR_IN[5] ;
  assign \IR_IN[5]  = IR_IN[5];
  assign imm26[4] = \IR_IN[4] ;
  assign imm16[4] = \IR_IN[4] ;
  assign \IR_IN[4]  = IR_IN[4];
  assign imm26[3] = \IR_IN[3] ;
  assign imm16[3] = \IR_IN[3] ;
  assign \IR_IN[3]  = IR_IN[3];
  assign imm26[2] = \IR_IN[2] ;
  assign imm16[2] = \IR_IN[2] ;
  assign \IR_IN[2]  = IR_IN[2];
  assign imm26[1] = \IR_IN[1] ;
  assign imm16[1] = \IR_IN[1] ;
  assign \IR_IN[1]  = IR_IN[1];
  assign imm26[0] = \IR_IN[0] ;
  assign imm16[0] = \IR_IN[0] ;
  assign \IR_IN[0]  = IR_IN[0];

  NOR4_X2 U2 ( .A1(IR_IN[26]), .A2(n8), .A3(IR_IN[30]), .A4(IR_IN[27]), .ZN(n3) );
  OR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(RD[4]) );
  MUX2_X1 U4 ( .A(\IR_IN[20] ), .B(\IR_IN[15] ), .S(n3), .Z(n2) );
  OR2_X1 U5 ( .A1(n1), .A2(n4), .ZN(RD[3]) );
  MUX2_X1 U6 ( .A(\IR_IN[19] ), .B(\IR_IN[14] ), .S(n3), .Z(n4) );
  OR2_X1 U7 ( .A1(n1), .A2(n5), .ZN(RD[2]) );
  MUX2_X1 U8 ( .A(\IR_IN[18] ), .B(\IR_IN[13] ), .S(n3), .Z(n5) );
  OR2_X1 U9 ( .A1(n1), .A2(n6), .ZN(RD[1]) );
  MUX2_X1 U10 ( .A(\IR_IN[17] ), .B(\IR_IN[12] ), .S(n3), .Z(n6) );
  OR2_X1 U11 ( .A1(n1), .A2(n7), .ZN(RD[0]) );
  MUX2_X1 U12 ( .A(\IR_IN[16] ), .B(\IR_IN[11] ), .S(n3), .Z(n7) );
  INV_X1 U13 ( .A(n9), .ZN(n8) );
  AND3_X1 U14 ( .A1(IR_IN[26]), .A2(n9), .A3(IR_IN[27]), .ZN(n1) );
  NOR3_X1 U15 ( .A1(IR_IN[31]), .A2(IR_IN[29]), .A3(IR_IN[28]), .ZN(n9) );
endmodule


module DU ( IR_IN, NPC, WR_ADDR_RF, DATAIN, EN1, RF1, RF2, WF1, CLK, RST, 
        SEL_IMM, NPC1_OUT, regA_OUT, regB_OUT, IMM_OUT, RD1_IN, RD1_OUT );
  input [31:0] IR_IN;
  input [31:0] NPC;
  input [4:0] WR_ADDR_RF;
  input [31:0] DATAIN;
  input [1:0] SEL_IMM;
  output [31:0] NPC1_OUT;
  output [31:0] regA_OUT;
  output [31:0] regB_OUT;
  output [31:0] IMM_OUT;
  output [4:0] RD1_IN;
  output [4:0] RD1_OUT;
  input EN1, RF1, RF2, WF1, CLK, RST;
  wire   imm1632_31, imm2632_31;
  wire   [14:0] imm1632;
  wire   [24:0] imm2632;
  wire   [4:0] RS1s;
  wire   [4:0] RS2s;
  wire   [31:0] registerA;
  wire   [31:0] registerB;
  wire   [31:0] immediate32;

  register_file_WORD_SIZE32_ADDR_SIZE5 RegisterFile ( .CLK(CLK), .RESET(RST), 
        .ENABLE(EN1), .RD1(RF1), .RD2(RF2), .WR(WF1), .ADD_WR(WR_ADDR_RF), 
        .ADD_RD1(RS1s), .ADD_RD2(RS2s), .DATAIN(DATAIN), .OUT1(registerA), 
        .OUT2(registerB) );
  regN_N32_0 NPC1reg ( .regIn(NPC), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(NPC1_OUT) );
  regN_N32_3 Areg ( .regIn(registerA), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(regA_OUT) );
  regN_N32_2 Breg ( .regIn(registerB), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(regB_OUT) );
  regN_N32_1 IMMreg ( .regIn(immediate32), .Clk(CLK), .Reset(RST), .Enable(EN1), .regOut(IMM_OUT) );
  regN_N5 RD1reg ( .regIn(RD1_IN), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(RD1_OUT) );
  MUX41_GENERIC_N32 MUXimm ( .SHIFTER_OUT({imm1632_31, imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632}), .ADD_OUT({imm2632_31, imm2632_31, 
        imm2632_31, imm2632_31, imm2632_31, imm2632_31, imm2632_31, imm2632}), 
        .CMP_OUT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, imm1632_31, imm1632}), 
        .LOGICALS_OUT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, imm2632_31, imm2632}), .SEL(SEL_IMM), .Y(immediate32) );
  IR_decoder_N32 DEC ( .IR_IN(IR_IN), .RS1(RS1s), .RS2(RS2s), .RD(RD1_IN), 
        .imm16({imm1632_31, imm1632}), .imm26({imm2632_31, imm2632}) );
endmodule

