
module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_2 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_3 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_4 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_5 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_7 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_8 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_9 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_10 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_11 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_12 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_13 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_14 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_15 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_16 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_17 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_18 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_19 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_20 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_21 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_22 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_23 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_24 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_25 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_26 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_27 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_28 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_29 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_30 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_31 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module register_file_WORD_SIZE32_ADDR_SIZE5 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N444,
         n1025, n1026, n1027, n1028, n1030, n1031, n1032, n1033, n1035, n1036,
         n1037, n1038, n1040, n1041, n1042, n1043, n1045, n1046, n1047, n1048,
         n1050, n1051, n1052, n1053, n1055, n1056, n1057, n1058, n1060, n1061,
         n1062, n1063, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5707, n5709, n5711, n5713, n5715, n5717, n5719, n5721,
         n5723, n5725, n5727, n5729, n5731, n5733, n5735, n5737, n5739, n5741,
         n5743, n5745, n5747, n5749, n5751, n5753, n5755, n5757, n5759, n5761,
         n5763, n5765;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n5673), .CK(n5671), .QN(n5287) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n5674), .CK(n5671), .QN(n5288) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n5675), .CK(n5671), .QN(n5289) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n5676), .CK(n5671), .QN(n5290) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n5677), .CK(n5671), .QN(n5291) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n5678), .CK(n5671), .QN(n5292) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n5679), .CK(n5671), .QN(n5293) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n5680), .CK(n5671), .QN(n5294) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n5681), .CK(n5671), .QN(n5295) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n5682), .CK(n5671), .QN(n5296) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n5683), .CK(n5671), .QN(n5297) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n5684), .CK(n5671), .QN(n5298) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n5685), .CK(n5671), .QN(n5299) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n5686), .CK(n5671), .QN(n5300) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n5687), .CK(n5671), .QN(n5301) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n5688), .CK(n5671), .QN(n5302) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n5689), .CK(n5671), .QN(n5303) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n5690), .CK(n5671), .QN(n5304) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n5691), .CK(n5671), .QN(n5305) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n5692), .CK(n5671), .QN(n5306) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n5693), .CK(n5671), .QN(n5307) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n5694), .CK(n5671), .QN(n5308) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n5695), .CK(n5671), .QN(n5309) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n5696), .CK(n5671), .QN(n5310) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n5697), .CK(n5671), .QN(n5311) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n5698), .CK(n5671), .QN(n5312) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n5699), .CK(n5671), .QN(n5313) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n5700), .CK(n5671), .QN(n5314) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n5701), .CK(n5671), .QN(n5315) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n5702), .CK(n5671), .QN(n5316) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n5703), .CK(n5671), .QN(n5317) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n5704), .CK(n5671), .QN(n5318) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n5673), .CK(n5725), .QN(n5159) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n5674), .CK(n5725), .QN(n5163) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n5675), .CK(n5725), .QN(n5167) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n5676), .CK(n5725), .QN(n5171) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n5677), .CK(n5725), .QN(n5175) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n5678), .CK(n5725), .QN(n5179) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n5679), .CK(n5725), .QN(n5183) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n5680), .CK(n5725), .QN(n5187) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n5681), .CK(n5725), .QN(n5191) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n5682), .CK(n5725), .QN(n5195) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n5683), .CK(n5725), .QN(n5199) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n5684), .CK(n5725), .QN(n5203) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n5685), .CK(n5725), .QN(n5207) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n5686), .CK(n5725), .QN(n5211) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n5687), .CK(n5725), .QN(n5215) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n5688), .CK(n5725), .QN(n5219) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n5689), .CK(n5725), .QN(n5223) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n5690), .CK(n5725), .QN(n5227) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n5691), .CK(n5725), .QN(n5231) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n5692), .CK(n5725), .QN(n5235) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n5693), .CK(n5725), .QN(n5239) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n5694), .CK(n5725), .QN(n5243) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n5695), .CK(n5725), .QN(n5247) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n5696), .CK(n5725), .QN(n5251) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n5697), .CK(n5725), .QN(n5255) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n5698), .CK(n5725), .QN(n5259) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n5699), .CK(n5725), .QN(n5263) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n5700), .CK(n5725), .QN(n5267) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n5701), .CK(n5725), .QN(n5271) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n5702), .CK(n5725), .QN(n5275) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n5703), .CK(n5725), .QN(n5279) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n5704), .CK(n5725), .QN(n5283) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n5673), .CK(n5747), .QN(n5319) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n5674), .CK(n5747), .QN(n5320) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n5675), .CK(n5747), .QN(n5321) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n5676), .CK(n5747), .QN(n5322) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n5677), .CK(n5747), .QN(n5323) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n5678), .CK(n5747), .QN(n5324) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n5679), .CK(n5747), .QN(n5325) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n5680), .CK(n5747), .QN(n5326) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n5681), .CK(n5747), .QN(n5327) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n5682), .CK(n5747), .QN(n5328) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n5683), .CK(n5747), .QN(n5329) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n5684), .CK(n5747), .QN(n5330) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n5685), .CK(n5747), .QN(n5331) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n5686), .CK(n5747), .QN(n5332) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n5687), .CK(n5747), .QN(n5333) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n5688), .CK(n5747), .QN(n5334) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n5689), .CK(n5747), .QN(n5335) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n5690), .CK(n5747), .QN(n5336) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n5691), .CK(n5747), .QN(n5337) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n5692), .CK(n5747), .QN(n5338) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n5693), .CK(n5747), .QN(n5339) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n5694), .CK(n5747), .QN(n5340) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n5695), .CK(n5747), .QN(n5341) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n5696), .CK(n5747), .QN(n5342) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n5697), .CK(n5747), .QN(n5343) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n5698), .CK(n5747), .QN(n5344) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n5699), .CK(n5747), .QN(n5345) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n5700), .CK(n5747), .QN(n5346) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n5701), .CK(n5747), .QN(n5347) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n5702), .CK(n5747), .QN(n5348) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n5703), .CK(n5747), .QN(n5349) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n5704), .CK(n5747), .QN(n5350) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n5673), .CK(n5753), .QN(n5351) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n5674), .CK(n5753), .QN(n5352) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n5675), .CK(n5753), .QN(n5353) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n5676), .CK(n5753), .QN(n5354) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n5677), .CK(n5753), .QN(n5355) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n5678), .CK(n5753), .QN(n5356) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n5679), .CK(n5753), .QN(n5357) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n5680), .CK(n5753), .QN(n5358) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n5681), .CK(n5753), .QN(n5359) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n5682), .CK(n5753), .QN(n5360) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n5683), .CK(n5753), .QN(n5361) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n5684), .CK(n5753), .QN(n5362) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n5685), .CK(n5753), .QN(n5363) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n5686), .CK(n5753), .QN(n5364) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n5687), .CK(n5753), .QN(n5365) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n5688), .CK(n5753), .QN(n5366) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n5689), .CK(n5753), .QN(n5367) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n5690), .CK(n5753), .QN(n5368) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n5691), .CK(n5753), .QN(n5369) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n5692), .CK(n5753), .QN(n5370) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n5693), .CK(n5753), .QN(n5371) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n5694), .CK(n5753), .QN(n5372) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n5695), .CK(n5753), .QN(n5373) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n5696), .CK(n5753), .QN(n5374) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n5697), .CK(n5753), .QN(n5375) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n5698), .CK(n5753), .QN(n5376) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n5699), .CK(n5753), .QN(n5377) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n5700), .CK(n5753), .QN(n5378) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n5701), .CK(n5753), .QN(n5379) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n5702), .CK(n5753), .QN(n5380) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n5703), .CK(n5753), .QN(n5381) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n5704), .CK(n5753), .QN(n5382) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n5673), .CK(n5755), .QN(n5383) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n5674), .CK(n5755), .QN(n5384) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n5675), .CK(n5755), .QN(n5385) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n5676), .CK(n5755), .QN(n5386) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n5677), .CK(n5755), .QN(n5387) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n5678), .CK(n5755), .QN(n5388) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n5679), .CK(n5755), .QN(n5389) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n5680), .CK(n5755), .QN(n5390) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n5681), .CK(n5755), .QN(n5391) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n5682), .CK(n5755), .QN(n5392) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n5683), .CK(n5755), .QN(n5393) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n5684), .CK(n5755), .QN(n5394) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n5685), .CK(n5755), .QN(n5395) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n5686), .CK(n5755), .QN(n5396) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n5687), .CK(n5755), .QN(n5397) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n5688), .CK(n5755), .QN(n5398) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n5689), .CK(n5755), .QN(n5399) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n5690), .CK(n5755), .QN(n5400) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n5691), .CK(n5755), .QN(n5401) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n5692), .CK(n5755), .QN(n5402) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n5693), .CK(n5755), .QN(n5403) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n5694), .CK(n5755), .QN(n5404) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n5695), .CK(n5755), .QN(n5405) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n5696), .CK(n5755), .QN(n5406) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n5697), .CK(n5755), .QN(n5407) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n5698), .CK(n5755), .QN(n5408) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n5699), .CK(n5755), .QN(n5409) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n5700), .CK(n5755), .QN(n5410) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n5701), .CK(n5755), .QN(n5411) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n5702), .CK(n5755), .QN(n5412) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n5703), .CK(n5755), .QN(n5413) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n5704), .CK(n5755), .QN(n5414) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n5673), .CK(n5757), .QN(n5415) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n5674), .CK(n5757), .QN(n5416) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n5675), .CK(n5757), .QN(n5417) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n5676), .CK(n5757), .QN(n5418) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n5677), .CK(n5757), .QN(n5419) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n5678), .CK(n5757), .QN(n5420) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n5679), .CK(n5757), .QN(n5421) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n5680), .CK(n5757), .QN(n5422) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n5681), .CK(n5757), .QN(n5423) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n5682), .CK(n5757), .QN(n5424) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n5683), .CK(n5757), .QN(n5425) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n5684), .CK(n5757), .QN(n5426) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n5685), .CK(n5757), .QN(n5427) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n5686), .CK(n5757), .QN(n5428) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n5687), .CK(n5757), .QN(n5429) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n5688), .CK(n5757), .QN(n5430) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n5689), .CK(n5757), .QN(n5431) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n5690), .CK(n5757), .QN(n5432) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n5691), .CK(n5757), .QN(n5433) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n5692), .CK(n5757), .QN(n5434) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n5693), .CK(n5757), .QN(n5435) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n5694), .CK(n5757), .QN(n5436) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n5695), .CK(n5757), .QN(n5437) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n5696), .CK(n5757), .QN(n5438) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n5697), .CK(n5757), .QN(n5439) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n5698), .CK(n5757), .QN(n5440) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n5699), .CK(n5757), .QN(n5441) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n5700), .CK(n5757), .QN(n5442) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n5701), .CK(n5757), .QN(n5443) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n5702), .CK(n5757), .QN(n5444) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n5703), .CK(n5757), .QN(n5445) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n5704), .CK(n5757), .QN(n5446) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n5673), .CK(n5759), .QN(n5447) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n5674), .CK(n5759), .QN(n5448) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n5675), .CK(n5759), .QN(n5449) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n5676), .CK(n5759), .QN(n5450) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n5677), .CK(n5759), .QN(n5451) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n5678), .CK(n5759), .QN(n5452) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n5679), .CK(n5759), .QN(n5453) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n5680), .CK(n5759), .QN(n5454) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n5681), .CK(n5759), .QN(n5455) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n5682), .CK(n5759), .QN(n5456) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n5683), .CK(n5759), .QN(n5457) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n5684), .CK(n5759), .QN(n5458) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n5685), .CK(n5759), .QN(n5459) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n5686), .CK(n5759), .QN(n5460) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n5687), .CK(n5759), .QN(n5461) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n5688), .CK(n5759), .QN(n5462) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n5689), .CK(n5759), .QN(n5463) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n5690), .CK(n5759), .QN(n5464) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n5691), .CK(n5759), .QN(n5465) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n5692), .CK(n5759), .QN(n5466) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n5693), .CK(n5759), .QN(n5467) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n5694), .CK(n5759), .QN(n5468) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n5695), .CK(n5759), .QN(n5469) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n5696), .CK(n5759), .QN(n5470) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n5697), .CK(n5759), .QN(n5471) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n5698), .CK(n5759), .QN(n5472) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n5699), .CK(n5759), .QN(n5473) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n5700), .CK(n5759), .QN(n5474) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n5701), .CK(n5759), .QN(n5475) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n5702), .CK(n5759), .QN(n5476) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n5703), .CK(n5759), .QN(n5477) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n5704), .CK(n5759), .QN(n5478) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n5673), .CK(n5761), .Q(n3536) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n5674), .CK(n5761), .Q(n3535) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n5675), .CK(n5761), .Q(n3534) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n5676), .CK(n5761), .Q(n3533) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n5677), .CK(n5761), .Q(n3532) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n5678), .CK(n5761), .Q(n3531) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n5679), .CK(n5761), .Q(n3530) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n5680), .CK(n5761), .Q(n3529) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n5681), .CK(n5761), .Q(n3528) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n5682), .CK(n5761), .Q(n3527) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n5683), .CK(n5761), .Q(n3526) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n5684), .CK(n5761), .Q(n3525) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n5685), .CK(n5761), .Q(n3524) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n5686), .CK(n5761), .Q(n3523) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n5687), .CK(n5761), .Q(n3522) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n5688), .CK(n5761), .Q(n3521) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n5689), .CK(n5761), .Q(n3520) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n5690), .CK(n5761), .Q(n3519) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n5691), .CK(n5761), .Q(n3518) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n5692), .CK(n5761), .Q(n3517) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n5693), .CK(n5761), .Q(n3516) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n5694), .CK(n5761), .Q(n3515) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n5695), .CK(n5761), .Q(n3514) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n5696), .CK(n5761), .Q(n3513) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n5697), .CK(n5761), .Q(n3512) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n5698), .CK(n5761), .Q(n3511) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n5699), .CK(n5761), .Q(n3510) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n5700), .CK(n5761), .Q(n3509) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n5701), .CK(n5761), .Q(n3508) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n5702), .CK(n5761), .Q(n3507) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n5703), .CK(n5761), .Q(n3506) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n5704), .CK(n5761), .Q(n3505) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n5673), .CK(n5763), .Q(n3504) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n5674), .CK(n5763), .Q(n3503) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n5675), .CK(n5763), .Q(n3502) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n5676), .CK(n5763), .Q(n3501) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n5677), .CK(n5763), .Q(n3500) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n5678), .CK(n5763), .Q(n3499) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n5679), .CK(n5763), .Q(n3498) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n5680), .CK(n5763), .Q(n3497) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n5681), .CK(n5763), .Q(n3496) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n5682), .CK(n5763), .Q(n3495) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n5683), .CK(n5763), .Q(n3494) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n5684), .CK(n5763), .Q(n3493) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n5685), .CK(n5763), .Q(n3492) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n5686), .CK(n5763), .Q(n3491) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n5687), .CK(n5763), .Q(n3490) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n5688), .CK(n5763), .Q(n3489) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n5689), .CK(n5763), .Q(n3488) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n5690), .CK(n5763), .Q(n3487) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n5691), .CK(n5763), .Q(n3486) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n5692), .CK(n5763), .Q(n3485) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n5693), .CK(n5763), .Q(n3484) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n5694), .CK(n5763), .Q(n3483) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n5695), .CK(n5763), .Q(n3482) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n5696), .CK(n5763), .Q(n3481) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n5697), .CK(n5763), .Q(n3480) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n5698), .CK(n5763), .Q(n3479) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n5699), .CK(n5763), .Q(n3478) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n5700), .CK(n5763), .Q(n3477) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n5701), .CK(n5763), .Q(n3476) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n5702), .CK(n5763), .Q(n3475) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n5703), .CK(n5763), .Q(n3474) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n5704), .CK(n5763), .Q(n3473) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n5673), .CK(n5765), .QN(n5479) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n5674), .CK(n5765), .QN(n5480) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n5675), .CK(n5765), .QN(n5481) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n5676), .CK(n5765), .QN(n5482) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n5677), .CK(n5765), .QN(n5483) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n5678), .CK(n5765), .QN(n5484) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n5679), .CK(n5765), .QN(n5485) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n5680), .CK(n5765), .QN(n5486) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n5681), .CK(n5765), .QN(n5487) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n5682), .CK(n5765), .QN(n5488) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n5683), .CK(n5765), .QN(n5489) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n5684), .CK(n5765), .QN(n5490) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n5685), .CK(n5765), .QN(n5491) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n5686), .CK(n5765), .QN(n5492) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n5687), .CK(n5765), .QN(n5493) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n5688), .CK(n5765), .QN(n5494) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n5689), .CK(n5765), .QN(n5495) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n5690), .CK(n5765), .QN(n5496) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n5691), .CK(n5765), .QN(n5497) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n5692), .CK(n5765), .QN(n5498) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n5693), .CK(n5765), .QN(n5499) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n5694), .CK(n5765), .QN(n5500) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n5695), .CK(n5765), .QN(n5501) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n5696), .CK(n5765), .QN(n5502) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n5697), .CK(n5765), .QN(n5503) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n5698), .CK(n5765), .QN(n5504) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n5699), .CK(n5765), .QN(n5505) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n5700), .CK(n5765), .QN(n5506) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n5701), .CK(n5765), .QN(n5507) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n5702), .CK(n5765), .QN(n5508) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n5703), .CK(n5765), .QN(n5509) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n5704), .CK(n5765), .QN(n5510) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n5673), .CK(n5705), .Q(n3440) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n5674), .CK(n5705), .Q(n3439) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n5675), .CK(n5705), .Q(n3438) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n5676), .CK(n5705), .Q(n3437) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n5677), .CK(n5705), .Q(n3436) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n5678), .CK(n5705), .Q(n3435) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n5679), .CK(n5705), .Q(n3434) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n5680), .CK(n5705), .Q(n3433) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n5681), .CK(n5705), .Q(n3432) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n5682), .CK(n5705), .Q(n3431) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n5683), .CK(n5705), .Q(n3430) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n5684), .CK(n5705), .Q(n3429) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n5685), .CK(n5705), .Q(n3428) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n5686), .CK(n5705), .Q(n3427) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n5687), .CK(n5705), .Q(n3426) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n5688), .CK(n5705), .Q(n3425) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n5689), .CK(n5705), .Q(n3424) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n5690), .CK(n5705), .Q(n3423) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n5691), .CK(n5705), .Q(n3422) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n5692), .CK(n5705), .Q(n3421) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n5693), .CK(n5705), .Q(n3420) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n5694), .CK(n5705), .Q(n3419) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n5695), .CK(n5705), .Q(n3418) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n5696), .CK(n5705), .Q(n3417) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n5697), .CK(n5705), .Q(n3416) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n5698), .CK(n5705), .Q(n3415) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n5699), .CK(n5705), .Q(n3414) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n5700), .CK(n5705), .Q(n3413) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n5701), .CK(n5705), .Q(n3412) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n5702), .CK(n5705), .Q(n3411) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n5703), .CK(n5705), .Q(n3410) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n5704), .CK(n5705), .Q(n3409) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n5673), .CK(n5707), .Q(n3408) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n5674), .CK(n5707), .Q(n3407) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n5675), .CK(n5707), .Q(n3406) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n5676), .CK(n5707), .Q(n3405) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n5677), .CK(n5707), .Q(n3404) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n5678), .CK(n5707), .Q(n3403) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n5679), .CK(n5707), .Q(n3402) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n5680), .CK(n5707), .Q(n3401) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n5681), .CK(n5707), .Q(n3400) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n5682), .CK(n5707), .Q(n3399) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n5683), .CK(n5707), .Q(n3398) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n5684), .CK(n5707), .Q(n3397) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n5685), .CK(n5707), .Q(n3396) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n5686), .CK(n5707), .Q(n3395) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n5687), .CK(n5707), .Q(n3394) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n5688), .CK(n5707), .Q(n3393) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n5689), .CK(n5707), .Q(n3392) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n5690), .CK(n5707), .Q(n3391) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n5691), .CK(n5707), .Q(n3390) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n5692), .CK(n5707), .Q(n3389) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n5693), .CK(n5707), .Q(n3388) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n5694), .CK(n5707), .Q(n3387) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n5695), .CK(n5707), .Q(n3386) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n5696), .CK(n5707), .Q(n3385) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n5697), .CK(n5707), .Q(n3384) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n5698), .CK(n5707), .Q(n3383) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n5699), .CK(n5707), .Q(n3382) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n5700), .CK(n5707), .Q(n3381) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n5701), .CK(n5707), .Q(n3380) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n5702), .CK(n5707), .Q(n3379) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n5703), .CK(n5707), .Q(n3378) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n5704), .CK(n5707), .Q(n3377) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n5673), .CK(n5709), .QN(n5511) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n5674), .CK(n5709), .QN(n5512) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n5675), .CK(n5709), .QN(n5513) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n5676), .CK(n5709), .QN(n5514) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n5677), .CK(n5709), .QN(n5515) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n5678), .CK(n5709), .QN(n5516) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n5679), .CK(n5709), .QN(n5517) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n5680), .CK(n5709), .QN(n5518) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n5681), .CK(n5709), .QN(n5519) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n5682), .CK(n5709), .QN(n5520) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n5683), .CK(n5709), .QN(n5521) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n5684), .CK(n5709), .QN(n5522) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n5685), .CK(n5709), .QN(n5523) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n5686), .CK(n5709), .QN(n5524) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n5687), .CK(n5709), .QN(n5525) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n5688), .CK(n5709), .QN(n5526) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n5689), .CK(n5709), .QN(n5527) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n5690), .CK(n5709), .QN(n5528) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n5691), .CK(n5709), .QN(n5529) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n5692), .CK(n5709), .QN(n5530) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n5693), .CK(n5709), .QN(n5531) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n5694), .CK(n5709), .QN(n5532) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n5695), .CK(n5709), .QN(n5533) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n5696), .CK(n5709), .QN(n5534) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n5697), .CK(n5709), .QN(n5535) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n5698), .CK(n5709), .QN(n5536) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n5699), .CK(n5709), .QN(n5537) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n5700), .CK(n5709), .QN(n5538) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n5701), .CK(n5709), .QN(n5539) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n5702), .CK(n5709), .QN(n5540) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n5703), .CK(n5709), .QN(n5541) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n5704), .CK(n5709), .QN(n5542) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n5673), .CK(n5711), .Q(n3344) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n5674), .CK(n5711), .Q(n3343) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n5675), .CK(n5711), .Q(n3342) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n5676), .CK(n5711), .Q(n3341) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n5677), .CK(n5711), .Q(n3340) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n5678), .CK(n5711), .Q(n3339) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n5679), .CK(n5711), .Q(n3338) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n5680), .CK(n5711), .Q(n3337) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n5681), .CK(n5711), .Q(n3336) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n5682), .CK(n5711), .Q(n3335) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n5683), .CK(n5711), .Q(n3334) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n5684), .CK(n5711), .Q(n3333) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n5685), .CK(n5711), .Q(n3332) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n5686), .CK(n5711), .Q(n3331) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n5687), .CK(n5711), .Q(n3330) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n5688), .CK(n5711), .Q(n3329) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n5689), .CK(n5711), .Q(n3328) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n5690), .CK(n5711), .Q(n3327) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n5691), .CK(n5711), .Q(n3326) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n5692), .CK(n5711), .Q(n3325) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n5693), .CK(n5711), .Q(n3324) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n5694), .CK(n5711), .Q(n3323) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n5695), .CK(n5711), .Q(n3322) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n5696), .CK(n5711), .Q(n3321) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n5697), .CK(n5711), .Q(n3320) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n5698), .CK(n5711), .Q(n3319) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n5699), .CK(n5711), .Q(n3318) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n5700), .CK(n5711), .Q(n3317) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n5701), .CK(n5711), .Q(n3316) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n5702), .CK(n5711), .Q(n3315) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n5703), .CK(n5711), .Q(n3314) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n5704), .CK(n5711), .Q(n3313) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n5673), .CK(n5713), .QN(n5160) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n5674), .CK(n5713), .QN(n5164) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n5675), .CK(n5713), .QN(n5168) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n5676), .CK(n5713), .QN(n5172) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n5677), .CK(n5713), .QN(n5176) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n5678), .CK(n5713), .QN(n5180) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n5679), .CK(n5713), .QN(n5184) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n5680), .CK(n5713), .QN(n5188) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n5681), .CK(n5713), .QN(n5192) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n5682), .CK(n5713), .QN(n5196) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n5683), .CK(n5713), .QN(n5200) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n5684), .CK(n5713), .QN(n5204) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n5685), .CK(n5713), .QN(n5208) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n5686), .CK(n5713), .QN(n5212) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n5687), .CK(n5713), .QN(n5216) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n5688), .CK(n5713), .QN(n5220) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n5689), .CK(n5713), .QN(n5224) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n5690), .CK(n5713), .QN(n5228) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n5691), .CK(n5713), .QN(n5232) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n5692), .CK(n5713), .QN(n5236) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n5693), .CK(n5713), .QN(n5240) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n5694), .CK(n5713), .QN(n5244) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n5695), .CK(n5713), .QN(n5248) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n5696), .CK(n5713), .QN(n5252) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n5697), .CK(n5713), .QN(n5256) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n5698), .CK(n5713), .QN(n5260) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n5699), .CK(n5713), .QN(n5264) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n5700), .CK(n5713), .QN(n5268) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n5701), .CK(n5713), .QN(n5272) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n5702), .CK(n5713), .QN(n5276) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n5703), .CK(n5713), .QN(n5280) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n5704), .CK(n5713), .QN(n5284) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n5673), .CK(n5715), .Q(n3280) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n5674), .CK(n5715), .Q(n3279) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n5675), .CK(n5715), .Q(n3278) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n5676), .CK(n5715), .Q(n3277) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n5677), .CK(n5715), .Q(n3276) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n5678), .CK(n5715), .Q(n3275) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n5679), .CK(n5715), .Q(n3274) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n5680), .CK(n5715), .Q(n3273) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n5681), .CK(n5715), .Q(n3272) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n5682), .CK(n5715), .Q(n3271) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n5683), .CK(n5715), .Q(n3270) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n5684), .CK(n5715), .Q(n3269) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n5685), .CK(n5715), .Q(n3268) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n5686), .CK(n5715), .Q(n3267) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n5687), .CK(n5715), .Q(n3266) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n5688), .CK(n5715), .Q(n3265) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n5689), .CK(n5715), .Q(n3264) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n5690), .CK(n5715), .Q(n3263) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n5691), .CK(n5715), .Q(n3262) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n5692), .CK(n5715), .Q(n3261) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n5693), .CK(n5715), .Q(n3260) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n5694), .CK(n5715), .Q(n3259) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n5695), .CK(n5715), .Q(n3258) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n5696), .CK(n5715), .Q(n3257) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n5697), .CK(n5715), .Q(n3256) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n5698), .CK(n5715), .Q(n3255) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n5699), .CK(n5715), .Q(n3254) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n5700), .CK(n5715), .Q(n3253) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n5701), .CK(n5715), .Q(n3252) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n5702), .CK(n5715), .Q(n3251) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n5703), .CK(n5715), .Q(n3250) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n5704), .CK(n5715), .Q(n3249) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n5673), .CK(n5717), .QN(n5543) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n5674), .CK(n5717), .QN(n5544) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n5675), .CK(n5717), .QN(n5545) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n5676), .CK(n5717), .QN(n5546) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n5677), .CK(n5717), .QN(n5547) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n5678), .CK(n5717), .QN(n5548) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n5679), .CK(n5717), .QN(n5549) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n5680), .CK(n5717), .QN(n5550) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n5681), .CK(n5717), .QN(n5551) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n5682), .CK(n5717), .QN(n5552) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n5683), .CK(n5717), .QN(n5553) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n5684), .CK(n5717), .QN(n5554) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n5685), .CK(n5717), .QN(n5555) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n5686), .CK(n5717), .QN(n5556) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n5687), .CK(n5717), .QN(n5557) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n5688), .CK(n5717), .QN(n5558) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n5689), .CK(n5717), .QN(n5559) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n5690), .CK(n5717), .QN(n5560) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n5691), .CK(n5717), .QN(n5561) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n5692), .CK(n5717), .QN(n5562) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n5693), .CK(n5717), .QN(n5563) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n5694), .CK(n5717), .QN(n5564) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n5695), .CK(n5717), .QN(n5565) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n5696), .CK(n5717), .QN(n5566) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n5697), .CK(n5717), .QN(n5567) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n5698), .CK(n5717), .QN(n5568) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n5699), .CK(n5717), .QN(n5569) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n5700), .CK(n5717), .QN(n5570) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n5701), .CK(n5717), .QN(n5571) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n5702), .CK(n5717), .QN(n5572) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n5703), .CK(n5717), .QN(n5573) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n5704), .CK(n5717), .QN(n5574) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n5673), .CK(n5719), .Q(n3216) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n5674), .CK(n5719), .Q(n3215) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n5675), .CK(n5719), .Q(n3214) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n5676), .CK(n5719), .Q(n3213) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n5677), .CK(n5719), .Q(n3212) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n5678), .CK(n5719), .Q(n3211) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n5679), .CK(n5719), .Q(n3210) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n5680), .CK(n5719), .Q(n3209) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n5681), .CK(n5719), .Q(n3208) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n5682), .CK(n5719), .Q(n3207) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n5683), .CK(n5719), .Q(n3206) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n5684), .CK(n5719), .Q(n3205) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n5685), .CK(n5719), .Q(n3204) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n5686), .CK(n5719), .Q(n3203) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n5687), .CK(n5719), .Q(n3202) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n5688), .CK(n5719), .Q(n3201) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n5689), .CK(n5719), .Q(n3200) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n5690), .CK(n5719), .Q(n3199) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n5691), .CK(n5719), .Q(n3198) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n5692), .CK(n5719), .Q(n3197) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n5693), .CK(n5719), .Q(n3196) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n5694), .CK(n5719), .Q(n3195) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n5695), .CK(n5719), .Q(n3194) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n5696), .CK(n5719), .Q(n3193) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n5697), .CK(n5719), .Q(n3192) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n5698), .CK(n5719), .Q(n3191) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n5699), .CK(n5719), .Q(n3190) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n5700), .CK(n5719), .Q(n3189) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n5701), .CK(n5719), .Q(n3188) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n5702), .CK(n5719), .Q(n3187) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n5703), .CK(n5719), .Q(n3186) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n5704), .CK(n5719), .Q(n3185) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n5673), .CK(n5721), .Q(n3184) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n5674), .CK(n5721), .Q(n3183) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n5675), .CK(n5721), .Q(n3182) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n5676), .CK(n5721), .Q(n3181) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n5677), .CK(n5721), .Q(n3180) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n5678), .CK(n5721), .Q(n3179) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n5679), .CK(n5721), .Q(n3178) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n5680), .CK(n5721), .Q(n3177) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n5681), .CK(n5721), .Q(n3176) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n5682), .CK(n5721), .Q(n3175) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n5683), .CK(n5721), .Q(n3174) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n5684), .CK(n5721), .Q(n3173) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n5685), .CK(n5721), .Q(n3172) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n5686), .CK(n5721), .Q(n3171) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n5687), .CK(n5721), .Q(n3170) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n5688), .CK(n5721), .Q(n3169) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n5689), .CK(n5721), .Q(n3168) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n5690), .CK(n5721), .Q(n3167) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n5691), .CK(n5721), .Q(n3166) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n5692), .CK(n5721), .Q(n3165) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n5693), .CK(n5721), .Q(n3164) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n5694), .CK(n5721), .Q(n3163) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n5695), .CK(n5721), .Q(n3162) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n5696), .CK(n5721), .Q(n3161) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n5697), .CK(n5721), .Q(n3160) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n5698), .CK(n5721), .Q(n3159) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n5699), .CK(n5721), .Q(n3158) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n5700), .CK(n5721), .Q(n3157) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n5701), .CK(n5721), .Q(n3156) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n5702), .CK(n5721), .Q(n3155) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n5703), .CK(n5721), .Q(n3154) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n5704), .CK(n5721), .Q(n3153) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n5673), .CK(n5723), .Q(n3152) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n5674), .CK(n5723), .Q(n3151) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n5675), .CK(n5723), .Q(n3150) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n5676), .CK(n5723), .Q(n3149) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n5677), .CK(n5723), .Q(n3148) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n5678), .CK(n5723), .Q(n3147) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n5679), .CK(n5723), .Q(n3146) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n5680), .CK(n5723), .Q(n3145) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n5681), .CK(n5723), .Q(n3144) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n5682), .CK(n5723), .Q(n3143) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n5683), .CK(n5723), .Q(n3142) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n5684), .CK(n5723), .Q(n3141) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n5685), .CK(n5723), .Q(n3140) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n5686), .CK(n5723), .Q(n3139) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n5687), .CK(n5723), .Q(n3138) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n5688), .CK(n5723), .Q(n3137) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n5689), .CK(n5723), .Q(n3136) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n5690), .CK(n5723), .Q(n3135) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n5691), .CK(n5723), .Q(n3134) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n5692), .CK(n5723), .Q(n3133) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n5693), .CK(n5723), .Q(n3132) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n5694), .CK(n5723), .Q(n3131) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n5695), .CK(n5723), .Q(n3130) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n5696), .CK(n5723), .Q(n3129) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n5697), .CK(n5723), .Q(n3128) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n5698), .CK(n5723), .Q(n3127) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n5699), .CK(n5723), .Q(n3126) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n5700), .CK(n5723), .Q(n3125) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n5701), .CK(n5723), .Q(n3124) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n5702), .CK(n5723), .Q(n3123) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n5703), .CK(n5723), .Q(n3122) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n5704), .CK(n5723), .Q(n3121) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n5673), .CK(n5727), .Q(n3120) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n5674), .CK(n5727), .Q(n3119) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n5675), .CK(n5727), .Q(n3118) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n5676), .CK(n5727), .Q(n3117) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n5677), .CK(n5727), .Q(n3116) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n5678), .CK(n5727), .Q(n3115) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n5679), .CK(n5727), .Q(n3114) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n5680), .CK(n5727), .Q(n3113) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n5681), .CK(n5727), .Q(n3112) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n5682), .CK(n5727), .Q(n3111) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n5683), .CK(n5727), .Q(n3110) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n5684), .CK(n5727), .Q(n3109) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n5685), .CK(n5727), .Q(n3108) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n5686), .CK(n5727), .Q(n3107) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n5687), .CK(n5727), .Q(n3106) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n5688), .CK(n5727), .Q(n3105) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n5689), .CK(n5727), .Q(n3104) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n5690), .CK(n5727), .Q(n3103) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n5691), .CK(n5727), .Q(n3102) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n5692), .CK(n5727), .Q(n3101) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n5693), .CK(n5727), .Q(n3100) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n5694), .CK(n5727), .Q(n3099) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n5695), .CK(n5727), .Q(n3098) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n5696), .CK(n5727), .Q(n3097) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n5697), .CK(n5727), .Q(n3096) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n5698), .CK(n5727), .Q(n3095) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n5699), .CK(n5727), .Q(n3094) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n5700), .CK(n5727), .Q(n3093) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n5701), .CK(n5727), .Q(n3092) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n5702), .CK(n5727), .Q(n3091) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n5703), .CK(n5727), .Q(n3090) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n5704), .CK(n5727), .Q(n3089) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n5673), .CK(n5729), .QN(n5575) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n5674), .CK(n5729), .QN(n5576) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n5675), .CK(n5729), .QN(n5577) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n5676), .CK(n5729), .QN(n5578) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n5677), .CK(n5729), .QN(n5579) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n5678), .CK(n5729), .QN(n5580) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n5679), .CK(n5729), .QN(n5581) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n5680), .CK(n5729), .QN(n5582) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n5681), .CK(n5729), .QN(n5583) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n5682), .CK(n5729), .QN(n5584) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n5683), .CK(n5729), .QN(n5585) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n5684), .CK(n5729), .QN(n5586) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n5685), .CK(n5729), .QN(n5587) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n5686), .CK(n5729), .QN(n5588) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n5687), .CK(n5729), .QN(n5589) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n5688), .CK(n5729), .QN(n5590) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n5689), .CK(n5729), .QN(n5591) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n5690), .CK(n5729), .QN(n5592) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n5691), .CK(n5729), .QN(n5593) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n5692), .CK(n5729), .QN(n5594) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n5693), .CK(n5729), .QN(n5595) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n5694), .CK(n5729), .QN(n5596) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n5695), .CK(n5729), .QN(n5597) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n5696), .CK(n5729), .QN(n5598) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n5697), .CK(n5729), .QN(n5599) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n5698), .CK(n5729), .QN(n5600) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n5699), .CK(n5729), .QN(n5601) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n5700), .CK(n5729), .QN(n5602) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n5701), .CK(n5729), .QN(n5603) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n5702), .CK(n5729), .QN(n5604) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n5703), .CK(n5729), .QN(n5605) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n5704), .CK(n5729), .QN(n5606) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n5673), .CK(n5731), .Q(n3056) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n5674), .CK(n5731), .Q(n3055) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n5675), .CK(n5731), .Q(n3054) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n5676), .CK(n5731), .Q(n3053) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n5677), .CK(n5731), .Q(n3052) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n5678), .CK(n5731), .Q(n3051) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n5679), .CK(n5731), .Q(n3050) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n5680), .CK(n5731), .Q(n3049) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n5681), .CK(n5731), .Q(n3048) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n5682), .CK(n5731), .Q(n3047) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n5683), .CK(n5731), .Q(n3046) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n5684), .CK(n5731), .Q(n3045) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n5685), .CK(n5731), .Q(n3044) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n5686), .CK(n5731), .Q(n3043) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n5687), .CK(n5731), .Q(n3042) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n5688), .CK(n5731), .Q(n3041) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n5689), .CK(n5731), .Q(n3040) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n5690), .CK(n5731), .Q(n3039) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n5691), .CK(n5731), .Q(n3038) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n5692), .CK(n5731), .Q(n3037) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n5693), .CK(n5731), .Q(n3036) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n5694), .CK(n5731), .Q(n3035) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n5695), .CK(n5731), .Q(n3034) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n5696), .CK(n5731), .Q(n3033) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n5697), .CK(n5731), .Q(n3032) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n5698), .CK(n5731), .Q(n3031) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n5699), .CK(n5731), .Q(n3030) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n5700), .CK(n5731), .Q(n3029) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n5701), .CK(n5731), .Q(n3028) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n5702), .CK(n5731), .Q(n3027) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n5703), .CK(n5731), .Q(n3026) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n5704), .CK(n5731), .Q(n3025) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5673), .CK(n5733), .QN(n5161) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5674), .CK(n5733), .QN(n5165) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5675), .CK(n5733), .QN(n5169) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5676), .CK(n5733), .QN(n5173) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5677), .CK(n5733), .QN(n5177) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5678), .CK(n5733), .QN(n5181) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5679), .CK(n5733), .QN(n5185) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5680), .CK(n5733), .QN(n5189) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5681), .CK(n5733), .QN(n5193) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5682), .CK(n5733), .QN(n5197) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5683), .CK(n5733), .QN(n5201) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5684), .CK(n5733), .QN(n5205) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5685), .CK(n5733), .QN(n5209) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5686), .CK(n5733), .QN(n5213) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5687), .CK(n5733), .QN(n5217) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5688), .CK(n5733), .QN(n5221) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5689), .CK(n5733), .QN(n5225) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5690), .CK(n5733), .QN(n5229) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5691), .CK(n5733), .QN(n5233) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5692), .CK(n5733), .QN(n5237) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5693), .CK(n5733), .QN(n5241) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5694), .CK(n5733), .QN(n5245) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5695), .CK(n5733), .QN(n5249) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5696), .CK(n5733), .QN(n5253) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5697), .CK(n5733), .QN(n5257) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5698), .CK(n5733), .QN(n5261) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5699), .CK(n5733), .QN(n5265) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5700), .CK(n5733), .QN(n5269) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5701), .CK(n5733), .QN(n5273) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5702), .CK(n5733), .QN(n5277) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5703), .CK(n5733), .QN(n5281) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5704), .CK(n5733), .QN(n5285) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5673), .CK(n5735), .Q(n2992) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5674), .CK(n5735), .Q(n2991) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5675), .CK(n5735), .Q(n2990) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5676), .CK(n5735), .Q(n2989) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5677), .CK(n5735), .Q(n2988) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5678), .CK(n5735), .Q(n2987) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5679), .CK(n5735), .Q(n2986) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5680), .CK(n5735), .Q(n2985) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5681), .CK(n5735), .Q(n2984) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5682), .CK(n5735), .Q(n2983) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5683), .CK(n5735), .Q(n2982) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5684), .CK(n5735), .Q(n2981) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5685), .CK(n5735), .Q(n2980) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5686), .CK(n5735), .Q(n2979) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5687), .CK(n5735), .Q(n2978) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5688), .CK(n5735), .Q(n2977) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5689), .CK(n5735), .Q(n2976) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5690), .CK(n5735), .Q(n2975) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5691), .CK(n5735), .Q(n2974) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5692), .CK(n5735), .Q(n2973) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5693), .CK(n5735), .Q(n2972) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5694), .CK(n5735), .Q(n2971) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5695), .CK(n5735), .Q(n2970) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5696), .CK(n5735), .Q(n2969) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5697), .CK(n5735), .Q(n2968) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5698), .CK(n5735), .Q(n2967) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5699), .CK(n5735), .Q(n2966) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5700), .CK(n5735), .Q(n2965) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5701), .CK(n5735), .Q(n2964) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5702), .CK(n5735), .Q(n2963) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5703), .CK(n5735), .Q(n2962) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5704), .CK(n5735), .Q(n2961) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5673), .CK(n5737), .Q(n2960) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5674), .CK(n5737), .Q(n2959) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5675), .CK(n5737), .Q(n2958) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5676), .CK(n5737), .Q(n2957) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5677), .CK(n5737), .Q(n2956) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5678), .CK(n5737), .Q(n2955) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5679), .CK(n5737), .Q(n2954) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5680), .CK(n5737), .Q(n2953) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5681), .CK(n5737), .Q(n2952) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5682), .CK(n5737), .Q(n2951) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5683), .CK(n5737), .Q(n2950) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5684), .CK(n5737), .Q(n2949) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5685), .CK(n5737), .Q(n2948) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5686), .CK(n5737), .Q(n2947) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5687), .CK(n5737), .Q(n2946) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5688), .CK(n5737), .Q(n2945) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5689), .CK(n5737), .Q(n2944) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5690), .CK(n5737), .Q(n2943) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5691), .CK(n5737), .Q(n2942) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5692), .CK(n5737), .Q(n2941) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5693), .CK(n5737), .Q(n2940) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5694), .CK(n5737), .Q(n2939) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5695), .CK(n5737), .Q(n2938) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5696), .CK(n5737), .Q(n2937) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5697), .CK(n5737), .Q(n2936) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5698), .CK(n5737), .Q(n2935) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5699), .CK(n5737), .Q(n2934) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5700), .CK(n5737), .Q(n2933) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5701), .CK(n5737), .Q(n2932) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5702), .CK(n5737), .Q(n2931) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5703), .CK(n5737), .Q(n2930) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5704), .CK(n5737), .Q(n2929) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5673), .CK(n5739), .QN(n5607) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5674), .CK(n5739), .QN(n5608) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5675), .CK(n5739), .QN(n5609) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5676), .CK(n5739), .QN(n5610) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5677), .CK(n5739), .QN(n5611) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5678), .CK(n5739), .QN(n5612) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5679), .CK(n5739), .QN(n5613) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5680), .CK(n5739), .QN(n5614) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5681), .CK(n5739), .QN(n5615) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5682), .CK(n5739), .QN(n5616) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5683), .CK(n5739), .QN(n5617) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5684), .CK(n5739), .QN(n5618) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5685), .CK(n5739), .QN(n5619) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5686), .CK(n5739), .QN(n5620) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5687), .CK(n5739), .QN(n5621) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5688), .CK(n5739), .QN(n5622) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5689), .CK(n5739), .QN(n5623) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5690), .CK(n5739), .QN(n5624) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5691), .CK(n5739), .QN(n5625) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5692), .CK(n5739), .QN(n5626) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5693), .CK(n5739), .QN(n5627) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5694), .CK(n5739), .QN(n5628) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5695), .CK(n5739), .QN(n5629) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5696), .CK(n5739), .QN(n5630) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5697), .CK(n5739), .QN(n5631) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5698), .CK(n5739), .QN(n5632) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5699), .CK(n5739), .QN(n5633) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5700), .CK(n5739), .QN(n5634) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5701), .CK(n5739), .QN(n5635) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5702), .CK(n5739), .QN(n5636) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5703), .CK(n5739), .QN(n5637) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5704), .CK(n5739), .QN(n5638) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5673), .CK(n5741), .QN(n5639) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5674), .CK(n5741), .QN(n5640) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5675), .CK(n5741), .QN(n5641) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5676), .CK(n5741), .QN(n5642) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5677), .CK(n5741), .QN(n5643) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5678), .CK(n5741), .QN(n5644) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5679), .CK(n5741), .QN(n5645) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5680), .CK(n5741), .QN(n5646) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5681), .CK(n5741), .QN(n5647) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5682), .CK(n5741), .QN(n5648) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5683), .CK(n5741), .QN(n5649) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5684), .CK(n5741), .QN(n5650) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5685), .CK(n5741), .QN(n5651) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5686), .CK(n5741), .QN(n5652) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5687), .CK(n5741), .QN(n5653) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5688), .CK(n5741), .QN(n5654) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5689), .CK(n5741), .QN(n5655) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5690), .CK(n5741), .QN(n5656) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5691), .CK(n5741), .QN(n5657) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5692), .CK(n5741), .QN(n5658) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5693), .CK(n5741), .QN(n5659) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5694), .CK(n5741), .QN(n5660) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5695), .CK(n5741), .QN(n5661) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5696), .CK(n5741), .QN(n5662) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5697), .CK(n5741), .QN(n5663) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5698), .CK(n5741), .QN(n5664) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5699), .CK(n5741), .QN(n5665) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5700), .CK(n5741), .QN(n5666) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5701), .CK(n5741), .QN(n5667) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5702), .CK(n5741), .QN(n5668) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5703), .CK(n5741), .QN(n5669) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5704), .CK(n5741), .QN(n5670) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5673), .CK(n5743), .Q(n2864) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5674), .CK(n5743), .Q(n2863) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5675), .CK(n5743), .Q(n2862) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5676), .CK(n5743), .Q(n2861) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5677), .CK(n5743), .Q(n2860) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5678), .CK(n5743), .Q(n2859) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5679), .CK(n5743), .Q(n2858) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5680), .CK(n5743), .Q(n2857) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5681), .CK(n5743), .Q(n2856) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5682), .CK(n5743), .Q(n2855) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5683), .CK(n5743), .Q(n2854) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5684), .CK(n5743), .Q(n2853) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5685), .CK(n5743), .Q(n2852) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5686), .CK(n5743), .Q(n2851) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5687), .CK(n5743), .Q(n2850) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5688), .CK(n5743), .Q(n2849) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5689), .CK(n5743), .Q(n2848) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5690), .CK(n5743), .Q(n2847) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5691), .CK(n5743), .Q(n2846) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5692), .CK(n5743), .Q(n2845) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5693), .CK(n5743), .Q(n2844) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5694), .CK(n5743), .Q(n2843) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5695), .CK(n5743), .Q(n2842) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5696), .CK(n5743), .Q(n2841) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5697), .CK(n5743), .Q(n2840) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5698), .CK(n5743), .Q(n2839) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5699), .CK(n5743), .Q(n2838) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5700), .CK(n5743), .Q(n2837) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5701), .CK(n5743), .Q(n2836) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5702), .CK(n5743), .Q(n2835) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5703), .CK(n5743), .Q(n2834) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5704), .CK(n5743), .Q(n2833) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5673), .CK(n5745), .Q(n2832) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5674), .CK(n5745), .Q(n2831) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5675), .CK(n5745), .Q(n2830) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5676), .CK(n5745), .Q(n2829) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5677), .CK(n5745), .Q(n2828) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5678), .CK(n5745), .Q(n2827) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5679), .CK(n5745), .Q(n2826) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5680), .CK(n5745), .Q(n2825) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5681), .CK(n5745), .Q(n2824) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5682), .CK(n5745), .Q(n2823) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5683), .CK(n5745), .Q(n2822) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5684), .CK(n5745), .Q(n2821) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5685), .CK(n5745), .Q(n2820) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5686), .CK(n5745), .Q(n2819) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5687), .CK(n5745), .Q(n2818) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5688), .CK(n5745), .Q(n2817) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5689), .CK(n5745), .Q(n2816) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5690), .CK(n5745), .Q(n2815) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5691), .CK(n5745), .Q(n2814) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5692), .CK(n5745), .Q(n2813) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5693), .CK(n5745), .Q(n2812) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5694), .CK(n5745), .Q(n2811) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5695), .CK(n5745), .Q(n2810) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5696), .CK(n5745), .Q(n2809) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5697), .CK(n5745), .Q(n2808) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5698), .CK(n5745), .Q(n2807) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5699), .CK(n5745), .Q(n2806) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5700), .CK(n5745), .Q(n2805) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5701), .CK(n5745), .Q(n2804) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5702), .CK(n5745), .Q(n2803) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5703), .CK(n5745), .Q(n2802) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5704), .CK(n5745), .Q(n2801) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5673), .CK(n5749), .QN(n5162) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5674), .CK(n5749), .QN(n5166) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5675), .CK(n5749), .QN(n5170) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5676), .CK(n5749), .QN(n5174) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5677), .CK(n5749), .QN(n5178) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5678), .CK(n5749), .QN(n5182) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5679), .CK(n5749), .QN(n5186) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5680), .CK(n5749), .QN(n5190) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5681), .CK(n5749), .QN(n5194) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5682), .CK(n5749), .QN(n5198) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5683), .CK(n5749), .QN(n5202) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5684), .CK(n5749), .QN(n5206) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5685), .CK(n5749), .QN(n5210) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5686), .CK(n5749), .QN(n5214) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5687), .CK(n5749), .QN(n5218) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5688), .CK(n5749), .QN(n5222) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5689), .CK(n5749), .QN(n5226) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5690), .CK(n5749), .QN(n5230) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5691), .CK(n5749), .QN(n5234) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5692), .CK(n5749), .QN(n5238) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5693), .CK(n5749), .QN(n5242) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5694), .CK(n5749), .QN(n5246) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5695), .CK(n5749), .QN(n5250) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5696), .CK(n5749), .QN(n5254) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5697), .CK(n5749), .QN(n5258) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5698), .CK(n5749), .QN(n5262) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5699), .CK(n5749), .QN(n5266) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5700), .CK(n5749), .QN(n5270) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5701), .CK(n5749), .QN(n5274) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5702), .CK(n5749), .QN(n5278) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5703), .CK(n5749), .QN(n5282) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5704), .CK(n5749), .QN(n5286) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5673), .CK(n5751), .Q(n2768) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5674), .CK(n5751), .Q(n2767) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5675), .CK(n5751), .Q(n2766) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5676), .CK(n5751), .Q(n2765) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5677), .CK(n5751), .Q(n2764) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5678), .CK(n5751), .Q(n2763) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5679), .CK(n5751), .Q(n2762) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5680), .CK(n5751), .Q(n2761) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5681), .CK(n5751), .Q(n2760) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5682), .CK(n5751), .Q(n2759) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5683), .CK(n5751), .Q(n2758) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5684), .CK(n5751), .Q(n2757) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5685), .CK(n5751), .Q(n2756) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5686), .CK(n5751), .Q(n2755) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5687), .CK(n5751), .Q(n2754) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5688), .CK(n5751), .Q(n2753) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5689), .CK(n5751), .Q(n2752) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5690), .CK(n5751), .Q(n2751) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5691), .CK(n5751), .Q(n2750) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5692), .CK(n5751), .Q(n2749) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5693), .CK(n5751), .Q(n2748) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5694), .CK(n5751), .Q(n2747) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5695), .CK(n5751), .Q(n2746) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5696), .CK(n5751), .Q(n2745) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5697), .CK(n5751), .Q(n2744) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5698), .CK(n5751), .Q(n2743) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5699), .CK(n5751), .Q(n2742) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5700), .CK(n5751), .Q(n2741) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5701), .CK(n5751), .Q(n2740) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5702), .CK(n5751), .Q(n2739) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5703), .CK(n5751), .Q(n2738) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5704), .CK(n5751), .Q(n2737) );
  DLH_X1 \OUT1_reg[31]  ( .G(N444), .D(N410), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N444), .D(N409), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N444), .D(N408), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N444), .D(N407), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N444), .D(N406), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N444), .D(N405), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N444), .D(N404), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N444), .D(N403), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N444), .D(N402), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N444), .D(N401), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N444), .D(N400), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N444), .D(N399), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N444), .D(N398), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N444), .D(N397), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N444), .D(N396), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N444), .D(N395), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N444), .D(N394), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N444), .D(N393), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N444), .D(N392), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N444), .D(N391), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N444), .D(N390), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N444), .D(N389), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N444), .D(N388), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N444), .D(N387), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N444), .D(N386), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N444), .D(N385), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N444), .D(N384), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N444), .D(N383), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N444), .D(N382), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N444), .D(N381), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N444), .D(N380), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N444), .D(N379), .Q(OUT1[0]) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_0 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(n1032), .ENCLK(n5765), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_1 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(n1027), .ENCLK(n5763), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_2 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(n1063), .ENCLK(n5761), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_3 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(n1058), .ENCLK(n5759), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_4 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(n1053), .ENCLK(n5757), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_5 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(n1048), .ENCLK(n5755), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_6 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(n1043), .ENCLK(n5753), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_7 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(n1060), .ENCLK(n5751), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_8 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(n1055), .ENCLK(n5749), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_9 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(n1038), .ENCLK(n5747), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_10 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(n1050), .ENCLK(n5745), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_11 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(n1045), .ENCLK(n5743), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_12 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(n1040), .ENCLK(n5741), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_13 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(n1035), .ENCLK(n5739), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_14 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(n1030), .ENCLK(n5737), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_15 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(n1025), .ENCLK(n5735), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_16 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(n1061), .ENCLK(n5733), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_17 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(n1056), .ENCLK(n5731), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_18 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(n1051), .ENCLK(n5729), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_19 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(n1046), .ENCLK(n5727), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_20 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(n1033), .ENCLK(n5725), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_21 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(n1041), .ENCLK(n5723), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_22 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(n1036), .ENCLK(n5721), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_23 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(n1031), .ENCLK(n5719), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_24 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(n1026), .ENCLK(n5717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_25 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(n1062), .ENCLK(n5715), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_26 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(n1057), .ENCLK(n5713), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_27 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(n1052), .ENCLK(n5711), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_28 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(n1047), .ENCLK(n5709), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_29 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(n1042), .ENCLK(n5707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_30 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(n1037), .ENCLK(n5705), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_31 \clk_gate_REGISTERS_reg[0]  ( 
        .CLK(CLK), .EN(n1028), .ENCLK(n5671), .TE(1'b0) );
  AND2_X2 U3 ( .A1(n5136), .A2(n5145), .ZN(n4579) );
  AND2_X2 U4 ( .A1(n5134), .A2(n5145), .ZN(n4574) );
  AND2_X2 U5 ( .A1(n5132), .A2(n5135), .ZN(n4584) );
  AND2_X2 U6 ( .A1(n5136), .A2(n5139), .ZN(n4550) );
  AND2_X2 U7 ( .A1(n5142), .A2(n5143), .ZN(n4555) );
  AND2_X2 U8 ( .A1(n5134), .A2(n5142), .ZN(n4569) );
  AND2_X2 U9 ( .A1(n5139), .A2(n5143), .ZN(n4560) );
  NAND2_X2 U10 ( .A1(n5132), .A2(n5145), .ZN(n4571) );
  NAND2_X2 U11 ( .A1(n5132), .A2(n5140), .ZN(n4576) );
  NAND2_X2 U12 ( .A1(n5137), .A2(n5143), .ZN(n4557) );
  NAND2_X2 U13 ( .A1(n5136), .A2(n5144), .ZN(n4570) );
  NAND2_X2 U14 ( .A1(n5134), .A2(n5139), .ZN(n4575) );
  AND2_X2 U15 ( .A1(n5132), .A2(n5133), .ZN(n4545) );
  NAND2_X2 U16 ( .A1(n5145), .A2(n5143), .ZN(n4552) );
  NAND2_X2 U17 ( .A1(n5134), .A2(n5137), .ZN(n4541) );
  NAND2_X2 U18 ( .A1(n5136), .A2(n5140), .ZN(n4546) );
  NAND2_X2 U19 ( .A1(n5132), .A2(n5137), .ZN(n4581) );
  NAND2_X2 U20 ( .A1(n5136), .A2(n5135), .ZN(n4542) );
  NAND2_X2 U21 ( .A1(n5140), .A2(n5143), .ZN(n4551) );
  NAND2_X2 U22 ( .A1(n5134), .A2(n5144), .ZN(n4565) );
  NAND2_X2 U23 ( .A1(n5132), .A2(n5139), .ZN(n4547) );
  NAND2_X2 U24 ( .A1(n5136), .A2(n5137), .ZN(n4580) );
  NAND2_X2 U25 ( .A1(n5133), .A2(n5143), .ZN(n4556) );
  AND2_X2 U26 ( .A1(n5134), .A2(n5140), .ZN(n4578) );
  NAND2_X2 U27 ( .A1(n5132), .A2(n5142), .ZN(n4566) );
  AND2_X2 U28 ( .A1(n5136), .A2(n5133), .ZN(n4583) );
  AND2_X2 U29 ( .A1(n5134), .A2(n5135), .ZN(n4544) );
  AND2_X2 U30 ( .A1(n5144), .A2(n5143), .ZN(n4554) );
  INV_X2 U31 ( .A(RESET), .ZN(n4507) );
  AND2_X2 U32 ( .A1(n5136), .A2(n5142), .ZN(n4568) );
  AND2_X2 U33 ( .A1(n5132), .A2(n5144), .ZN(n4573) );
  AND2_X2 U34 ( .A1(n5134), .A2(n5133), .ZN(n4549) );
  AND2_X2 U35 ( .A1(n5135), .A2(n5143), .ZN(n4559) );
  AND2_X1 U36 ( .A1(DATAIN[31]), .A2(n4507), .ZN(n5673) );
  AND2_X1 U37 ( .A1(DATAIN[30]), .A2(n4507), .ZN(n5674) );
  AND2_X1 U38 ( .A1(DATAIN[29]), .A2(n4507), .ZN(n5675) );
  AND2_X1 U39 ( .A1(DATAIN[28]), .A2(n4507), .ZN(n5676) );
  AND2_X1 U40 ( .A1(DATAIN[27]), .A2(n4507), .ZN(n5677) );
  AND2_X1 U41 ( .A1(DATAIN[26]), .A2(n4507), .ZN(n5678) );
  AND2_X1 U42 ( .A1(DATAIN[25]), .A2(n4507), .ZN(n5679) );
  AND2_X1 U43 ( .A1(DATAIN[24]), .A2(n4507), .ZN(n5680) );
  AND2_X1 U44 ( .A1(DATAIN[23]), .A2(n4507), .ZN(n5681) );
  AND2_X1 U45 ( .A1(DATAIN[22]), .A2(n4507), .ZN(n5682) );
  AND2_X1 U46 ( .A1(DATAIN[21]), .A2(n4507), .ZN(n5683) );
  AND2_X1 U47 ( .A1(DATAIN[20]), .A2(n4507), .ZN(n5684) );
  AND2_X1 U48 ( .A1(DATAIN[19]), .A2(n4507), .ZN(n5685) );
  AND2_X1 U49 ( .A1(DATAIN[18]), .A2(n4507), .ZN(n5686) );
  AND2_X1 U50 ( .A1(DATAIN[17]), .A2(n4507), .ZN(n5687) );
  AND2_X1 U51 ( .A1(DATAIN[16]), .A2(n4507), .ZN(n5688) );
  AND2_X1 U52 ( .A1(DATAIN[15]), .A2(n4507), .ZN(n5689) );
  AND2_X1 U53 ( .A1(DATAIN[14]), .A2(n4507), .ZN(n5690) );
  AND2_X1 U54 ( .A1(DATAIN[13]), .A2(n4507), .ZN(n5691) );
  AND2_X1 U55 ( .A1(DATAIN[12]), .A2(n4507), .ZN(n5692) );
  AND2_X1 U56 ( .A1(DATAIN[11]), .A2(n4507), .ZN(n5693) );
  AND2_X1 U57 ( .A1(DATAIN[10]), .A2(n4507), .ZN(n5694) );
  AND2_X1 U58 ( .A1(DATAIN[9]), .A2(n4507), .ZN(n5695) );
  AND2_X1 U59 ( .A1(DATAIN[8]), .A2(n4507), .ZN(n5696) );
  AND2_X1 U60 ( .A1(DATAIN[7]), .A2(n4507), .ZN(n5697) );
  AND2_X1 U61 ( .A1(DATAIN[6]), .A2(n4507), .ZN(n5698) );
  AND2_X1 U62 ( .A1(DATAIN[5]), .A2(n4507), .ZN(n5699) );
  AND2_X1 U63 ( .A1(DATAIN[4]), .A2(n4507), .ZN(n5700) );
  AND2_X1 U64 ( .A1(DATAIN[3]), .A2(n4507), .ZN(n5701) );
  AND2_X1 U65 ( .A1(DATAIN[2]), .A2(n4507), .ZN(n5702) );
  AND2_X1 U66 ( .A1(DATAIN[1]), .A2(n4507), .ZN(n5703) );
  AND2_X1 U67 ( .A1(DATAIN[0]), .A2(n4507), .ZN(n5704) );
  NOR2_X1 U68 ( .A1(n4508), .A2(n4509), .ZN(n1063) );
  NOR2_X1 U69 ( .A1(n4510), .A2(n4509), .ZN(n1062) );
  NOR2_X1 U70 ( .A1(n4511), .A2(n4509), .ZN(n1061) );
  NOR2_X1 U71 ( .A1(n4512), .A2(n4509), .ZN(n1060) );
  OAI21_X1 U72 ( .B1(RESET), .B2(n4513), .A(n4514), .ZN(n4509) );
  NOR2_X1 U73 ( .A1(n4508), .A2(n4515), .ZN(n1058) );
  NOR2_X1 U74 ( .A1(n4510), .A2(n4515), .ZN(n1057) );
  NOR2_X1 U75 ( .A1(n4511), .A2(n4515), .ZN(n1056) );
  NOR2_X1 U76 ( .A1(n4512), .A2(n4515), .ZN(n1055) );
  OAI21_X1 U77 ( .B1(RESET), .B2(n4513), .A(n4516), .ZN(n4515) );
  NOR2_X1 U78 ( .A1(n4517), .A2(n4518), .ZN(n4513) );
  NOR2_X1 U79 ( .A1(n4508), .A2(n4519), .ZN(n1053) );
  NOR2_X1 U80 ( .A1(n4510), .A2(n4519), .ZN(n1052) );
  NOR2_X1 U81 ( .A1(n4511), .A2(n4519), .ZN(n1051) );
  NOR2_X1 U82 ( .A1(n4512), .A2(n4519), .ZN(n1050) );
  OAI21_X1 U83 ( .B1(RESET), .B2(n4520), .A(n4514), .ZN(n4519) );
  NOR2_X1 U84 ( .A1(n4508), .A2(n4521), .ZN(n1048) );
  NOR2_X1 U85 ( .A1(n4510), .A2(n4521), .ZN(n1047) );
  NOR2_X1 U86 ( .A1(n4511), .A2(n4521), .ZN(n1046) );
  NOR2_X1 U87 ( .A1(n4512), .A2(n4521), .ZN(n1045) );
  OAI21_X1 U88 ( .B1(RESET), .B2(n4520), .A(n4516), .ZN(n4521) );
  NOR2_X1 U89 ( .A1(n4517), .A2(ADD_WR[1]), .ZN(n4520) );
  INV_X1 U90 ( .A(ADD_WR[2]), .ZN(n4517) );
  NOR2_X1 U91 ( .A1(n4508), .A2(n4522), .ZN(n1043) );
  NOR2_X1 U92 ( .A1(n4510), .A2(n4522), .ZN(n1042) );
  NOR2_X1 U93 ( .A1(n4511), .A2(n4522), .ZN(n1041) );
  NOR2_X1 U94 ( .A1(n4512), .A2(n4522), .ZN(n1040) );
  OAI21_X1 U95 ( .B1(RESET), .B2(n4523), .A(n4514), .ZN(n4522) );
  NOR2_X1 U96 ( .A1(n4508), .A2(n4524), .ZN(n1038) );
  NOR2_X1 U97 ( .A1(n4510), .A2(n4524), .ZN(n1037) );
  NOR2_X1 U98 ( .A1(n4511), .A2(n4524), .ZN(n1036) );
  NOR2_X1 U99 ( .A1(n4512), .A2(n4524), .ZN(n1035) );
  OAI21_X1 U100 ( .B1(RESET), .B2(n4523), .A(n4516), .ZN(n4524) );
  NOR2_X1 U101 ( .A1(n4518), .A2(ADD_WR[2]), .ZN(n4523) );
  INV_X1 U102 ( .A(ADD_WR[1]), .ZN(n4518) );
  NOR2_X1 U103 ( .A1(n4508), .A2(n4525), .ZN(n1033) );
  NOR2_X1 U104 ( .A1(n4510), .A2(n4525), .ZN(n1032) );
  NOR2_X1 U105 ( .A1(n4511), .A2(n4525), .ZN(n1031) );
  NOR2_X1 U106 ( .A1(n4512), .A2(n4525), .ZN(n1030) );
  OAI21_X1 U107 ( .B1(RESET), .B2(n4526), .A(n4514), .ZN(n4525) );
  OR2_X1 U108 ( .A1(ADD_WR[0]), .A2(RESET), .ZN(n4514) );
  NOR2_X1 U109 ( .A1(n4508), .A2(n4527), .ZN(n1028) );
  AND2_X1 U110 ( .A1(n4507), .A2(n4528), .ZN(n4508) );
  NAND3_X1 U111 ( .A1(n4529), .A2(n4530), .A3(n4531), .ZN(n4528) );
  NOR2_X1 U112 ( .A1(n4510), .A2(n4527), .ZN(n1027) );
  AND2_X1 U113 ( .A1(n4507), .A2(n4532), .ZN(n4510) );
  NAND3_X1 U114 ( .A1(n4531), .A2(n4530), .A3(ADD_WR[3]), .ZN(n4532) );
  INV_X1 U115 ( .A(ADD_WR[4]), .ZN(n4530) );
  NOR2_X1 U116 ( .A1(n4511), .A2(n4527), .ZN(n1026) );
  AND2_X1 U117 ( .A1(n4507), .A2(n4533), .ZN(n4511) );
  NAND3_X1 U118 ( .A1(n4531), .A2(n4529), .A3(ADD_WR[4]), .ZN(n4533) );
  INV_X1 U119 ( .A(ADD_WR[3]), .ZN(n4529) );
  NOR2_X1 U120 ( .A1(n4512), .A2(n4527), .ZN(n1025) );
  OAI21_X1 U121 ( .B1(RESET), .B2(n4526), .A(n4516), .ZN(n4527) );
  NAND2_X1 U122 ( .A1(ADD_WR[0]), .A2(n4507), .ZN(n4516) );
  NOR2_X1 U123 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n4526) );
  AND2_X1 U124 ( .A1(n4507), .A2(n4534), .ZN(n4512) );
  NAND3_X1 U125 ( .A1(ADD_WR[3]), .A2(n4531), .A3(ADD_WR[4]), .ZN(n4534) );
  AND2_X1 U126 ( .A1(WR), .A2(ENABLE), .ZN(n4531) );
  AND2_X1 U127 ( .A1(RD1), .A2(ENABLE), .ZN(N444) );
  NAND2_X1 U128 ( .A1(n4535), .A2(n4536), .ZN(N410) );
  NOR4_X1 U129 ( .A1(n4537), .A2(n4538), .A3(n4539), .A4(n4540), .ZN(n4536) );
  OAI221_X1 U130 ( .B1(n5351), .B2(n4541), .C1(n5479), .C2(n4542), .A(n4543), 
        .ZN(n4540) );
  AOI22_X1 U131 ( .A1(n4544), .A2(n3408), .B1(n4545), .B2(n3184), .ZN(n4543)
         );
  OAI221_X1 U132 ( .B1(n5415), .B2(n4546), .C1(n5607), .C2(n4547), .A(n4548), 
        .ZN(n4539) );
  AOI22_X1 U133 ( .A1(n4549), .A2(n3152), .B1(n4550), .B2(n2960), .ZN(n4548)
         );
  OAI221_X1 U134 ( .B1(n5383), .B2(n4551), .C1(n5511), .C2(n4552), .A(n4553), 
        .ZN(n4538) );
  AOI22_X1 U135 ( .A1(n4554), .A2(n3120), .B1(n4555), .B2(n2864), .ZN(n4553)
         );
  OAI221_X1 U136 ( .B1(n5543), .B2(n4556), .C1(n5287), .C2(n4557), .A(n4558), 
        .ZN(n4537) );
  AOI22_X1 U137 ( .A1(n4559), .A2(n3504), .B1(n4560), .B2(n2992), .ZN(n4558)
         );
  NOR4_X1 U138 ( .A1(n4561), .A2(n4562), .A3(n4563), .A4(n4564), .ZN(n4535) );
  OAI221_X1 U139 ( .B1(n5161), .B2(n4565), .C1(n5162), .C2(n4566), .A(n4567), 
        .ZN(n4564) );
  AOI22_X1 U140 ( .A1(n4568), .A2(n2832), .B1(n4569), .B2(n2768), .ZN(n4567)
         );
  OAI221_X1 U141 ( .B1(n5575), .B2(n4570), .C1(n5160), .C2(n4571), .A(n4572), 
        .ZN(n4563) );
  AOI22_X1 U142 ( .A1(n4573), .A2(n3056), .B1(n4574), .B2(n3280), .ZN(n4572)
         );
  OAI221_X1 U143 ( .B1(n5639), .B2(n4575), .C1(n5447), .C2(n4576), .A(n4577), 
        .ZN(n4562) );
  AOI22_X1 U144 ( .A1(n4578), .A2(n3536), .B1(n4579), .B2(n3344), .ZN(n4577)
         );
  OAI221_X1 U145 ( .B1(n5159), .B2(n4580), .C1(n5319), .C2(n4581), .A(n4582), 
        .ZN(n4561) );
  AOI22_X1 U146 ( .A1(n4583), .A2(n3216), .B1(n4584), .B2(n3440), .ZN(n4582)
         );
  NAND2_X1 U147 ( .A1(n4585), .A2(n4586), .ZN(N409) );
  NOR4_X1 U148 ( .A1(n4587), .A2(n4588), .A3(n4589), .A4(n4590), .ZN(n4586) );
  OAI221_X1 U149 ( .B1(n5352), .B2(n4541), .C1(n5480), .C2(n4542), .A(n4591), 
        .ZN(n4590) );
  AOI22_X1 U150 ( .A1(n4544), .A2(n3407), .B1(n4545), .B2(n3183), .ZN(n4591)
         );
  OAI221_X1 U151 ( .B1(n5416), .B2(n4546), .C1(n5608), .C2(n4547), .A(n4592), 
        .ZN(n4589) );
  AOI22_X1 U152 ( .A1(n4549), .A2(n3151), .B1(n4550), .B2(n2959), .ZN(n4592)
         );
  OAI221_X1 U153 ( .B1(n5384), .B2(n4551), .C1(n5512), .C2(n4552), .A(n4593), 
        .ZN(n4588) );
  AOI22_X1 U154 ( .A1(n4554), .A2(n3119), .B1(n4555), .B2(n2863), .ZN(n4593)
         );
  OAI221_X1 U155 ( .B1(n5544), .B2(n4556), .C1(n5288), .C2(n4557), .A(n4594), 
        .ZN(n4587) );
  AOI22_X1 U156 ( .A1(n4559), .A2(n3503), .B1(n4560), .B2(n2991), .ZN(n4594)
         );
  NOR4_X1 U157 ( .A1(n4595), .A2(n4596), .A3(n4597), .A4(n4598), .ZN(n4585) );
  OAI221_X1 U158 ( .B1(n5165), .B2(n4565), .C1(n5166), .C2(n4566), .A(n4599), 
        .ZN(n4598) );
  AOI22_X1 U159 ( .A1(n4568), .A2(n2831), .B1(n4569), .B2(n2767), .ZN(n4599)
         );
  OAI221_X1 U160 ( .B1(n5576), .B2(n4570), .C1(n5164), .C2(n4571), .A(n4600), 
        .ZN(n4597) );
  AOI22_X1 U161 ( .A1(n4573), .A2(n3055), .B1(n4574), .B2(n3279), .ZN(n4600)
         );
  OAI221_X1 U162 ( .B1(n5640), .B2(n4575), .C1(n5448), .C2(n4576), .A(n4601), 
        .ZN(n4596) );
  AOI22_X1 U163 ( .A1(n4578), .A2(n3535), .B1(n4579), .B2(n3343), .ZN(n4601)
         );
  OAI221_X1 U164 ( .B1(n5163), .B2(n4580), .C1(n5320), .C2(n4581), .A(n4602), 
        .ZN(n4595) );
  AOI22_X1 U165 ( .A1(n4583), .A2(n3215), .B1(n4584), .B2(n3439), .ZN(n4602)
         );
  NAND2_X1 U166 ( .A1(n4603), .A2(n4604), .ZN(N408) );
  NOR4_X1 U167 ( .A1(n4605), .A2(n4606), .A3(n4607), .A4(n4608), .ZN(n4604) );
  OAI221_X1 U168 ( .B1(n5353), .B2(n4541), .C1(n5481), .C2(n4542), .A(n4609), 
        .ZN(n4608) );
  AOI22_X1 U169 ( .A1(n4544), .A2(n3406), .B1(n4545), .B2(n3182), .ZN(n4609)
         );
  OAI221_X1 U170 ( .B1(n5417), .B2(n4546), .C1(n5609), .C2(n4547), .A(n4610), 
        .ZN(n4607) );
  AOI22_X1 U171 ( .A1(n4549), .A2(n3150), .B1(n4550), .B2(n2958), .ZN(n4610)
         );
  OAI221_X1 U172 ( .B1(n5385), .B2(n4551), .C1(n5513), .C2(n4552), .A(n4611), 
        .ZN(n4606) );
  AOI22_X1 U173 ( .A1(n4554), .A2(n3118), .B1(n4555), .B2(n2862), .ZN(n4611)
         );
  OAI221_X1 U174 ( .B1(n5545), .B2(n4556), .C1(n5289), .C2(n4557), .A(n4612), 
        .ZN(n4605) );
  AOI22_X1 U175 ( .A1(n4559), .A2(n3502), .B1(n4560), .B2(n2990), .ZN(n4612)
         );
  NOR4_X1 U176 ( .A1(n4613), .A2(n4614), .A3(n4615), .A4(n4616), .ZN(n4603) );
  OAI221_X1 U177 ( .B1(n5169), .B2(n4565), .C1(n5170), .C2(n4566), .A(n4617), 
        .ZN(n4616) );
  AOI22_X1 U178 ( .A1(n4568), .A2(n2830), .B1(n4569), .B2(n2766), .ZN(n4617)
         );
  OAI221_X1 U179 ( .B1(n5577), .B2(n4570), .C1(n5168), .C2(n4571), .A(n4618), 
        .ZN(n4615) );
  AOI22_X1 U180 ( .A1(n4573), .A2(n3054), .B1(n4574), .B2(n3278), .ZN(n4618)
         );
  OAI221_X1 U181 ( .B1(n5641), .B2(n4575), .C1(n5449), .C2(n4576), .A(n4619), 
        .ZN(n4614) );
  AOI22_X1 U182 ( .A1(n4578), .A2(n3534), .B1(n4579), .B2(n3342), .ZN(n4619)
         );
  OAI221_X1 U183 ( .B1(n5167), .B2(n4580), .C1(n5321), .C2(n4581), .A(n4620), 
        .ZN(n4613) );
  AOI22_X1 U184 ( .A1(n4583), .A2(n3214), .B1(n4584), .B2(n3438), .ZN(n4620)
         );
  NAND2_X1 U185 ( .A1(n4621), .A2(n4622), .ZN(N407) );
  NOR4_X1 U186 ( .A1(n4623), .A2(n4624), .A3(n4625), .A4(n4626), .ZN(n4622) );
  OAI221_X1 U187 ( .B1(n5354), .B2(n4541), .C1(n5482), .C2(n4542), .A(n4627), 
        .ZN(n4626) );
  AOI22_X1 U188 ( .A1(n4544), .A2(n3405), .B1(n4545), .B2(n3181), .ZN(n4627)
         );
  OAI221_X1 U189 ( .B1(n5418), .B2(n4546), .C1(n5610), .C2(n4547), .A(n4628), 
        .ZN(n4625) );
  AOI22_X1 U190 ( .A1(n4549), .A2(n3149), .B1(n4550), .B2(n2957), .ZN(n4628)
         );
  OAI221_X1 U191 ( .B1(n5386), .B2(n4551), .C1(n5514), .C2(n4552), .A(n4629), 
        .ZN(n4624) );
  AOI22_X1 U192 ( .A1(n4554), .A2(n3117), .B1(n4555), .B2(n2861), .ZN(n4629)
         );
  OAI221_X1 U193 ( .B1(n5546), .B2(n4556), .C1(n5290), .C2(n4557), .A(n4630), 
        .ZN(n4623) );
  AOI22_X1 U194 ( .A1(n4559), .A2(n3501), .B1(n4560), .B2(n2989), .ZN(n4630)
         );
  NOR4_X1 U195 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n4621) );
  OAI221_X1 U196 ( .B1(n5173), .B2(n4565), .C1(n5174), .C2(n4566), .A(n4635), 
        .ZN(n4634) );
  AOI22_X1 U197 ( .A1(n4568), .A2(n2829), .B1(n4569), .B2(n2765), .ZN(n4635)
         );
  OAI221_X1 U198 ( .B1(n5578), .B2(n4570), .C1(n5172), .C2(n4571), .A(n4636), 
        .ZN(n4633) );
  AOI22_X1 U199 ( .A1(n4573), .A2(n3053), .B1(n4574), .B2(n3277), .ZN(n4636)
         );
  OAI221_X1 U200 ( .B1(n5642), .B2(n4575), .C1(n5450), .C2(n4576), .A(n4637), 
        .ZN(n4632) );
  AOI22_X1 U201 ( .A1(n4578), .A2(n3533), .B1(n4579), .B2(n3341), .ZN(n4637)
         );
  OAI221_X1 U202 ( .B1(n5171), .B2(n4580), .C1(n5322), .C2(n4581), .A(n4638), 
        .ZN(n4631) );
  AOI22_X1 U203 ( .A1(n4583), .A2(n3213), .B1(n4584), .B2(n3437), .ZN(n4638)
         );
  NAND2_X1 U204 ( .A1(n4639), .A2(n4640), .ZN(N406) );
  NOR4_X1 U205 ( .A1(n4641), .A2(n4642), .A3(n4643), .A4(n4644), .ZN(n4640) );
  OAI221_X1 U206 ( .B1(n5355), .B2(n4541), .C1(n5483), .C2(n4542), .A(n4645), 
        .ZN(n4644) );
  AOI22_X1 U207 ( .A1(n4544), .A2(n3404), .B1(n4545), .B2(n3180), .ZN(n4645)
         );
  OAI221_X1 U208 ( .B1(n5419), .B2(n4546), .C1(n5611), .C2(n4547), .A(n4646), 
        .ZN(n4643) );
  AOI22_X1 U209 ( .A1(n4549), .A2(n3148), .B1(n4550), .B2(n2956), .ZN(n4646)
         );
  OAI221_X1 U210 ( .B1(n5387), .B2(n4551), .C1(n5515), .C2(n4552), .A(n4647), 
        .ZN(n4642) );
  AOI22_X1 U211 ( .A1(n4554), .A2(n3116), .B1(n4555), .B2(n2860), .ZN(n4647)
         );
  OAI221_X1 U212 ( .B1(n5547), .B2(n4556), .C1(n5291), .C2(n4557), .A(n4648), 
        .ZN(n4641) );
  AOI22_X1 U213 ( .A1(n4559), .A2(n3500), .B1(n4560), .B2(n2988), .ZN(n4648)
         );
  NOR4_X1 U214 ( .A1(n4649), .A2(n4650), .A3(n4651), .A4(n4652), .ZN(n4639) );
  OAI221_X1 U215 ( .B1(n5177), .B2(n4565), .C1(n5178), .C2(n4566), .A(n4653), 
        .ZN(n4652) );
  AOI22_X1 U216 ( .A1(n4568), .A2(n2828), .B1(n4569), .B2(n2764), .ZN(n4653)
         );
  OAI221_X1 U217 ( .B1(n5579), .B2(n4570), .C1(n5176), .C2(n4571), .A(n4654), 
        .ZN(n4651) );
  AOI22_X1 U218 ( .A1(n4573), .A2(n3052), .B1(n4574), .B2(n3276), .ZN(n4654)
         );
  OAI221_X1 U219 ( .B1(n5643), .B2(n4575), .C1(n5451), .C2(n4576), .A(n4655), 
        .ZN(n4650) );
  AOI22_X1 U220 ( .A1(n4578), .A2(n3532), .B1(n4579), .B2(n3340), .ZN(n4655)
         );
  OAI221_X1 U221 ( .B1(n5175), .B2(n4580), .C1(n5323), .C2(n4581), .A(n4656), 
        .ZN(n4649) );
  AOI22_X1 U222 ( .A1(n4583), .A2(n3212), .B1(n4584), .B2(n3436), .ZN(n4656)
         );
  NAND2_X1 U223 ( .A1(n4657), .A2(n4658), .ZN(N405) );
  NOR4_X1 U224 ( .A1(n4659), .A2(n4660), .A3(n4661), .A4(n4662), .ZN(n4658) );
  OAI221_X1 U225 ( .B1(n5356), .B2(n4541), .C1(n5484), .C2(n4542), .A(n4663), 
        .ZN(n4662) );
  AOI22_X1 U226 ( .A1(n4544), .A2(n3403), .B1(n4545), .B2(n3179), .ZN(n4663)
         );
  OAI221_X1 U227 ( .B1(n5420), .B2(n4546), .C1(n5612), .C2(n4547), .A(n4664), 
        .ZN(n4661) );
  AOI22_X1 U228 ( .A1(n4549), .A2(n3147), .B1(n4550), .B2(n2955), .ZN(n4664)
         );
  OAI221_X1 U229 ( .B1(n5388), .B2(n4551), .C1(n5516), .C2(n4552), .A(n4665), 
        .ZN(n4660) );
  AOI22_X1 U230 ( .A1(n4554), .A2(n3115), .B1(n4555), .B2(n2859), .ZN(n4665)
         );
  OAI221_X1 U231 ( .B1(n5548), .B2(n4556), .C1(n5292), .C2(n4557), .A(n4666), 
        .ZN(n4659) );
  AOI22_X1 U232 ( .A1(n4559), .A2(n3499), .B1(n4560), .B2(n2987), .ZN(n4666)
         );
  NOR4_X1 U233 ( .A1(n4667), .A2(n4668), .A3(n4669), .A4(n4670), .ZN(n4657) );
  OAI221_X1 U234 ( .B1(n5181), .B2(n4565), .C1(n5182), .C2(n4566), .A(n4671), 
        .ZN(n4670) );
  AOI22_X1 U235 ( .A1(n4568), .A2(n2827), .B1(n4569), .B2(n2763), .ZN(n4671)
         );
  OAI221_X1 U236 ( .B1(n5580), .B2(n4570), .C1(n5180), .C2(n4571), .A(n4672), 
        .ZN(n4669) );
  AOI22_X1 U237 ( .A1(n4573), .A2(n3051), .B1(n4574), .B2(n3275), .ZN(n4672)
         );
  OAI221_X1 U238 ( .B1(n5644), .B2(n4575), .C1(n5452), .C2(n4576), .A(n4673), 
        .ZN(n4668) );
  AOI22_X1 U239 ( .A1(n4578), .A2(n3531), .B1(n4579), .B2(n3339), .ZN(n4673)
         );
  OAI221_X1 U240 ( .B1(n5179), .B2(n4580), .C1(n5324), .C2(n4581), .A(n4674), 
        .ZN(n4667) );
  AOI22_X1 U241 ( .A1(n4583), .A2(n3211), .B1(n4584), .B2(n3435), .ZN(n4674)
         );
  NAND2_X1 U242 ( .A1(n4675), .A2(n4676), .ZN(N404) );
  NOR4_X1 U243 ( .A1(n4677), .A2(n4678), .A3(n4679), .A4(n4680), .ZN(n4676) );
  OAI221_X1 U244 ( .B1(n5357), .B2(n4541), .C1(n5485), .C2(n4542), .A(n4681), 
        .ZN(n4680) );
  AOI22_X1 U245 ( .A1(n4544), .A2(n3402), .B1(n4545), .B2(n3178), .ZN(n4681)
         );
  OAI221_X1 U246 ( .B1(n5421), .B2(n4546), .C1(n5613), .C2(n4547), .A(n4682), 
        .ZN(n4679) );
  AOI22_X1 U247 ( .A1(n4549), .A2(n3146), .B1(n4550), .B2(n2954), .ZN(n4682)
         );
  OAI221_X1 U248 ( .B1(n5389), .B2(n4551), .C1(n5517), .C2(n4552), .A(n4683), 
        .ZN(n4678) );
  AOI22_X1 U249 ( .A1(n4554), .A2(n3114), .B1(n4555), .B2(n2858), .ZN(n4683)
         );
  OAI221_X1 U250 ( .B1(n5549), .B2(n4556), .C1(n5293), .C2(n4557), .A(n4684), 
        .ZN(n4677) );
  AOI22_X1 U251 ( .A1(n4559), .A2(n3498), .B1(n4560), .B2(n2986), .ZN(n4684)
         );
  NOR4_X1 U252 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .ZN(n4675) );
  OAI221_X1 U253 ( .B1(n5185), .B2(n4565), .C1(n5186), .C2(n4566), .A(n4689), 
        .ZN(n4688) );
  AOI22_X1 U254 ( .A1(n4568), .A2(n2826), .B1(n4569), .B2(n2762), .ZN(n4689)
         );
  OAI221_X1 U255 ( .B1(n5581), .B2(n4570), .C1(n5184), .C2(n4571), .A(n4690), 
        .ZN(n4687) );
  AOI22_X1 U256 ( .A1(n4573), .A2(n3050), .B1(n4574), .B2(n3274), .ZN(n4690)
         );
  OAI221_X1 U257 ( .B1(n5645), .B2(n4575), .C1(n5453), .C2(n4576), .A(n4691), 
        .ZN(n4686) );
  AOI22_X1 U258 ( .A1(n4578), .A2(n3530), .B1(n4579), .B2(n3338), .ZN(n4691)
         );
  OAI221_X1 U259 ( .B1(n5183), .B2(n4580), .C1(n5325), .C2(n4581), .A(n4692), 
        .ZN(n4685) );
  AOI22_X1 U260 ( .A1(n4583), .A2(n3210), .B1(n4584), .B2(n3434), .ZN(n4692)
         );
  NAND2_X1 U261 ( .A1(n4693), .A2(n4694), .ZN(N403) );
  NOR4_X1 U262 ( .A1(n4695), .A2(n4696), .A3(n4697), .A4(n4698), .ZN(n4694) );
  OAI221_X1 U263 ( .B1(n5358), .B2(n4541), .C1(n5486), .C2(n4542), .A(n4699), 
        .ZN(n4698) );
  AOI22_X1 U264 ( .A1(n4544), .A2(n3401), .B1(n4545), .B2(n3177), .ZN(n4699)
         );
  OAI221_X1 U265 ( .B1(n5422), .B2(n4546), .C1(n5614), .C2(n4547), .A(n4700), 
        .ZN(n4697) );
  AOI22_X1 U266 ( .A1(n4549), .A2(n3145), .B1(n4550), .B2(n2953), .ZN(n4700)
         );
  OAI221_X1 U267 ( .B1(n5390), .B2(n4551), .C1(n5518), .C2(n4552), .A(n4701), 
        .ZN(n4696) );
  AOI22_X1 U268 ( .A1(n4554), .A2(n3113), .B1(n4555), .B2(n2857), .ZN(n4701)
         );
  OAI221_X1 U269 ( .B1(n5550), .B2(n4556), .C1(n5294), .C2(n4557), .A(n4702), 
        .ZN(n4695) );
  AOI22_X1 U270 ( .A1(n4559), .A2(n3497), .B1(n4560), .B2(n2985), .ZN(n4702)
         );
  NOR4_X1 U271 ( .A1(n4703), .A2(n4704), .A3(n4705), .A4(n4706), .ZN(n4693) );
  OAI221_X1 U272 ( .B1(n5189), .B2(n4565), .C1(n5190), .C2(n4566), .A(n4707), 
        .ZN(n4706) );
  AOI22_X1 U273 ( .A1(n4568), .A2(n2825), .B1(n4569), .B2(n2761), .ZN(n4707)
         );
  OAI221_X1 U274 ( .B1(n5582), .B2(n4570), .C1(n5188), .C2(n4571), .A(n4708), 
        .ZN(n4705) );
  AOI22_X1 U275 ( .A1(n4573), .A2(n3049), .B1(n4574), .B2(n3273), .ZN(n4708)
         );
  OAI221_X1 U276 ( .B1(n5646), .B2(n4575), .C1(n5454), .C2(n4576), .A(n4709), 
        .ZN(n4704) );
  AOI22_X1 U277 ( .A1(n4578), .A2(n3529), .B1(n4579), .B2(n3337), .ZN(n4709)
         );
  OAI221_X1 U278 ( .B1(n5187), .B2(n4580), .C1(n5326), .C2(n4581), .A(n4710), 
        .ZN(n4703) );
  AOI22_X1 U279 ( .A1(n4583), .A2(n3209), .B1(n4584), .B2(n3433), .ZN(n4710)
         );
  NAND2_X1 U280 ( .A1(n4711), .A2(n4712), .ZN(N402) );
  NOR4_X1 U281 ( .A1(n4713), .A2(n4714), .A3(n4715), .A4(n4716), .ZN(n4712) );
  OAI221_X1 U282 ( .B1(n5359), .B2(n4541), .C1(n5487), .C2(n4542), .A(n4717), 
        .ZN(n4716) );
  AOI22_X1 U283 ( .A1(n4544), .A2(n3400), .B1(n4545), .B2(n3176), .ZN(n4717)
         );
  OAI221_X1 U284 ( .B1(n5423), .B2(n4546), .C1(n5615), .C2(n4547), .A(n4718), 
        .ZN(n4715) );
  AOI22_X1 U285 ( .A1(n4549), .A2(n3144), .B1(n4550), .B2(n2952), .ZN(n4718)
         );
  OAI221_X1 U286 ( .B1(n5391), .B2(n4551), .C1(n5519), .C2(n4552), .A(n4719), 
        .ZN(n4714) );
  AOI22_X1 U287 ( .A1(n4554), .A2(n3112), .B1(n4555), .B2(n2856), .ZN(n4719)
         );
  OAI221_X1 U288 ( .B1(n5551), .B2(n4556), .C1(n5295), .C2(n4557), .A(n4720), 
        .ZN(n4713) );
  AOI22_X1 U289 ( .A1(n4559), .A2(n3496), .B1(n4560), .B2(n2984), .ZN(n4720)
         );
  NOR4_X1 U290 ( .A1(n4721), .A2(n4722), .A3(n4723), .A4(n4724), .ZN(n4711) );
  OAI221_X1 U291 ( .B1(n5193), .B2(n4565), .C1(n5194), .C2(n4566), .A(n4725), 
        .ZN(n4724) );
  AOI22_X1 U292 ( .A1(n4568), .A2(n2824), .B1(n4569), .B2(n2760), .ZN(n4725)
         );
  OAI221_X1 U293 ( .B1(n5583), .B2(n4570), .C1(n5192), .C2(n4571), .A(n4726), 
        .ZN(n4723) );
  AOI22_X1 U294 ( .A1(n4573), .A2(n3048), .B1(n4574), .B2(n3272), .ZN(n4726)
         );
  OAI221_X1 U295 ( .B1(n5647), .B2(n4575), .C1(n5455), .C2(n4576), .A(n4727), 
        .ZN(n4722) );
  AOI22_X1 U296 ( .A1(n4578), .A2(n3528), .B1(n4579), .B2(n3336), .ZN(n4727)
         );
  OAI221_X1 U297 ( .B1(n5191), .B2(n4580), .C1(n5327), .C2(n4581), .A(n4728), 
        .ZN(n4721) );
  AOI22_X1 U298 ( .A1(n4583), .A2(n3208), .B1(n4584), .B2(n3432), .ZN(n4728)
         );
  NAND2_X1 U299 ( .A1(n4729), .A2(n4730), .ZN(N401) );
  NOR4_X1 U300 ( .A1(n4731), .A2(n4732), .A3(n4733), .A4(n4734), .ZN(n4730) );
  OAI221_X1 U301 ( .B1(n5360), .B2(n4541), .C1(n5488), .C2(n4542), .A(n4735), 
        .ZN(n4734) );
  AOI22_X1 U302 ( .A1(n4544), .A2(n3399), .B1(n4545), .B2(n3175), .ZN(n4735)
         );
  OAI221_X1 U303 ( .B1(n5424), .B2(n4546), .C1(n5616), .C2(n4547), .A(n4736), 
        .ZN(n4733) );
  AOI22_X1 U304 ( .A1(n4549), .A2(n3143), .B1(n4550), .B2(n2951), .ZN(n4736)
         );
  OAI221_X1 U305 ( .B1(n5392), .B2(n4551), .C1(n5520), .C2(n4552), .A(n4737), 
        .ZN(n4732) );
  AOI22_X1 U306 ( .A1(n4554), .A2(n3111), .B1(n4555), .B2(n2855), .ZN(n4737)
         );
  OAI221_X1 U307 ( .B1(n5552), .B2(n4556), .C1(n5296), .C2(n4557), .A(n4738), 
        .ZN(n4731) );
  AOI22_X1 U308 ( .A1(n4559), .A2(n3495), .B1(n4560), .B2(n2983), .ZN(n4738)
         );
  NOR4_X1 U309 ( .A1(n4739), .A2(n4740), .A3(n4741), .A4(n4742), .ZN(n4729) );
  OAI221_X1 U310 ( .B1(n5197), .B2(n4565), .C1(n5198), .C2(n4566), .A(n4743), 
        .ZN(n4742) );
  AOI22_X1 U311 ( .A1(n4568), .A2(n2823), .B1(n4569), .B2(n2759), .ZN(n4743)
         );
  OAI221_X1 U312 ( .B1(n5584), .B2(n4570), .C1(n5196), .C2(n4571), .A(n4744), 
        .ZN(n4741) );
  AOI22_X1 U313 ( .A1(n4573), .A2(n3047), .B1(n4574), .B2(n3271), .ZN(n4744)
         );
  OAI221_X1 U314 ( .B1(n5648), .B2(n4575), .C1(n5456), .C2(n4576), .A(n4745), 
        .ZN(n4740) );
  AOI22_X1 U315 ( .A1(n4578), .A2(n3527), .B1(n4579), .B2(n3335), .ZN(n4745)
         );
  OAI221_X1 U316 ( .B1(n5195), .B2(n4580), .C1(n5328), .C2(n4581), .A(n4746), 
        .ZN(n4739) );
  AOI22_X1 U317 ( .A1(n4583), .A2(n3207), .B1(n4584), .B2(n3431), .ZN(n4746)
         );
  NAND2_X1 U318 ( .A1(n4747), .A2(n4748), .ZN(N400) );
  NOR4_X1 U319 ( .A1(n4749), .A2(n4750), .A3(n4751), .A4(n4752), .ZN(n4748) );
  OAI221_X1 U320 ( .B1(n5361), .B2(n4541), .C1(n5489), .C2(n4542), .A(n4753), 
        .ZN(n4752) );
  AOI22_X1 U321 ( .A1(n4544), .A2(n3398), .B1(n4545), .B2(n3174), .ZN(n4753)
         );
  OAI221_X1 U322 ( .B1(n5425), .B2(n4546), .C1(n5617), .C2(n4547), .A(n4754), 
        .ZN(n4751) );
  AOI22_X1 U323 ( .A1(n4549), .A2(n3142), .B1(n4550), .B2(n2950), .ZN(n4754)
         );
  OAI221_X1 U324 ( .B1(n5393), .B2(n4551), .C1(n5521), .C2(n4552), .A(n4755), 
        .ZN(n4750) );
  AOI22_X1 U325 ( .A1(n4554), .A2(n3110), .B1(n4555), .B2(n2854), .ZN(n4755)
         );
  OAI221_X1 U326 ( .B1(n5553), .B2(n4556), .C1(n5297), .C2(n4557), .A(n4756), 
        .ZN(n4749) );
  AOI22_X1 U327 ( .A1(n4559), .A2(n3494), .B1(n4560), .B2(n2982), .ZN(n4756)
         );
  NOR4_X1 U328 ( .A1(n4757), .A2(n4758), .A3(n4759), .A4(n4760), .ZN(n4747) );
  OAI221_X1 U329 ( .B1(n5201), .B2(n4565), .C1(n5202), .C2(n4566), .A(n4761), 
        .ZN(n4760) );
  AOI22_X1 U330 ( .A1(n4568), .A2(n2822), .B1(n4569), .B2(n2758), .ZN(n4761)
         );
  OAI221_X1 U331 ( .B1(n5585), .B2(n4570), .C1(n5200), .C2(n4571), .A(n4762), 
        .ZN(n4759) );
  AOI22_X1 U332 ( .A1(n4573), .A2(n3046), .B1(n4574), .B2(n3270), .ZN(n4762)
         );
  OAI221_X1 U333 ( .B1(n5649), .B2(n4575), .C1(n5457), .C2(n4576), .A(n4763), 
        .ZN(n4758) );
  AOI22_X1 U334 ( .A1(n4578), .A2(n3526), .B1(n4579), .B2(n3334), .ZN(n4763)
         );
  OAI221_X1 U335 ( .B1(n5199), .B2(n4580), .C1(n5329), .C2(n4581), .A(n4764), 
        .ZN(n4757) );
  AOI22_X1 U336 ( .A1(n4583), .A2(n3206), .B1(n4584), .B2(n3430), .ZN(n4764)
         );
  NAND2_X1 U337 ( .A1(n4765), .A2(n4766), .ZN(N399) );
  NOR4_X1 U338 ( .A1(n4767), .A2(n4768), .A3(n4769), .A4(n4770), .ZN(n4766) );
  OAI221_X1 U339 ( .B1(n5362), .B2(n4541), .C1(n5490), .C2(n4542), .A(n4771), 
        .ZN(n4770) );
  AOI22_X1 U340 ( .A1(n4544), .A2(n3397), .B1(n4545), .B2(n3173), .ZN(n4771)
         );
  OAI221_X1 U341 ( .B1(n5426), .B2(n4546), .C1(n5618), .C2(n4547), .A(n4772), 
        .ZN(n4769) );
  AOI22_X1 U342 ( .A1(n4549), .A2(n3141), .B1(n4550), .B2(n2949), .ZN(n4772)
         );
  OAI221_X1 U343 ( .B1(n5394), .B2(n4551), .C1(n5522), .C2(n4552), .A(n4773), 
        .ZN(n4768) );
  AOI22_X1 U344 ( .A1(n4554), .A2(n3109), .B1(n4555), .B2(n2853), .ZN(n4773)
         );
  OAI221_X1 U345 ( .B1(n5554), .B2(n4556), .C1(n5298), .C2(n4557), .A(n4774), 
        .ZN(n4767) );
  AOI22_X1 U346 ( .A1(n4559), .A2(n3493), .B1(n4560), .B2(n2981), .ZN(n4774)
         );
  NOR4_X1 U347 ( .A1(n4775), .A2(n4776), .A3(n4777), .A4(n4778), .ZN(n4765) );
  OAI221_X1 U348 ( .B1(n5205), .B2(n4565), .C1(n5206), .C2(n4566), .A(n4779), 
        .ZN(n4778) );
  AOI22_X1 U349 ( .A1(n4568), .A2(n2821), .B1(n4569), .B2(n2757), .ZN(n4779)
         );
  OAI221_X1 U350 ( .B1(n5586), .B2(n4570), .C1(n5204), .C2(n4571), .A(n4780), 
        .ZN(n4777) );
  AOI22_X1 U351 ( .A1(n4573), .A2(n3045), .B1(n4574), .B2(n3269), .ZN(n4780)
         );
  OAI221_X1 U352 ( .B1(n5650), .B2(n4575), .C1(n5458), .C2(n4576), .A(n4781), 
        .ZN(n4776) );
  AOI22_X1 U353 ( .A1(n4578), .A2(n3525), .B1(n4579), .B2(n3333), .ZN(n4781)
         );
  OAI221_X1 U354 ( .B1(n5203), .B2(n4580), .C1(n5330), .C2(n4581), .A(n4782), 
        .ZN(n4775) );
  AOI22_X1 U355 ( .A1(n4583), .A2(n3205), .B1(n4584), .B2(n3429), .ZN(n4782)
         );
  NAND2_X1 U356 ( .A1(n4783), .A2(n4784), .ZN(N398) );
  NOR4_X1 U357 ( .A1(n4785), .A2(n4786), .A3(n4787), .A4(n4788), .ZN(n4784) );
  OAI221_X1 U358 ( .B1(n5363), .B2(n4541), .C1(n5491), .C2(n4542), .A(n4789), 
        .ZN(n4788) );
  AOI22_X1 U359 ( .A1(n4544), .A2(n3396), .B1(n4545), .B2(n3172), .ZN(n4789)
         );
  OAI221_X1 U360 ( .B1(n5427), .B2(n4546), .C1(n5619), .C2(n4547), .A(n4790), 
        .ZN(n4787) );
  AOI22_X1 U361 ( .A1(n4549), .A2(n3140), .B1(n4550), .B2(n2948), .ZN(n4790)
         );
  OAI221_X1 U362 ( .B1(n5395), .B2(n4551), .C1(n5523), .C2(n4552), .A(n4791), 
        .ZN(n4786) );
  AOI22_X1 U363 ( .A1(n4554), .A2(n3108), .B1(n4555), .B2(n2852), .ZN(n4791)
         );
  OAI221_X1 U364 ( .B1(n5555), .B2(n4556), .C1(n5299), .C2(n4557), .A(n4792), 
        .ZN(n4785) );
  AOI22_X1 U365 ( .A1(n4559), .A2(n3492), .B1(n4560), .B2(n2980), .ZN(n4792)
         );
  NOR4_X1 U366 ( .A1(n4793), .A2(n4794), .A3(n4795), .A4(n4796), .ZN(n4783) );
  OAI221_X1 U367 ( .B1(n5209), .B2(n4565), .C1(n5210), .C2(n4566), .A(n4797), 
        .ZN(n4796) );
  AOI22_X1 U368 ( .A1(n4568), .A2(n2820), .B1(n4569), .B2(n2756), .ZN(n4797)
         );
  OAI221_X1 U369 ( .B1(n5587), .B2(n4570), .C1(n5208), .C2(n4571), .A(n4798), 
        .ZN(n4795) );
  AOI22_X1 U370 ( .A1(n4573), .A2(n3044), .B1(n4574), .B2(n3268), .ZN(n4798)
         );
  OAI221_X1 U371 ( .B1(n5651), .B2(n4575), .C1(n5459), .C2(n4576), .A(n4799), 
        .ZN(n4794) );
  AOI22_X1 U372 ( .A1(n4578), .A2(n3524), .B1(n4579), .B2(n3332), .ZN(n4799)
         );
  OAI221_X1 U373 ( .B1(n5207), .B2(n4580), .C1(n5331), .C2(n4581), .A(n4800), 
        .ZN(n4793) );
  AOI22_X1 U374 ( .A1(n4583), .A2(n3204), .B1(n4584), .B2(n3428), .ZN(n4800)
         );
  NAND2_X1 U375 ( .A1(n4801), .A2(n4802), .ZN(N397) );
  NOR4_X1 U376 ( .A1(n4803), .A2(n4804), .A3(n4805), .A4(n4806), .ZN(n4802) );
  OAI221_X1 U377 ( .B1(n5364), .B2(n4541), .C1(n5492), .C2(n4542), .A(n4807), 
        .ZN(n4806) );
  AOI22_X1 U378 ( .A1(n4544), .A2(n3395), .B1(n4545), .B2(n3171), .ZN(n4807)
         );
  OAI221_X1 U379 ( .B1(n5428), .B2(n4546), .C1(n5620), .C2(n4547), .A(n4808), 
        .ZN(n4805) );
  AOI22_X1 U380 ( .A1(n4549), .A2(n3139), .B1(n4550), .B2(n2947), .ZN(n4808)
         );
  OAI221_X1 U381 ( .B1(n5396), .B2(n4551), .C1(n5524), .C2(n4552), .A(n4809), 
        .ZN(n4804) );
  AOI22_X1 U382 ( .A1(n4554), .A2(n3107), .B1(n4555), .B2(n2851), .ZN(n4809)
         );
  OAI221_X1 U383 ( .B1(n5556), .B2(n4556), .C1(n5300), .C2(n4557), .A(n4810), 
        .ZN(n4803) );
  AOI22_X1 U384 ( .A1(n4559), .A2(n3491), .B1(n4560), .B2(n2979), .ZN(n4810)
         );
  NOR4_X1 U385 ( .A1(n4811), .A2(n4812), .A3(n4813), .A4(n4814), .ZN(n4801) );
  OAI221_X1 U386 ( .B1(n5213), .B2(n4565), .C1(n5214), .C2(n4566), .A(n4815), 
        .ZN(n4814) );
  AOI22_X1 U387 ( .A1(n4568), .A2(n2819), .B1(n4569), .B2(n2755), .ZN(n4815)
         );
  OAI221_X1 U388 ( .B1(n5588), .B2(n4570), .C1(n5212), .C2(n4571), .A(n4816), 
        .ZN(n4813) );
  AOI22_X1 U389 ( .A1(n4573), .A2(n3043), .B1(n4574), .B2(n3267), .ZN(n4816)
         );
  OAI221_X1 U390 ( .B1(n5652), .B2(n4575), .C1(n5460), .C2(n4576), .A(n4817), 
        .ZN(n4812) );
  AOI22_X1 U391 ( .A1(n4578), .A2(n3523), .B1(n4579), .B2(n3331), .ZN(n4817)
         );
  OAI221_X1 U392 ( .B1(n5211), .B2(n4580), .C1(n5332), .C2(n4581), .A(n4818), 
        .ZN(n4811) );
  AOI22_X1 U393 ( .A1(n4583), .A2(n3203), .B1(n4584), .B2(n3427), .ZN(n4818)
         );
  NAND2_X1 U394 ( .A1(n4819), .A2(n4820), .ZN(N396) );
  NOR4_X1 U395 ( .A1(n4821), .A2(n4822), .A3(n4823), .A4(n4824), .ZN(n4820) );
  OAI221_X1 U396 ( .B1(n5365), .B2(n4541), .C1(n5493), .C2(n4542), .A(n4825), 
        .ZN(n4824) );
  AOI22_X1 U397 ( .A1(n4544), .A2(n3394), .B1(n4545), .B2(n3170), .ZN(n4825)
         );
  OAI221_X1 U398 ( .B1(n5429), .B2(n4546), .C1(n5621), .C2(n4547), .A(n4826), 
        .ZN(n4823) );
  AOI22_X1 U399 ( .A1(n4549), .A2(n3138), .B1(n4550), .B2(n2946), .ZN(n4826)
         );
  OAI221_X1 U400 ( .B1(n5397), .B2(n4551), .C1(n5525), .C2(n4552), .A(n4827), 
        .ZN(n4822) );
  AOI22_X1 U401 ( .A1(n4554), .A2(n3106), .B1(n4555), .B2(n2850), .ZN(n4827)
         );
  OAI221_X1 U402 ( .B1(n5557), .B2(n4556), .C1(n5301), .C2(n4557), .A(n4828), 
        .ZN(n4821) );
  AOI22_X1 U403 ( .A1(n4559), .A2(n3490), .B1(n4560), .B2(n2978), .ZN(n4828)
         );
  NOR4_X1 U404 ( .A1(n4829), .A2(n4830), .A3(n4831), .A4(n4832), .ZN(n4819) );
  OAI221_X1 U405 ( .B1(n5217), .B2(n4565), .C1(n5218), .C2(n4566), .A(n4833), 
        .ZN(n4832) );
  AOI22_X1 U406 ( .A1(n4568), .A2(n2818), .B1(n4569), .B2(n2754), .ZN(n4833)
         );
  OAI221_X1 U407 ( .B1(n5589), .B2(n4570), .C1(n5216), .C2(n4571), .A(n4834), 
        .ZN(n4831) );
  AOI22_X1 U408 ( .A1(n4573), .A2(n3042), .B1(n4574), .B2(n3266), .ZN(n4834)
         );
  OAI221_X1 U409 ( .B1(n5653), .B2(n4575), .C1(n5461), .C2(n4576), .A(n4835), 
        .ZN(n4830) );
  AOI22_X1 U410 ( .A1(n4578), .A2(n3522), .B1(n4579), .B2(n3330), .ZN(n4835)
         );
  OAI221_X1 U411 ( .B1(n5215), .B2(n4580), .C1(n5333), .C2(n4581), .A(n4836), 
        .ZN(n4829) );
  AOI22_X1 U412 ( .A1(n4583), .A2(n3202), .B1(n4584), .B2(n3426), .ZN(n4836)
         );
  NAND2_X1 U413 ( .A1(n4837), .A2(n4838), .ZN(N395) );
  NOR4_X1 U414 ( .A1(n4839), .A2(n4840), .A3(n4841), .A4(n4842), .ZN(n4838) );
  OAI221_X1 U415 ( .B1(n5366), .B2(n4541), .C1(n5494), .C2(n4542), .A(n4843), 
        .ZN(n4842) );
  AOI22_X1 U416 ( .A1(n4544), .A2(n3393), .B1(n4545), .B2(n3169), .ZN(n4843)
         );
  OAI221_X1 U417 ( .B1(n5430), .B2(n4546), .C1(n5622), .C2(n4547), .A(n4844), 
        .ZN(n4841) );
  AOI22_X1 U418 ( .A1(n4549), .A2(n3137), .B1(n4550), .B2(n2945), .ZN(n4844)
         );
  OAI221_X1 U419 ( .B1(n5398), .B2(n4551), .C1(n5526), .C2(n4552), .A(n4845), 
        .ZN(n4840) );
  AOI22_X1 U420 ( .A1(n4554), .A2(n3105), .B1(n4555), .B2(n2849), .ZN(n4845)
         );
  OAI221_X1 U421 ( .B1(n5558), .B2(n4556), .C1(n5302), .C2(n4557), .A(n4846), 
        .ZN(n4839) );
  AOI22_X1 U422 ( .A1(n4559), .A2(n3489), .B1(n4560), .B2(n2977), .ZN(n4846)
         );
  NOR4_X1 U423 ( .A1(n4847), .A2(n4848), .A3(n4849), .A4(n4850), .ZN(n4837) );
  OAI221_X1 U424 ( .B1(n5221), .B2(n4565), .C1(n5222), .C2(n4566), .A(n4851), 
        .ZN(n4850) );
  AOI22_X1 U425 ( .A1(n4568), .A2(n2817), .B1(n4569), .B2(n2753), .ZN(n4851)
         );
  OAI221_X1 U426 ( .B1(n5590), .B2(n4570), .C1(n5220), .C2(n4571), .A(n4852), 
        .ZN(n4849) );
  AOI22_X1 U427 ( .A1(n4573), .A2(n3041), .B1(n4574), .B2(n3265), .ZN(n4852)
         );
  OAI221_X1 U428 ( .B1(n5654), .B2(n4575), .C1(n5462), .C2(n4576), .A(n4853), 
        .ZN(n4848) );
  AOI22_X1 U429 ( .A1(n4578), .A2(n3521), .B1(n4579), .B2(n3329), .ZN(n4853)
         );
  OAI221_X1 U430 ( .B1(n5219), .B2(n4580), .C1(n5334), .C2(n4581), .A(n4854), 
        .ZN(n4847) );
  AOI22_X1 U431 ( .A1(n4583), .A2(n3201), .B1(n4584), .B2(n3425), .ZN(n4854)
         );
  NAND2_X1 U432 ( .A1(n4855), .A2(n4856), .ZN(N394) );
  NOR4_X1 U433 ( .A1(n4857), .A2(n4858), .A3(n4859), .A4(n4860), .ZN(n4856) );
  OAI221_X1 U434 ( .B1(n5367), .B2(n4541), .C1(n5495), .C2(n4542), .A(n4861), 
        .ZN(n4860) );
  AOI22_X1 U435 ( .A1(n4544), .A2(n3392), .B1(n4545), .B2(n3168), .ZN(n4861)
         );
  OAI221_X1 U436 ( .B1(n5431), .B2(n4546), .C1(n5623), .C2(n4547), .A(n4862), 
        .ZN(n4859) );
  AOI22_X1 U437 ( .A1(n4549), .A2(n3136), .B1(n4550), .B2(n2944), .ZN(n4862)
         );
  OAI221_X1 U438 ( .B1(n5399), .B2(n4551), .C1(n5527), .C2(n4552), .A(n4863), 
        .ZN(n4858) );
  AOI22_X1 U439 ( .A1(n4554), .A2(n3104), .B1(n4555), .B2(n2848), .ZN(n4863)
         );
  OAI221_X1 U440 ( .B1(n5559), .B2(n4556), .C1(n5303), .C2(n4557), .A(n4864), 
        .ZN(n4857) );
  AOI22_X1 U441 ( .A1(n4559), .A2(n3488), .B1(n4560), .B2(n2976), .ZN(n4864)
         );
  NOR4_X1 U442 ( .A1(n4865), .A2(n4866), .A3(n4867), .A4(n4868), .ZN(n4855) );
  OAI221_X1 U443 ( .B1(n5225), .B2(n4565), .C1(n5226), .C2(n4566), .A(n4869), 
        .ZN(n4868) );
  AOI22_X1 U444 ( .A1(n4568), .A2(n2816), .B1(n4569), .B2(n2752), .ZN(n4869)
         );
  OAI221_X1 U445 ( .B1(n5591), .B2(n4570), .C1(n5224), .C2(n4571), .A(n4870), 
        .ZN(n4867) );
  AOI22_X1 U446 ( .A1(n4573), .A2(n3040), .B1(n4574), .B2(n3264), .ZN(n4870)
         );
  OAI221_X1 U447 ( .B1(n5655), .B2(n4575), .C1(n5463), .C2(n4576), .A(n4871), 
        .ZN(n4866) );
  AOI22_X1 U448 ( .A1(n4578), .A2(n3520), .B1(n4579), .B2(n3328), .ZN(n4871)
         );
  OAI221_X1 U449 ( .B1(n5223), .B2(n4580), .C1(n5335), .C2(n4581), .A(n4872), 
        .ZN(n4865) );
  AOI22_X1 U450 ( .A1(n4583), .A2(n3200), .B1(n4584), .B2(n3424), .ZN(n4872)
         );
  NAND2_X1 U451 ( .A1(n4873), .A2(n4874), .ZN(N393) );
  NOR4_X1 U452 ( .A1(n4875), .A2(n4876), .A3(n4877), .A4(n4878), .ZN(n4874) );
  OAI221_X1 U453 ( .B1(n5368), .B2(n4541), .C1(n5496), .C2(n4542), .A(n4879), 
        .ZN(n4878) );
  AOI22_X1 U454 ( .A1(n4544), .A2(n3391), .B1(n4545), .B2(n3167), .ZN(n4879)
         );
  OAI221_X1 U455 ( .B1(n5432), .B2(n4546), .C1(n5624), .C2(n4547), .A(n4880), 
        .ZN(n4877) );
  AOI22_X1 U456 ( .A1(n4549), .A2(n3135), .B1(n4550), .B2(n2943), .ZN(n4880)
         );
  OAI221_X1 U457 ( .B1(n5400), .B2(n4551), .C1(n5528), .C2(n4552), .A(n4881), 
        .ZN(n4876) );
  AOI22_X1 U458 ( .A1(n4554), .A2(n3103), .B1(n4555), .B2(n2847), .ZN(n4881)
         );
  OAI221_X1 U459 ( .B1(n5560), .B2(n4556), .C1(n5304), .C2(n4557), .A(n4882), 
        .ZN(n4875) );
  AOI22_X1 U460 ( .A1(n4559), .A2(n3487), .B1(n4560), .B2(n2975), .ZN(n4882)
         );
  NOR4_X1 U461 ( .A1(n4883), .A2(n4884), .A3(n4885), .A4(n4886), .ZN(n4873) );
  OAI221_X1 U462 ( .B1(n5229), .B2(n4565), .C1(n5230), .C2(n4566), .A(n4887), 
        .ZN(n4886) );
  AOI22_X1 U463 ( .A1(n4568), .A2(n2815), .B1(n4569), .B2(n2751), .ZN(n4887)
         );
  OAI221_X1 U464 ( .B1(n5592), .B2(n4570), .C1(n5228), .C2(n4571), .A(n4888), 
        .ZN(n4885) );
  AOI22_X1 U465 ( .A1(n4573), .A2(n3039), .B1(n4574), .B2(n3263), .ZN(n4888)
         );
  OAI221_X1 U466 ( .B1(n5656), .B2(n4575), .C1(n5464), .C2(n4576), .A(n4889), 
        .ZN(n4884) );
  AOI22_X1 U467 ( .A1(n4578), .A2(n3519), .B1(n4579), .B2(n3327), .ZN(n4889)
         );
  OAI221_X1 U468 ( .B1(n5227), .B2(n4580), .C1(n5336), .C2(n4581), .A(n4890), 
        .ZN(n4883) );
  AOI22_X1 U469 ( .A1(n4583), .A2(n3199), .B1(n4584), .B2(n3423), .ZN(n4890)
         );
  NAND2_X1 U470 ( .A1(n4891), .A2(n4892), .ZN(N392) );
  NOR4_X1 U471 ( .A1(n4893), .A2(n4894), .A3(n4895), .A4(n4896), .ZN(n4892) );
  OAI221_X1 U472 ( .B1(n5369), .B2(n4541), .C1(n5497), .C2(n4542), .A(n4897), 
        .ZN(n4896) );
  AOI22_X1 U473 ( .A1(n4544), .A2(n3390), .B1(n4545), .B2(n3166), .ZN(n4897)
         );
  OAI221_X1 U474 ( .B1(n5433), .B2(n4546), .C1(n5625), .C2(n4547), .A(n4898), 
        .ZN(n4895) );
  AOI22_X1 U475 ( .A1(n4549), .A2(n3134), .B1(n4550), .B2(n2942), .ZN(n4898)
         );
  OAI221_X1 U476 ( .B1(n5401), .B2(n4551), .C1(n5529), .C2(n4552), .A(n4899), 
        .ZN(n4894) );
  AOI22_X1 U477 ( .A1(n4554), .A2(n3102), .B1(n4555), .B2(n2846), .ZN(n4899)
         );
  OAI221_X1 U478 ( .B1(n5561), .B2(n4556), .C1(n5305), .C2(n4557), .A(n4900), 
        .ZN(n4893) );
  AOI22_X1 U479 ( .A1(n4559), .A2(n3486), .B1(n4560), .B2(n2974), .ZN(n4900)
         );
  NOR4_X1 U480 ( .A1(n4901), .A2(n4902), .A3(n4903), .A4(n4904), .ZN(n4891) );
  OAI221_X1 U481 ( .B1(n5233), .B2(n4565), .C1(n5234), .C2(n4566), .A(n4905), 
        .ZN(n4904) );
  AOI22_X1 U482 ( .A1(n4568), .A2(n2814), .B1(n4569), .B2(n2750), .ZN(n4905)
         );
  OAI221_X1 U483 ( .B1(n5593), .B2(n4570), .C1(n5232), .C2(n4571), .A(n4906), 
        .ZN(n4903) );
  AOI22_X1 U484 ( .A1(n4573), .A2(n3038), .B1(n4574), .B2(n3262), .ZN(n4906)
         );
  OAI221_X1 U485 ( .B1(n5657), .B2(n4575), .C1(n5465), .C2(n4576), .A(n4907), 
        .ZN(n4902) );
  AOI22_X1 U486 ( .A1(n4578), .A2(n3518), .B1(n4579), .B2(n3326), .ZN(n4907)
         );
  OAI221_X1 U487 ( .B1(n5231), .B2(n4580), .C1(n5337), .C2(n4581), .A(n4908), 
        .ZN(n4901) );
  AOI22_X1 U488 ( .A1(n4583), .A2(n3198), .B1(n4584), .B2(n3422), .ZN(n4908)
         );
  NAND2_X1 U489 ( .A1(n4909), .A2(n4910), .ZN(N391) );
  NOR4_X1 U490 ( .A1(n4911), .A2(n4912), .A3(n4913), .A4(n4914), .ZN(n4910) );
  OAI221_X1 U491 ( .B1(n5370), .B2(n4541), .C1(n5498), .C2(n4542), .A(n4915), 
        .ZN(n4914) );
  AOI22_X1 U492 ( .A1(n4544), .A2(n3389), .B1(n4545), .B2(n3165), .ZN(n4915)
         );
  OAI221_X1 U493 ( .B1(n5434), .B2(n4546), .C1(n5626), .C2(n4547), .A(n4916), 
        .ZN(n4913) );
  AOI22_X1 U494 ( .A1(n4549), .A2(n3133), .B1(n4550), .B2(n2941), .ZN(n4916)
         );
  OAI221_X1 U495 ( .B1(n5402), .B2(n4551), .C1(n5530), .C2(n4552), .A(n4917), 
        .ZN(n4912) );
  AOI22_X1 U496 ( .A1(n4554), .A2(n3101), .B1(n4555), .B2(n2845), .ZN(n4917)
         );
  OAI221_X1 U497 ( .B1(n5562), .B2(n4556), .C1(n5306), .C2(n4557), .A(n4918), 
        .ZN(n4911) );
  AOI22_X1 U498 ( .A1(n4559), .A2(n3485), .B1(n4560), .B2(n2973), .ZN(n4918)
         );
  NOR4_X1 U499 ( .A1(n4919), .A2(n4920), .A3(n4921), .A4(n4922), .ZN(n4909) );
  OAI221_X1 U500 ( .B1(n5237), .B2(n4565), .C1(n5238), .C2(n4566), .A(n4923), 
        .ZN(n4922) );
  AOI22_X1 U501 ( .A1(n4568), .A2(n2813), .B1(n4569), .B2(n2749), .ZN(n4923)
         );
  OAI221_X1 U502 ( .B1(n5594), .B2(n4570), .C1(n5236), .C2(n4571), .A(n4924), 
        .ZN(n4921) );
  AOI22_X1 U503 ( .A1(n4573), .A2(n3037), .B1(n4574), .B2(n3261), .ZN(n4924)
         );
  OAI221_X1 U504 ( .B1(n5658), .B2(n4575), .C1(n5466), .C2(n4576), .A(n4925), 
        .ZN(n4920) );
  AOI22_X1 U505 ( .A1(n4578), .A2(n3517), .B1(n4579), .B2(n3325), .ZN(n4925)
         );
  OAI221_X1 U506 ( .B1(n5235), .B2(n4580), .C1(n5338), .C2(n4581), .A(n4926), 
        .ZN(n4919) );
  AOI22_X1 U507 ( .A1(n4583), .A2(n3197), .B1(n4584), .B2(n3421), .ZN(n4926)
         );
  NAND2_X1 U508 ( .A1(n4927), .A2(n4928), .ZN(N390) );
  NOR4_X1 U509 ( .A1(n4929), .A2(n4930), .A3(n4931), .A4(n4932), .ZN(n4928) );
  OAI221_X1 U510 ( .B1(n5371), .B2(n4541), .C1(n5499), .C2(n4542), .A(n4933), 
        .ZN(n4932) );
  AOI22_X1 U511 ( .A1(n4544), .A2(n3388), .B1(n4545), .B2(n3164), .ZN(n4933)
         );
  OAI221_X1 U512 ( .B1(n5435), .B2(n4546), .C1(n5627), .C2(n4547), .A(n4934), 
        .ZN(n4931) );
  AOI22_X1 U513 ( .A1(n4549), .A2(n3132), .B1(n4550), .B2(n2940), .ZN(n4934)
         );
  OAI221_X1 U514 ( .B1(n5403), .B2(n4551), .C1(n5531), .C2(n4552), .A(n4935), 
        .ZN(n4930) );
  AOI22_X1 U515 ( .A1(n4554), .A2(n3100), .B1(n4555), .B2(n2844), .ZN(n4935)
         );
  OAI221_X1 U516 ( .B1(n5563), .B2(n4556), .C1(n5307), .C2(n4557), .A(n4936), 
        .ZN(n4929) );
  AOI22_X1 U517 ( .A1(n4559), .A2(n3484), .B1(n4560), .B2(n2972), .ZN(n4936)
         );
  NOR4_X1 U518 ( .A1(n4937), .A2(n4938), .A3(n4939), .A4(n4940), .ZN(n4927) );
  OAI221_X1 U519 ( .B1(n5241), .B2(n4565), .C1(n5242), .C2(n4566), .A(n4941), 
        .ZN(n4940) );
  AOI22_X1 U520 ( .A1(n4568), .A2(n2812), .B1(n4569), .B2(n2748), .ZN(n4941)
         );
  OAI221_X1 U521 ( .B1(n5595), .B2(n4570), .C1(n5240), .C2(n4571), .A(n4942), 
        .ZN(n4939) );
  AOI22_X1 U522 ( .A1(n4573), .A2(n3036), .B1(n4574), .B2(n3260), .ZN(n4942)
         );
  OAI221_X1 U523 ( .B1(n5659), .B2(n4575), .C1(n5467), .C2(n4576), .A(n4943), 
        .ZN(n4938) );
  AOI22_X1 U524 ( .A1(n4578), .A2(n3516), .B1(n4579), .B2(n3324), .ZN(n4943)
         );
  OAI221_X1 U525 ( .B1(n5239), .B2(n4580), .C1(n5339), .C2(n4581), .A(n4944), 
        .ZN(n4937) );
  AOI22_X1 U526 ( .A1(n4583), .A2(n3196), .B1(n4584), .B2(n3420), .ZN(n4944)
         );
  NAND2_X1 U527 ( .A1(n4945), .A2(n4946), .ZN(N389) );
  NOR4_X1 U528 ( .A1(n4947), .A2(n4948), .A3(n4949), .A4(n4950), .ZN(n4946) );
  OAI221_X1 U529 ( .B1(n5372), .B2(n4541), .C1(n5500), .C2(n4542), .A(n4951), 
        .ZN(n4950) );
  AOI22_X1 U530 ( .A1(n4544), .A2(n3387), .B1(n4545), .B2(n3163), .ZN(n4951)
         );
  OAI221_X1 U531 ( .B1(n5436), .B2(n4546), .C1(n5628), .C2(n4547), .A(n4952), 
        .ZN(n4949) );
  AOI22_X1 U532 ( .A1(n4549), .A2(n3131), .B1(n4550), .B2(n2939), .ZN(n4952)
         );
  OAI221_X1 U533 ( .B1(n5404), .B2(n4551), .C1(n5532), .C2(n4552), .A(n4953), 
        .ZN(n4948) );
  AOI22_X1 U534 ( .A1(n4554), .A2(n3099), .B1(n4555), .B2(n2843), .ZN(n4953)
         );
  OAI221_X1 U535 ( .B1(n5564), .B2(n4556), .C1(n5308), .C2(n4557), .A(n4954), 
        .ZN(n4947) );
  AOI22_X1 U536 ( .A1(n4559), .A2(n3483), .B1(n4560), .B2(n2971), .ZN(n4954)
         );
  NOR4_X1 U537 ( .A1(n4955), .A2(n4956), .A3(n4957), .A4(n4958), .ZN(n4945) );
  OAI221_X1 U538 ( .B1(n5245), .B2(n4565), .C1(n5246), .C2(n4566), .A(n4959), 
        .ZN(n4958) );
  AOI22_X1 U539 ( .A1(n4568), .A2(n2811), .B1(n4569), .B2(n2747), .ZN(n4959)
         );
  OAI221_X1 U540 ( .B1(n5596), .B2(n4570), .C1(n5244), .C2(n4571), .A(n4960), 
        .ZN(n4957) );
  AOI22_X1 U541 ( .A1(n4573), .A2(n3035), .B1(n4574), .B2(n3259), .ZN(n4960)
         );
  OAI221_X1 U542 ( .B1(n5660), .B2(n4575), .C1(n5468), .C2(n4576), .A(n4961), 
        .ZN(n4956) );
  AOI22_X1 U543 ( .A1(n4578), .A2(n3515), .B1(n4579), .B2(n3323), .ZN(n4961)
         );
  OAI221_X1 U544 ( .B1(n5243), .B2(n4580), .C1(n5340), .C2(n4581), .A(n4962), 
        .ZN(n4955) );
  AOI22_X1 U545 ( .A1(n4583), .A2(n3195), .B1(n4584), .B2(n3419), .ZN(n4962)
         );
  NAND2_X1 U546 ( .A1(n4963), .A2(n4964), .ZN(N388) );
  NOR4_X1 U547 ( .A1(n4965), .A2(n4966), .A3(n4967), .A4(n4968), .ZN(n4964) );
  OAI221_X1 U548 ( .B1(n5373), .B2(n4541), .C1(n5501), .C2(n4542), .A(n4969), 
        .ZN(n4968) );
  AOI22_X1 U549 ( .A1(n4544), .A2(n3386), .B1(n4545), .B2(n3162), .ZN(n4969)
         );
  OAI221_X1 U550 ( .B1(n5437), .B2(n4546), .C1(n5629), .C2(n4547), .A(n4970), 
        .ZN(n4967) );
  AOI22_X1 U551 ( .A1(n4549), .A2(n3130), .B1(n4550), .B2(n2938), .ZN(n4970)
         );
  OAI221_X1 U552 ( .B1(n5405), .B2(n4551), .C1(n5533), .C2(n4552), .A(n4971), 
        .ZN(n4966) );
  AOI22_X1 U553 ( .A1(n4554), .A2(n3098), .B1(n4555), .B2(n2842), .ZN(n4971)
         );
  OAI221_X1 U554 ( .B1(n5565), .B2(n4556), .C1(n5309), .C2(n4557), .A(n4972), 
        .ZN(n4965) );
  AOI22_X1 U555 ( .A1(n4559), .A2(n3482), .B1(n4560), .B2(n2970), .ZN(n4972)
         );
  NOR4_X1 U556 ( .A1(n4973), .A2(n4974), .A3(n4975), .A4(n4976), .ZN(n4963) );
  OAI221_X1 U557 ( .B1(n5249), .B2(n4565), .C1(n5250), .C2(n4566), .A(n4977), 
        .ZN(n4976) );
  AOI22_X1 U558 ( .A1(n4568), .A2(n2810), .B1(n4569), .B2(n2746), .ZN(n4977)
         );
  OAI221_X1 U559 ( .B1(n5597), .B2(n4570), .C1(n5248), .C2(n4571), .A(n4978), 
        .ZN(n4975) );
  AOI22_X1 U560 ( .A1(n4573), .A2(n3034), .B1(n4574), .B2(n3258), .ZN(n4978)
         );
  OAI221_X1 U561 ( .B1(n5661), .B2(n4575), .C1(n5469), .C2(n4576), .A(n4979), 
        .ZN(n4974) );
  AOI22_X1 U562 ( .A1(n4578), .A2(n3514), .B1(n4579), .B2(n3322), .ZN(n4979)
         );
  OAI221_X1 U563 ( .B1(n5247), .B2(n4580), .C1(n5341), .C2(n4581), .A(n4980), 
        .ZN(n4973) );
  AOI22_X1 U564 ( .A1(n4583), .A2(n3194), .B1(n4584), .B2(n3418), .ZN(n4980)
         );
  NAND2_X1 U565 ( .A1(n4981), .A2(n4982), .ZN(N387) );
  NOR4_X1 U566 ( .A1(n4983), .A2(n4984), .A3(n4985), .A4(n4986), .ZN(n4982) );
  OAI221_X1 U567 ( .B1(n5374), .B2(n4541), .C1(n5502), .C2(n4542), .A(n4987), 
        .ZN(n4986) );
  AOI22_X1 U568 ( .A1(n4544), .A2(n3385), .B1(n4545), .B2(n3161), .ZN(n4987)
         );
  OAI221_X1 U569 ( .B1(n5438), .B2(n4546), .C1(n5630), .C2(n4547), .A(n4988), 
        .ZN(n4985) );
  AOI22_X1 U570 ( .A1(n4549), .A2(n3129), .B1(n4550), .B2(n2937), .ZN(n4988)
         );
  OAI221_X1 U571 ( .B1(n5406), .B2(n4551), .C1(n5534), .C2(n4552), .A(n4989), 
        .ZN(n4984) );
  AOI22_X1 U572 ( .A1(n4554), .A2(n3097), .B1(n4555), .B2(n2841), .ZN(n4989)
         );
  OAI221_X1 U573 ( .B1(n5566), .B2(n4556), .C1(n5310), .C2(n4557), .A(n4990), 
        .ZN(n4983) );
  AOI22_X1 U574 ( .A1(n4559), .A2(n3481), .B1(n4560), .B2(n2969), .ZN(n4990)
         );
  NOR4_X1 U575 ( .A1(n4991), .A2(n4992), .A3(n4993), .A4(n4994), .ZN(n4981) );
  OAI221_X1 U576 ( .B1(n5253), .B2(n4565), .C1(n5254), .C2(n4566), .A(n4995), 
        .ZN(n4994) );
  AOI22_X1 U577 ( .A1(n4568), .A2(n2809), .B1(n4569), .B2(n2745), .ZN(n4995)
         );
  OAI221_X1 U578 ( .B1(n5598), .B2(n4570), .C1(n5252), .C2(n4571), .A(n4996), 
        .ZN(n4993) );
  AOI22_X1 U579 ( .A1(n4573), .A2(n3033), .B1(n4574), .B2(n3257), .ZN(n4996)
         );
  OAI221_X1 U580 ( .B1(n5662), .B2(n4575), .C1(n5470), .C2(n4576), .A(n4997), 
        .ZN(n4992) );
  AOI22_X1 U581 ( .A1(n4578), .A2(n3513), .B1(n4579), .B2(n3321), .ZN(n4997)
         );
  OAI221_X1 U582 ( .B1(n5251), .B2(n4580), .C1(n5342), .C2(n4581), .A(n4998), 
        .ZN(n4991) );
  AOI22_X1 U583 ( .A1(n4583), .A2(n3193), .B1(n4584), .B2(n3417), .ZN(n4998)
         );
  NAND2_X1 U584 ( .A1(n4999), .A2(n5000), .ZN(N386) );
  NOR4_X1 U585 ( .A1(n5001), .A2(n5002), .A3(n5003), .A4(n5004), .ZN(n5000) );
  OAI221_X1 U586 ( .B1(n5375), .B2(n4541), .C1(n5503), .C2(n4542), .A(n5005), 
        .ZN(n5004) );
  AOI22_X1 U587 ( .A1(n4544), .A2(n3384), .B1(n4545), .B2(n3160), .ZN(n5005)
         );
  OAI221_X1 U588 ( .B1(n5439), .B2(n4546), .C1(n5631), .C2(n4547), .A(n5006), 
        .ZN(n5003) );
  AOI22_X1 U589 ( .A1(n4549), .A2(n3128), .B1(n4550), .B2(n2936), .ZN(n5006)
         );
  OAI221_X1 U590 ( .B1(n5407), .B2(n4551), .C1(n5535), .C2(n4552), .A(n5007), 
        .ZN(n5002) );
  AOI22_X1 U591 ( .A1(n4554), .A2(n3096), .B1(n4555), .B2(n2840), .ZN(n5007)
         );
  OAI221_X1 U592 ( .B1(n5567), .B2(n4556), .C1(n5311), .C2(n4557), .A(n5008), 
        .ZN(n5001) );
  AOI22_X1 U593 ( .A1(n4559), .A2(n3480), .B1(n4560), .B2(n2968), .ZN(n5008)
         );
  NOR4_X1 U594 ( .A1(n5009), .A2(n5010), .A3(n5011), .A4(n5012), .ZN(n4999) );
  OAI221_X1 U595 ( .B1(n5257), .B2(n4565), .C1(n5258), .C2(n4566), .A(n5013), 
        .ZN(n5012) );
  AOI22_X1 U596 ( .A1(n4568), .A2(n2808), .B1(n4569), .B2(n2744), .ZN(n5013)
         );
  OAI221_X1 U597 ( .B1(n5599), .B2(n4570), .C1(n5256), .C2(n4571), .A(n5014), 
        .ZN(n5011) );
  AOI22_X1 U598 ( .A1(n4573), .A2(n3032), .B1(n4574), .B2(n3256), .ZN(n5014)
         );
  OAI221_X1 U599 ( .B1(n5663), .B2(n4575), .C1(n5471), .C2(n4576), .A(n5015), 
        .ZN(n5010) );
  AOI22_X1 U600 ( .A1(n4578), .A2(n3512), .B1(n4579), .B2(n3320), .ZN(n5015)
         );
  OAI221_X1 U601 ( .B1(n5255), .B2(n4580), .C1(n5343), .C2(n4581), .A(n5016), 
        .ZN(n5009) );
  AOI22_X1 U602 ( .A1(n4583), .A2(n3192), .B1(n4584), .B2(n3416), .ZN(n5016)
         );
  NAND2_X1 U603 ( .A1(n5017), .A2(n5018), .ZN(N385) );
  NOR4_X1 U604 ( .A1(n5019), .A2(n5020), .A3(n5021), .A4(n5022), .ZN(n5018) );
  OAI221_X1 U605 ( .B1(n5376), .B2(n4541), .C1(n5504), .C2(n4542), .A(n5023), 
        .ZN(n5022) );
  AOI22_X1 U606 ( .A1(n4544), .A2(n3383), .B1(n4545), .B2(n3159), .ZN(n5023)
         );
  OAI221_X1 U607 ( .B1(n5440), .B2(n4546), .C1(n5632), .C2(n4547), .A(n5024), 
        .ZN(n5021) );
  AOI22_X1 U608 ( .A1(n4549), .A2(n3127), .B1(n4550), .B2(n2935), .ZN(n5024)
         );
  OAI221_X1 U609 ( .B1(n5408), .B2(n4551), .C1(n5536), .C2(n4552), .A(n5025), 
        .ZN(n5020) );
  AOI22_X1 U610 ( .A1(n4554), .A2(n3095), .B1(n4555), .B2(n2839), .ZN(n5025)
         );
  OAI221_X1 U611 ( .B1(n5568), .B2(n4556), .C1(n5312), .C2(n4557), .A(n5026), 
        .ZN(n5019) );
  AOI22_X1 U612 ( .A1(n4559), .A2(n3479), .B1(n4560), .B2(n2967), .ZN(n5026)
         );
  NOR4_X1 U613 ( .A1(n5027), .A2(n5028), .A3(n5029), .A4(n5030), .ZN(n5017) );
  OAI221_X1 U614 ( .B1(n5261), .B2(n4565), .C1(n5262), .C2(n4566), .A(n5031), 
        .ZN(n5030) );
  AOI22_X1 U615 ( .A1(n4568), .A2(n2807), .B1(n4569), .B2(n2743), .ZN(n5031)
         );
  OAI221_X1 U616 ( .B1(n5600), .B2(n4570), .C1(n5260), .C2(n4571), .A(n5032), 
        .ZN(n5029) );
  AOI22_X1 U617 ( .A1(n4573), .A2(n3031), .B1(n4574), .B2(n3255), .ZN(n5032)
         );
  OAI221_X1 U618 ( .B1(n5664), .B2(n4575), .C1(n5472), .C2(n4576), .A(n5033), 
        .ZN(n5028) );
  AOI22_X1 U619 ( .A1(n4578), .A2(n3511), .B1(n4579), .B2(n3319), .ZN(n5033)
         );
  OAI221_X1 U620 ( .B1(n5259), .B2(n4580), .C1(n5344), .C2(n4581), .A(n5034), 
        .ZN(n5027) );
  AOI22_X1 U621 ( .A1(n4583), .A2(n3191), .B1(n4584), .B2(n3415), .ZN(n5034)
         );
  NAND2_X1 U622 ( .A1(n5035), .A2(n5036), .ZN(N384) );
  NOR4_X1 U623 ( .A1(n5037), .A2(n5038), .A3(n5039), .A4(n5040), .ZN(n5036) );
  OAI221_X1 U624 ( .B1(n5377), .B2(n4541), .C1(n5505), .C2(n4542), .A(n5041), 
        .ZN(n5040) );
  AOI22_X1 U625 ( .A1(n4544), .A2(n3382), .B1(n4545), .B2(n3158), .ZN(n5041)
         );
  OAI221_X1 U626 ( .B1(n5441), .B2(n4546), .C1(n5633), .C2(n4547), .A(n5042), 
        .ZN(n5039) );
  AOI22_X1 U627 ( .A1(n4549), .A2(n3126), .B1(n4550), .B2(n2934), .ZN(n5042)
         );
  OAI221_X1 U628 ( .B1(n5409), .B2(n4551), .C1(n5537), .C2(n4552), .A(n5043), 
        .ZN(n5038) );
  AOI22_X1 U629 ( .A1(n4554), .A2(n3094), .B1(n4555), .B2(n2838), .ZN(n5043)
         );
  OAI221_X1 U630 ( .B1(n5569), .B2(n4556), .C1(n5313), .C2(n4557), .A(n5044), 
        .ZN(n5037) );
  AOI22_X1 U631 ( .A1(n4559), .A2(n3478), .B1(n4560), .B2(n2966), .ZN(n5044)
         );
  NOR4_X1 U632 ( .A1(n5045), .A2(n5046), .A3(n5047), .A4(n5048), .ZN(n5035) );
  OAI221_X1 U633 ( .B1(n5265), .B2(n4565), .C1(n5266), .C2(n4566), .A(n5049), 
        .ZN(n5048) );
  AOI22_X1 U634 ( .A1(n4568), .A2(n2806), .B1(n4569), .B2(n2742), .ZN(n5049)
         );
  OAI221_X1 U635 ( .B1(n5601), .B2(n4570), .C1(n5264), .C2(n4571), .A(n5050), 
        .ZN(n5047) );
  AOI22_X1 U636 ( .A1(n4573), .A2(n3030), .B1(n4574), .B2(n3254), .ZN(n5050)
         );
  OAI221_X1 U637 ( .B1(n5665), .B2(n4575), .C1(n5473), .C2(n4576), .A(n5051), 
        .ZN(n5046) );
  AOI22_X1 U638 ( .A1(n4578), .A2(n3510), .B1(n4579), .B2(n3318), .ZN(n5051)
         );
  OAI221_X1 U639 ( .B1(n5263), .B2(n4580), .C1(n5345), .C2(n4581), .A(n5052), 
        .ZN(n5045) );
  AOI22_X1 U640 ( .A1(n4583), .A2(n3190), .B1(n4584), .B2(n3414), .ZN(n5052)
         );
  NAND2_X1 U641 ( .A1(n5053), .A2(n5054), .ZN(N383) );
  NOR4_X1 U642 ( .A1(n5055), .A2(n5056), .A3(n5057), .A4(n5058), .ZN(n5054) );
  OAI221_X1 U643 ( .B1(n5378), .B2(n4541), .C1(n5506), .C2(n4542), .A(n5059), 
        .ZN(n5058) );
  AOI22_X1 U644 ( .A1(n4544), .A2(n3381), .B1(n4545), .B2(n3157), .ZN(n5059)
         );
  OAI221_X1 U645 ( .B1(n5442), .B2(n4546), .C1(n5634), .C2(n4547), .A(n5060), 
        .ZN(n5057) );
  AOI22_X1 U646 ( .A1(n4549), .A2(n3125), .B1(n4550), .B2(n2933), .ZN(n5060)
         );
  OAI221_X1 U647 ( .B1(n5410), .B2(n4551), .C1(n5538), .C2(n4552), .A(n5061), 
        .ZN(n5056) );
  AOI22_X1 U648 ( .A1(n4554), .A2(n3093), .B1(n4555), .B2(n2837), .ZN(n5061)
         );
  OAI221_X1 U649 ( .B1(n5570), .B2(n4556), .C1(n5314), .C2(n4557), .A(n5062), 
        .ZN(n5055) );
  AOI22_X1 U650 ( .A1(n4559), .A2(n3477), .B1(n4560), .B2(n2965), .ZN(n5062)
         );
  NOR4_X1 U651 ( .A1(n5063), .A2(n5064), .A3(n5065), .A4(n5066), .ZN(n5053) );
  OAI221_X1 U652 ( .B1(n5269), .B2(n4565), .C1(n5270), .C2(n4566), .A(n5067), 
        .ZN(n5066) );
  AOI22_X1 U653 ( .A1(n4568), .A2(n2805), .B1(n4569), .B2(n2741), .ZN(n5067)
         );
  OAI221_X1 U654 ( .B1(n5602), .B2(n4570), .C1(n5268), .C2(n4571), .A(n5068), 
        .ZN(n5065) );
  AOI22_X1 U655 ( .A1(n4573), .A2(n3029), .B1(n4574), .B2(n3253), .ZN(n5068)
         );
  OAI221_X1 U656 ( .B1(n5666), .B2(n4575), .C1(n5474), .C2(n4576), .A(n5069), 
        .ZN(n5064) );
  AOI22_X1 U657 ( .A1(n4578), .A2(n3509), .B1(n4579), .B2(n3317), .ZN(n5069)
         );
  OAI221_X1 U658 ( .B1(n5267), .B2(n4580), .C1(n5346), .C2(n4581), .A(n5070), 
        .ZN(n5063) );
  AOI22_X1 U659 ( .A1(n4583), .A2(n3189), .B1(n4584), .B2(n3413), .ZN(n5070)
         );
  NAND2_X1 U660 ( .A1(n5071), .A2(n5072), .ZN(N382) );
  NOR4_X1 U661 ( .A1(n5073), .A2(n5074), .A3(n5075), .A4(n5076), .ZN(n5072) );
  OAI221_X1 U662 ( .B1(n5379), .B2(n4541), .C1(n5507), .C2(n4542), .A(n5077), 
        .ZN(n5076) );
  AOI22_X1 U663 ( .A1(n4544), .A2(n3380), .B1(n4545), .B2(n3156), .ZN(n5077)
         );
  OAI221_X1 U664 ( .B1(n5443), .B2(n4546), .C1(n5635), .C2(n4547), .A(n5078), 
        .ZN(n5075) );
  AOI22_X1 U665 ( .A1(n4549), .A2(n3124), .B1(n4550), .B2(n2932), .ZN(n5078)
         );
  OAI221_X1 U666 ( .B1(n5411), .B2(n4551), .C1(n5539), .C2(n4552), .A(n5079), 
        .ZN(n5074) );
  AOI22_X1 U667 ( .A1(n4554), .A2(n3092), .B1(n4555), .B2(n2836), .ZN(n5079)
         );
  OAI221_X1 U668 ( .B1(n5571), .B2(n4556), .C1(n5315), .C2(n4557), .A(n5080), 
        .ZN(n5073) );
  AOI22_X1 U669 ( .A1(n4559), .A2(n3476), .B1(n4560), .B2(n2964), .ZN(n5080)
         );
  NOR4_X1 U670 ( .A1(n5081), .A2(n5082), .A3(n5083), .A4(n5084), .ZN(n5071) );
  OAI221_X1 U671 ( .B1(n5273), .B2(n4565), .C1(n5274), .C2(n4566), .A(n5085), 
        .ZN(n5084) );
  AOI22_X1 U672 ( .A1(n4568), .A2(n2804), .B1(n4569), .B2(n2740), .ZN(n5085)
         );
  OAI221_X1 U673 ( .B1(n5603), .B2(n4570), .C1(n5272), .C2(n4571), .A(n5086), 
        .ZN(n5083) );
  AOI22_X1 U674 ( .A1(n4573), .A2(n3028), .B1(n4574), .B2(n3252), .ZN(n5086)
         );
  OAI221_X1 U675 ( .B1(n5667), .B2(n4575), .C1(n5475), .C2(n4576), .A(n5087), 
        .ZN(n5082) );
  AOI22_X1 U676 ( .A1(n4578), .A2(n3508), .B1(n4579), .B2(n3316), .ZN(n5087)
         );
  OAI221_X1 U677 ( .B1(n5271), .B2(n4580), .C1(n5347), .C2(n4581), .A(n5088), 
        .ZN(n5081) );
  AOI22_X1 U678 ( .A1(n4583), .A2(n3188), .B1(n4584), .B2(n3412), .ZN(n5088)
         );
  NAND2_X1 U679 ( .A1(n5089), .A2(n5090), .ZN(N381) );
  NOR4_X1 U680 ( .A1(n5091), .A2(n5092), .A3(n5093), .A4(n5094), .ZN(n5090) );
  OAI221_X1 U681 ( .B1(n5380), .B2(n4541), .C1(n5508), .C2(n4542), .A(n5095), 
        .ZN(n5094) );
  AOI22_X1 U682 ( .A1(n4544), .A2(n3379), .B1(n4545), .B2(n3155), .ZN(n5095)
         );
  OAI221_X1 U683 ( .B1(n5444), .B2(n4546), .C1(n5636), .C2(n4547), .A(n5096), 
        .ZN(n5093) );
  AOI22_X1 U684 ( .A1(n4549), .A2(n3123), .B1(n4550), .B2(n2931), .ZN(n5096)
         );
  OAI221_X1 U685 ( .B1(n5412), .B2(n4551), .C1(n5540), .C2(n4552), .A(n5097), 
        .ZN(n5092) );
  AOI22_X1 U686 ( .A1(n4554), .A2(n3091), .B1(n4555), .B2(n2835), .ZN(n5097)
         );
  OAI221_X1 U687 ( .B1(n5572), .B2(n4556), .C1(n5316), .C2(n4557), .A(n5098), 
        .ZN(n5091) );
  AOI22_X1 U688 ( .A1(n4559), .A2(n3475), .B1(n4560), .B2(n2963), .ZN(n5098)
         );
  NOR4_X1 U689 ( .A1(n5099), .A2(n5100), .A3(n5101), .A4(n5102), .ZN(n5089) );
  OAI221_X1 U690 ( .B1(n5277), .B2(n4565), .C1(n5278), .C2(n4566), .A(n5103), 
        .ZN(n5102) );
  AOI22_X1 U691 ( .A1(n4568), .A2(n2803), .B1(n4569), .B2(n2739), .ZN(n5103)
         );
  OAI221_X1 U692 ( .B1(n5604), .B2(n4570), .C1(n5276), .C2(n4571), .A(n5104), 
        .ZN(n5101) );
  AOI22_X1 U693 ( .A1(n4573), .A2(n3027), .B1(n4574), .B2(n3251), .ZN(n5104)
         );
  OAI221_X1 U694 ( .B1(n5668), .B2(n4575), .C1(n5476), .C2(n4576), .A(n5105), 
        .ZN(n5100) );
  AOI22_X1 U695 ( .A1(n4578), .A2(n3507), .B1(n4579), .B2(n3315), .ZN(n5105)
         );
  OAI221_X1 U696 ( .B1(n5275), .B2(n4580), .C1(n5348), .C2(n4581), .A(n5106), 
        .ZN(n5099) );
  AOI22_X1 U697 ( .A1(n4583), .A2(n3187), .B1(n4584), .B2(n3411), .ZN(n5106)
         );
  NAND2_X1 U698 ( .A1(n5107), .A2(n5108), .ZN(N380) );
  NOR4_X1 U699 ( .A1(n5109), .A2(n5110), .A3(n5111), .A4(n5112), .ZN(n5108) );
  OAI221_X1 U700 ( .B1(n5381), .B2(n4541), .C1(n5509), .C2(n4542), .A(n5113), 
        .ZN(n5112) );
  AOI22_X1 U701 ( .A1(n4544), .A2(n3378), .B1(n4545), .B2(n3154), .ZN(n5113)
         );
  OAI221_X1 U702 ( .B1(n5445), .B2(n4546), .C1(n5637), .C2(n4547), .A(n5114), 
        .ZN(n5111) );
  AOI22_X1 U703 ( .A1(n4549), .A2(n3122), .B1(n4550), .B2(n2930), .ZN(n5114)
         );
  OAI221_X1 U704 ( .B1(n5413), .B2(n4551), .C1(n5541), .C2(n4552), .A(n5115), 
        .ZN(n5110) );
  AOI22_X1 U705 ( .A1(n4554), .A2(n3090), .B1(n4555), .B2(n2834), .ZN(n5115)
         );
  OAI221_X1 U706 ( .B1(n5573), .B2(n4556), .C1(n5317), .C2(n4557), .A(n5116), 
        .ZN(n5109) );
  AOI22_X1 U707 ( .A1(n4559), .A2(n3474), .B1(n4560), .B2(n2962), .ZN(n5116)
         );
  NOR4_X1 U708 ( .A1(n5117), .A2(n5118), .A3(n5119), .A4(n5120), .ZN(n5107) );
  OAI221_X1 U709 ( .B1(n5281), .B2(n4565), .C1(n5282), .C2(n4566), .A(n5121), 
        .ZN(n5120) );
  AOI22_X1 U710 ( .A1(n4568), .A2(n2802), .B1(n4569), .B2(n2738), .ZN(n5121)
         );
  OAI221_X1 U711 ( .B1(n5605), .B2(n4570), .C1(n5280), .C2(n4571), .A(n5122), 
        .ZN(n5119) );
  AOI22_X1 U712 ( .A1(n4573), .A2(n3026), .B1(n4574), .B2(n3250), .ZN(n5122)
         );
  OAI221_X1 U713 ( .B1(n5669), .B2(n4575), .C1(n5477), .C2(n4576), .A(n5123), 
        .ZN(n5118) );
  AOI22_X1 U714 ( .A1(n4578), .A2(n3506), .B1(n4579), .B2(n3314), .ZN(n5123)
         );
  OAI221_X1 U715 ( .B1(n5279), .B2(n4580), .C1(n5349), .C2(n4581), .A(n5124), 
        .ZN(n5117) );
  AOI22_X1 U716 ( .A1(n4583), .A2(n3186), .B1(n4584), .B2(n3410), .ZN(n5124)
         );
  NAND2_X1 U717 ( .A1(n5125), .A2(n5126), .ZN(N379) );
  NOR4_X1 U718 ( .A1(n5127), .A2(n5128), .A3(n5129), .A4(n5130), .ZN(n5126) );
  OAI221_X1 U719 ( .B1(n5382), .B2(n4541), .C1(n5510), .C2(n4542), .A(n5131), 
        .ZN(n5130) );
  AOI22_X1 U720 ( .A1(n4544), .A2(n3377), .B1(n4545), .B2(n3153), .ZN(n5131)
         );
  OAI221_X1 U721 ( .B1(n5446), .B2(n4546), .C1(n5638), .C2(n4547), .A(n5138), 
        .ZN(n5129) );
  AOI22_X1 U722 ( .A1(n4549), .A2(n3121), .B1(n4550), .B2(n2929), .ZN(n5138)
         );
  OAI221_X1 U723 ( .B1(n5414), .B2(n4551), .C1(n5542), .C2(n4552), .A(n5141), 
        .ZN(n5128) );
  AOI22_X1 U724 ( .A1(n4554), .A2(n3089), .B1(n4555), .B2(n2833), .ZN(n5141)
         );
  OAI221_X1 U725 ( .B1(n5574), .B2(n4556), .C1(n5318), .C2(n4557), .A(n5146), 
        .ZN(n5127) );
  AOI22_X1 U726 ( .A1(n4559), .A2(n3473), .B1(n4560), .B2(n2961), .ZN(n5146)
         );
  NOR2_X1 U727 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[0]), .ZN(n5143) );
  NOR4_X1 U728 ( .A1(n5147), .A2(n5148), .A3(n5149), .A4(n5150), .ZN(n5125) );
  OAI221_X1 U729 ( .B1(n5285), .B2(n4565), .C1(n5286), .C2(n4566), .A(n5151), 
        .ZN(n5150) );
  AOI22_X1 U730 ( .A1(n4568), .A2(n2801), .B1(n4569), .B2(n2737), .ZN(n5151)
         );
  AND3_X1 U731 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[2]), .ZN(n5142)
         );
  OAI221_X1 U732 ( .B1(n5606), .B2(n4570), .C1(n5284), .C2(n4571), .A(n5152), 
        .ZN(n5149) );
  AOI22_X1 U733 ( .A1(n4573), .A2(n3025), .B1(n4574), .B2(n3249), .ZN(n5152)
         );
  AND3_X1 U734 ( .A1(ADD_RD1[4]), .A2(n5153), .A3(ADD_RD1[2]), .ZN(n5144) );
  OAI221_X1 U735 ( .B1(n5670), .B2(n4575), .C1(n5478), .C2(n4576), .A(n5154), 
        .ZN(n5148) );
  AOI22_X1 U736 ( .A1(n4578), .A2(n3505), .B1(n4579), .B2(n3313), .ZN(n5154)
         );
  AND3_X1 U737 ( .A1(ADD_RD1[3]), .A2(n5155), .A3(ADD_RD1[2]), .ZN(n5145) );
  AND3_X1 U738 ( .A1(n5153), .A2(n5155), .A3(ADD_RD1[2]), .ZN(n5140) );
  NOR3_X1 U739 ( .A1(n5155), .A2(ADD_RD1[2]), .A3(n5153), .ZN(n5139) );
  NOR2_X1 U740 ( .A1(n5156), .A2(n5157), .ZN(n5134) );
  OAI221_X1 U741 ( .B1(n5283), .B2(n4580), .C1(n5350), .C2(n4581), .A(n5158), 
        .ZN(n5147) );
  AOI22_X1 U742 ( .A1(n4583), .A2(n3185), .B1(n4584), .B2(n3409), .ZN(n5158)
         );
  NOR3_X1 U743 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[4]), .A3(n5153), .ZN(n5135) );
  INV_X1 U744 ( .A(ADD_RD1[3]), .ZN(n5153) );
  NOR3_X1 U745 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[3]), .A3(n5155), .ZN(n5133) );
  INV_X1 U746 ( .A(ADD_RD1[4]), .ZN(n5155) );
  NOR2_X1 U747 ( .A1(n5156), .A2(ADD_RD1[0]), .ZN(n5132) );
  INV_X1 U748 ( .A(ADD_RD1[1]), .ZN(n5156) );
  NOR3_X1 U749 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[2]), .ZN(n5137)
         );
  NOR2_X1 U750 ( .A1(n5157), .A2(ADD_RD1[1]), .ZN(n5136) );
  INV_X1 U751 ( .A(ADD_RD1[0]), .ZN(n5157) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   n1, n4;

  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(n4) );
  INV_X1 U1 ( .A(n4), .ZN(n1) );
  INV_X4 U2 ( .A(n1), .ZN(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   n1, n4;

  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(n4) );
  INV_X1 U1 ( .A(n4), .ZN(n1) );
  INV_X4 U2 ( .A(n1), .ZN(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   n1, n4;

  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(n4) );
  INV_X1 U1 ( .A(n4), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(ENCLK) );
endmodule


module dlx ( RST, CLK );
  input RST, CLK;
  wire   \cw_dec[2] , \cw_mem[4] , \unit_control/n153 , \unit_control/n152 ,
         \unit_control/cw1delay[9] , \unit_control/next_state[1] ,
         \unit_control/next_state[0] , \unit_fetch/pc_regout[2] ,
         \unit_fetch/pc_regout[3] , \unit_fetch/pc_regout[4] ,
         \unit_fetch/pc_regout[5] , \unit_fetch/pc_regout[6] ,
         \unit_fetch/pc_regout[7] , \unit_fetch/pc_regout[8] ,
         \unit_fetch/pc_regout[10] , \unit_fetch/pc_regout[12] ,
         \unit_fetch/pc_regout[13] , \unit_fetch/pc_regout[14] ,
         \unit_fetch/pc_regout[15] , \unit_fetch/pc_regout[18] ,
         \unit_fetch/pc_regout[19] , \unit_fetch/pc_regout[20] ,
         \unit_fetch/pc_regout[22] , \unit_fetch/pc_regout[24] ,
         \unit_fetch/pc_regout[25] , \unit_fetch/pc_regout[26] ,
         \unit_fetch/pc_regout[27] , \unit_fetch/pc_regout[28] ,
         \unit_fetch/pc_regout[29] , \unit_fetch/pc_regout[30] ,
         \unit_decode/registerA[31] , \unit_decode/registerA[30] ,
         \unit_decode/registerA[29] , \unit_decode/registerA[28] ,
         \unit_decode/registerA[27] , \unit_decode/registerA[26] ,
         \unit_decode/registerA[25] , \unit_decode/registerA[24] ,
         \unit_decode/registerA[23] , \unit_decode/registerA[22] ,
         \unit_decode/registerA[21] , \unit_decode/registerA[20] ,
         \unit_decode/registerA[19] , \unit_decode/registerA[18] ,
         \unit_decode/registerA[17] , \unit_decode/registerA[16] ,
         \unit_decode/registerA[15] , \unit_decode/registerA[14] ,
         \unit_decode/registerA[13] , \unit_decode/registerA[12] ,
         \unit_decode/registerA[11] , \unit_decode/registerA[10] ,
         \unit_decode/registerA[9] , \unit_decode/registerA[8] ,
         \unit_decode/registerA[7] , \unit_decode/registerA[6] ,
         \unit_decode/registerA[5] , \unit_decode/registerA[4] ,
         \unit_decode/registerA[3] , \unit_decode/registerA[2] ,
         \unit_decode/registerA[1] , \unit_decode/registerA[0] ,
         \unit_decode/RS1s[4] , \unit_decode/RS1s[3] , \unit_decode/RS1s[2] ,
         \unit_decode/RS1s[1] , \unit_fetch/unit_instructionRegister/n98 ,
         \unit_fetch/unit_instructionRegister/n97 ,
         \unit_fetch/unit_instructionRegister/n96 ,
         \unit_fetch/unit_instructionRegister/n95 ,
         \unit_fetch/unit_instructionRegister/n94 ,
         \unit_fetch/unit_instructionRegister/n93 ,
         \unit_fetch/unit_instructionRegister/n90 ,
         \unit_fetch/unit_instructionRegister/n89 ,
         \unit_fetch/unit_instructionRegister/n88 ,
         \unit_fetch/unit_instructionRegister/n87 ,
         \unit_fetch/unit_instructionRegister/n82 ,
         \unit_fetch/unit_instructionRegister/n81 ,
         \unit_fetch/unit_instructionRegister/n80 ,
         \unit_fetch/unit_instructionRegister/n79 ,
         \unit_fetch/unit_instructionRegister/n78 ,
         \unit_fetch/unit_instructionRegister/n77 ,
         \unit_fetch/unit_instructionRegister/n75 ,
         \unit_fetch/unit_instructionRegister/n74 ,
         \unit_fetch/unit_instructionRegister/n73 ,
         \unit_fetch/unit_instructionRegister/n72 ,
         \unit_fetch/unit_instructionRegister/n71 ,
         \unit_fetch/unit_instructionRegister/n70 ,
         \unit_fetch/unit_instructionRegister/n68 ,
         \unit_fetch/unit_instructionRegister/n66 ,
         \unit_fetch/unit_instructionRegister/n65 ,
         \unit_fetch/unit_instructionRegister/n64 ,
         \unit_fetch/unit_instructionRegister/n63 ,
         \unit_fetch/unit_instructionRegister/n62 ,
         \unit_fetch/unit_instructionRegister/n61 ,
         \unit_fetch/unit_instructionRegister/n60 ,
         \unit_fetch/unit_instructionRegister/n59 ,
         \unit_fetch/unit_instructionRegister/n57 ,
         \unit_fetch/unit_instructionRegister/n56 ,
         \unit_fetch/unit_instructionRegister/n55 ,
         \unit_fetch/unit_instructionRegister/n54 ,
         \unit_fetch/unit_instructionRegister/n53 ,
         \unit_fetch/unit_instructionRegister/n52 ,
         \unit_fetch/unit_instructionRegister/n51 ,
         \unit_fetch/unit_instructionRegister/n49 ,
         \unit_fetch/unit_instructionRegister/n48 ,
         \unit_fetch/unit_instructionRegister/n47 ,
         \unit_fetch/unit_instructionRegister/n46 ,
         \unit_fetch/unit_instructionRegister/n45 ,
         \unit_fetch/unit_instructionRegister/n44 ,
         \unit_fetch/unit_instructionRegister/n43 ,
         \unit_fetch/unit_instructionRegister/n41 ,
         \unit_fetch/unit_instructionRegister/n40 ,
         \unit_fetch/unit_instructionRegister/n39 ,
         \unit_fetch/unit_instructionRegister/n38 ,
         \unit_decode/RD1reg/ffi_0/n4 , \unit_decode/RD1reg/ffi_1/n4 ,
         \unit_decode/RD1reg/ffi_2/n4 , \unit_decode/RD1reg/ffi_3/n4 ,
         \unit_decode/RD1reg/ffi_4/n4 , \unit_decode/IMMreg/ffi_0/n4 ,
         \unit_decode/IMMreg/ffi_1/n4 , \unit_decode/IMMreg/ffi_2/n4 ,
         \unit_decode/IMMreg/ffi_3/n4 , \unit_decode/IMMreg/ffi_4/n4 ,
         \unit_decode/IMMreg/ffi_5/n4 , \unit_decode/IMMreg/ffi_6/n4 ,
         \unit_decode/IMMreg/ffi_7/n4 , \unit_decode/IMMreg/ffi_8/n4 ,
         \unit_decode/IMMreg/ffi_9/n4 , \unit_decode/IMMreg/ffi_10/n4 ,
         \unit_decode/IMMreg/ffi_11/n4 , \unit_decode/IMMreg/ffi_12/n4 ,
         \unit_decode/IMMreg/ffi_13/n4 , \unit_decode/IMMreg/ffi_14/n4 ,
         \unit_decode/IMMreg/ffi_15/n4 , \unit_decode/IMMreg/ffi_16/n4 ,
         \unit_decode/IMMreg/ffi_17/n4 , \unit_decode/IMMreg/ffi_18/n4 ,
         \unit_decode/IMMreg/ffi_19/n4 , \unit_decode/IMMreg/ffi_20/n4 ,
         \unit_decode/IMMreg/ffi_21/n4 , \unit_decode/IMMreg/ffi_22/n4 ,
         \unit_decode/IMMreg/ffi_23/n4 , \unit_decode/IMMreg/ffi_24/n4 ,
         \unit_decode/IMMreg/ffi_25/n4 , \unit_decode/IMMreg/ffi_26/n4 ,
         \unit_decode/IMMreg/ffi_27/n4 , \unit_decode/IMMreg/ffi_28/n4 ,
         \unit_decode/IMMreg/ffi_29/n4 , \unit_decode/IMMreg/ffi_30/n4 ,
         \unit_decode/IMMreg/ffi_31/n4 , \unit_decode/Areg/ffi_0/n4 ,
         \unit_decode/Areg/ffi_1/n4 , \unit_decode/Areg/ffi_2/n4 ,
         \unit_decode/Areg/ffi_3/n4 , \unit_decode/Areg/ffi_4/n4 ,
         \unit_decode/Areg/ffi_5/n4 , \unit_decode/Areg/ffi_6/n4 ,
         \unit_decode/Areg/ffi_7/n4 , \unit_decode/Areg/ffi_8/n4 ,
         \unit_decode/Areg/ffi_9/n4 , \unit_decode/Areg/ffi_10/n4 ,
         \unit_decode/Areg/ffi_11/n4 , \unit_decode/Areg/ffi_12/n4 ,
         \unit_decode/Areg/ffi_13/n4 , \unit_decode/Areg/ffi_14/n4 ,
         \unit_decode/Areg/ffi_15/n4 , \unit_decode/Areg/ffi_16/n4 ,
         \unit_decode/Areg/ffi_17/n4 , \unit_decode/Areg/ffi_18/n4 ,
         \unit_decode/Areg/ffi_19/n4 , \unit_decode/Areg/ffi_20/n4 ,
         \unit_decode/Areg/ffi_21/n4 , \unit_decode/Areg/ffi_22/n4 ,
         \unit_decode/Areg/ffi_23/n4 , \unit_decode/Areg/ffi_24/n4 ,
         \unit_decode/Areg/ffi_25/n4 , \unit_decode/Areg/ffi_26/n4 ,
         \unit_decode/Areg/ffi_27/n4 , \unit_decode/Areg/ffi_28/n4 ,
         \unit_decode/Areg/ffi_29/n4 , \unit_decode/Areg/ffi_30/n4 ,
         \unit_decode/Areg/ffi_31/n4 , \unit_decode/NPC1reg/ffi_0/n4 ,
         \unit_decode/NPC1reg/ffi_1/n4 , \unit_decode/NPC1reg/ffi_2/n4 ,
         \unit_decode/NPC1reg/ffi_3/n4 , \unit_decode/NPC1reg/ffi_4/n4 ,
         \unit_decode/NPC1reg/ffi_5/n4 , \unit_decode/NPC1reg/ffi_6/n4 ,
         \unit_decode/NPC1reg/ffi_7/n4 , \unit_decode/NPC1reg/ffi_8/n4 ,
         \unit_decode/NPC1reg/ffi_9/n4 , \unit_decode/NPC1reg/ffi_10/n4 ,
         \unit_decode/NPC1reg/ffi_11/n4 , \unit_decode/NPC1reg/ffi_12/n4 ,
         \unit_decode/NPC1reg/ffi_13/n4 , \unit_decode/NPC1reg/ffi_14/n4 ,
         \unit_decode/NPC1reg/ffi_15/n4 , \unit_decode/NPC1reg/ffi_16/n4 ,
         \unit_decode/NPC1reg/ffi_17/n4 , \unit_decode/NPC1reg/ffi_18/n4 ,
         \unit_decode/NPC1reg/ffi_19/n4 , \unit_decode/NPC1reg/ffi_20/n4 ,
         \unit_decode/NPC1reg/ffi_21/n4 , \unit_decode/NPC1reg/ffi_22/n4 ,
         \unit_decode/NPC1reg/ffi_23/n4 , \unit_decode/NPC1reg/ffi_24/n4 ,
         \unit_decode/NPC1reg/ffi_25/n4 , \unit_decode/NPC1reg/ffi_26/n4 ,
         \unit_decode/NPC1reg/ffi_27/n4 , \unit_decode/NPC1reg/ffi_28/n4 ,
         \unit_decode/NPC1reg/ffi_29/n4 , \unit_decode/NPC1reg/ffi_30/n4 ,
         \unit_decode/NPC1reg/ffi_31/n4 ,
         \unit_fetch/unit_npcregister/ffi_0/n4 ,
         \unit_fetch/unit_npcregister/ffi_1/n4 ,
         \unit_fetch/unit_npcregister/ffi_2/n4 ,
         \unit_fetch/unit_npcregister/ffi_3/n4 ,
         \unit_fetch/unit_npcregister/ffi_4/n4 ,
         \unit_fetch/unit_npcregister/ffi_5/n4 ,
         \unit_fetch/unit_npcregister/ffi_6/n4 ,
         \unit_fetch/unit_npcregister/ffi_7/n4 ,
         \unit_fetch/unit_npcregister/ffi_8/n4 ,
         \unit_fetch/unit_npcregister/ffi_9/n4 ,
         \unit_fetch/unit_npcregister/ffi_10/n4 ,
         \unit_fetch/unit_npcregister/ffi_11/n4 ,
         \unit_fetch/unit_npcregister/ffi_12/n4 ,
         \unit_fetch/unit_npcregister/ffi_13/n4 ,
         \unit_fetch/unit_npcregister/ffi_14/n4 ,
         \unit_fetch/unit_npcregister/ffi_15/n4 ,
         \unit_fetch/unit_npcregister/ffi_16/n4 ,
         \unit_fetch/unit_npcregister/ffi_17/n4 ,
         \unit_fetch/unit_npcregister/ffi_18/n4 ,
         \unit_fetch/unit_npcregister/ffi_19/n4 ,
         \unit_fetch/unit_npcregister/ffi_20/n4 ,
         \unit_fetch/unit_npcregister/ffi_21/n4 ,
         \unit_fetch/unit_npcregister/ffi_22/n4 ,
         \unit_fetch/unit_npcregister/ffi_23/n4 ,
         \unit_fetch/unit_npcregister/ffi_24/n4 ,
         \unit_fetch/unit_npcregister/ffi_25/n4 ,
         \unit_fetch/unit_npcregister/ffi_26/n4 ,
         \unit_fetch/unit_npcregister/ffi_27/n4 ,
         \unit_fetch/unit_npcregister/ffi_28/n4 ,
         \unit_fetch/unit_npcregister/ffi_29/n4 ,
         \unit_fetch/unit_npcregister/ffi_30/n4 ,
         \unit_fetch/unit_npcregister/ffi_31/n4 ,
         \unit_fetch/unit_programCounter/ffi_0/n5 ,
         \unit_fetch/unit_programCounter/ffi_0/n4 ,
         \unit_fetch/unit_programCounter/ffi_1/n5 ,
         \unit_fetch/unit_programCounter/ffi_1/n4 ,
         \unit_fetch/unit_programCounter/ffi_3/n5 ,
         \unit_fetch/unit_programCounter/ffi_4/n5 ,
         \unit_fetch/unit_programCounter/ffi_6/n5 ,
         \unit_fetch/unit_programCounter/ffi_8/n5 ,
         \unit_fetch/unit_programCounter/ffi_10/n5 ,
         \unit_fetch/unit_programCounter/ffi_12/n5 ,
         \unit_fetch/unit_programCounter/ffi_14/n5 ,
         \unit_fetch/unit_programCounter/ffi_16/n5 ,
         \unit_fetch/unit_programCounter/ffi_18/n5 ,
         \unit_fetch/unit_programCounter/ffi_19/n5 ,
         \unit_fetch/unit_programCounter/ffi_20/n5 ,
         \unit_fetch/unit_programCounter/ffi_22/n5 ,
         \unit_fetch/unit_programCounter/ffi_24/n5 ,
         \unit_fetch/unit_programCounter/ffi_26/n5 ,
         \unit_fetch/unit_programCounter/ffi_28/n5 ,
         \unit_fetch/unit_programCounter/ffi_29/n5 ,
         \unit_fetch/unit_programCounter/ffi_31/n5 ,
         \unit_control/uut_fourth_stage/ffi_3/n6 ,
         \unit_control/uut_fourth_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_3/n5 ,
         \unit_control/uut_third_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_9/n6 ,
         \unit_control/uut_third_stage/ffi_10/n5 ,
         \unit_control/uut_third_stage/ffi_12/n5 ,
         \unit_control/uut_third_stage/ffi_13/n5 ,
         \unit_control/uut_third_stage/ffi_14/n5 ,
         \unit_control/uut_third_stage/ffi_15/n5 ,
         \unit_control/uut_third_stage/ffi_17/n6 ,
         \unit_control/uut_third_stage/ffi_17/n5 ,
         \unit_control/uut_third_stage/ffi_19/n5 ,
         \unit_control/uut_second_stage/ffi_10/n5 ,
         \unit_control/uut_second_stage/ffi_12/n5 ,
         \unit_control/uut_second_stage/ffi_13/n5 ,
         \unit_control/uut_second_stage/ffi_17/n5 , n1337, n1394, n2598, n2599,
         n2600, n2617, n2618, n2619, n2620, n2621, n2912, n3095, n3676, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064;
  wire   [4:0] wr_address;
  wire   [31:0] wr_data;

  DFFR_X1 \unit_control/current_state_reg[1]  ( .D(
        \unit_control/next_state[1] ), .CK(CLK), .RN(n2912), .Q(
        \unit_control/n152 ) );
  DFFR_X1 \unit_control/current_state_reg[0]  ( .D(
        \unit_control/next_state[0] ), .CK(CLK), .RN(n2912), .Q(
        \unit_control/n153 ) );
  register_file_WORD_SIZE32_ADDR_SIZE5 \unit_decode/RegisterFile  ( .CLK(CLK), 
        .RESET(RST), .ENABLE(\cw_dec[2] ), .RD1(\unit_control/cw1delay[9] ), 
        .RD2(1'b0), .WR(\cw_mem[4] ), .ADD_WR(wr_address), .ADD_RD1({
        \unit_decode/RS1s[4] , \unit_decode/RS1s[3] , \unit_decode/RS1s[2] , 
        \unit_decode/RS1s[1] , n1394}), .ADD_RD2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATAIN(wr_data), .OUT1({\unit_decode/registerA[31] , 
        \unit_decode/registerA[30] , \unit_decode/registerA[29] , 
        \unit_decode/registerA[28] , \unit_decode/registerA[27] , 
        \unit_decode/registerA[26] , \unit_decode/registerA[25] , 
        \unit_decode/registerA[24] , \unit_decode/registerA[23] , 
        \unit_decode/registerA[22] , \unit_decode/registerA[21] , 
        \unit_decode/registerA[20] , \unit_decode/registerA[19] , 
        \unit_decode/registerA[18] , \unit_decode/registerA[17] , 
        \unit_decode/registerA[16] , \unit_decode/registerA[15] , 
        \unit_decode/registerA[14] , \unit_decode/registerA[13] , 
        \unit_decode/registerA[12] , \unit_decode/registerA[11] , 
        \unit_decode/registerA[10] , \unit_decode/registerA[9] , 
        \unit_decode/registerA[8] , \unit_decode/registerA[7] , 
        \unit_decode/registerA[6] , \unit_decode/registerA[5] , 
        \unit_decode/registerA[4] , \unit_decode/registerA[3] , 
        \unit_decode/registerA[2] , \unit_decode/registerA[1] , 
        \unit_decode/registerA[0] }) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[0]  ( .D(
        \unit_fetch/unit_instructionRegister/n98 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n38 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[1]  ( .D(
        \unit_fetch/unit_instructionRegister/n97 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n39 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[2]  ( .D(
        \unit_fetch/unit_instructionRegister/n96 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n40 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[3]  ( .D(
        \unit_fetch/unit_instructionRegister/n95 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n41 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[5]  ( .D(
        \unit_fetch/unit_instructionRegister/n93 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n43 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[6]  ( .D(
        \unit_fetch/unit_instructionRegister/n94 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n44 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[7]  ( .D(n2619), .CK(
        CLK), .QN(\unit_fetch/unit_instructionRegister/n45 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[8]  ( .D(
        \unit_fetch/unit_instructionRegister/n90 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n46 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[9]  ( .D(
        \unit_fetch/unit_instructionRegister/n89 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n47 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[10]  ( .D(
        \unit_fetch/unit_instructionRegister/n88 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n48 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[11]  ( .D(
        \unit_fetch/unit_instructionRegister/n87 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n49 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[13]  ( .D(n3770), 
        .CK(CLK), .QN(\unit_fetch/unit_instructionRegister/n51 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[14]  ( .D(n2617), 
        .CK(CLK), .QN(\unit_fetch/unit_instructionRegister/n52 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[15]  ( .D(n2618), 
        .CK(CLK), .Q(n3799), .QN(\unit_fetch/unit_instructionRegister/n53 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[16]  ( .D(
        \unit_fetch/unit_instructionRegister/n82 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n54 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[18]  ( .D(
        \unit_fetch/unit_instructionRegister/n80 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n56 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[19]  ( .D(
        \unit_fetch/unit_instructionRegister/n79 ), .CK(CLK), .Q(n3801), .QN(
        \unit_fetch/unit_instructionRegister/n57 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[21]  ( .D(
        \unit_fetch/unit_instructionRegister/n77 ), .CK(CLK), .Q(n1394), .QN(
        \unit_fetch/unit_instructionRegister/n59 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[23]  ( .D(n2621), 
        .CK(CLK), .Q(\unit_decode/RS1s[2] ), .QN(
        \unit_fetch/unit_instructionRegister/n61 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[24]  ( .D(
        \unit_fetch/unit_instructionRegister/n75 ), .CK(CLK), .Q(
        \unit_decode/RS1s[3] ), .QN(\unit_fetch/unit_instructionRegister/n62 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[25]  ( .D(
        \unit_fetch/unit_instructionRegister/n74 ), .CK(CLK), .Q(
        \unit_decode/RS1s[4] ), .QN(\unit_fetch/unit_instructionRegister/n63 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[26]  ( .D(
        \unit_fetch/unit_instructionRegister/n68 ), .CK(CLK), .QN(n4863) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[27]  ( .D(
        \unit_fetch/unit_instructionRegister/n73 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n64 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[28]  ( .D(
        \unit_fetch/unit_instructionRegister/n70 ), .CK(CLK), .QN(n3798) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[29]  ( .D(
        \unit_fetch/unit_instructionRegister/n72 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n65 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[31]  ( .D(
        \unit_fetch/unit_instructionRegister/n71 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n66 ) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_0/Q_reg  ( .D(n4900), .CK(n4969), 
        .Q(wr_address[0]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_1/Q_reg  ( .D(n4901), .CK(n4969), 
        .Q(wr_address[1]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_2/Q_reg  ( .D(n4902), .CK(n4969), 
        .Q(wr_address[2]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_3/Q_reg  ( .D(n4903), .CK(n4969), 
        .Q(wr_address[3]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_4/Q_reg  ( .D(n4904), .CK(n4969), 
        .Q(wr_address[4]) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_0/Q_reg  ( .D(n4905), .CK(n4969), 
        .Q(n4851) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_2/Q_reg  ( .D(n4906), .CK(n4969), 
        .Q(n4807) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_3/Q_reg  ( .D(n4907), .CK(n4969), 
        .Q(n4801) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_4/Q_reg  ( .D(n4908), .CK(n4969), 
        .Q(n4799) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_5/Q_reg  ( .D(n4909), .CK(n4969), 
        .Q(n4797) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_6/Q_reg  ( .D(n4910), .CK(n4969), 
        .Q(n4795) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_7/Q_reg  ( .D(n4911), .CK(n4969), 
        .Q(n4793) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_8/Q_reg  ( .D(n4912), .CK(n4969), 
        .Q(n4791) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_9/Q_reg  ( .D(n4913), .CK(n4969), 
        .Q(n4789) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_10/Q_reg  ( .D(n4914), .CK(n4969), .Q(n4849) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_11/Q_reg  ( .D(n4915), .CK(n4969), .Q(n4847) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_12/Q_reg  ( .D(n4916), .CK(n4969), .Q(n4845) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_13/Q_reg  ( .D(n4917), .CK(n4969), .Q(n4843) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_14/Q_reg  ( .D(n4918), .CK(n4969), .Q(n4841) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_15/Q_reg  ( .D(n4919), .CK(n4969), .Q(n4839) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_16/Q_reg  ( .D(n4920), .CK(n4969), .Q(n4837) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_17/Q_reg  ( .D(n4921), .CK(n4969), .Q(n4835) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_18/Q_reg  ( .D(n4922), .CK(n4969), .Q(n4833) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_19/Q_reg  ( .D(n4923), .CK(n4969), .Q(n4831) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_20/Q_reg  ( .D(n4924), .CK(n4969), .Q(n4827) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_21/Q_reg  ( .D(n4925), .CK(n4969), .Q(n4825) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_22/Q_reg  ( .D(n4926), .CK(n4969), .Q(n4823) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_23/Q_reg  ( .D(n4927), .CK(n4969), .Q(n4821) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_24/Q_reg  ( .D(n4928), .CK(n4969), .Q(n4819) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_25/Q_reg  ( .D(n4929), .CK(n4969), .Q(n4817) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_26/Q_reg  ( .D(n4930), .CK(n4969), .Q(n4815) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_27/Q_reg  ( .D(n4931), .CK(n4969), .Q(n4813) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_28/Q_reg  ( .D(n4932), .CK(n4969), .Q(n4811) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_29/Q_reg  ( .D(n4933), .CK(n4969), .Q(n4809) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_30/Q_reg  ( .D(n4934), .CK(n4969), .Q(n4805) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_31/Q_reg  ( .D(n4935), .CK(n4969), .Q(n4803) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_0/Q_reg  ( .D(n4936), .CK(n4969), .Q(
        n4852) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_1/Q_reg  ( .D(n4937), .CK(n4969), .Q(
        n4830) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_2/Q_reg  ( .D(n4938), .CK(n4969), .Q(
        n4808) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_3/Q_reg  ( .D(n4939), .CK(n4969), .Q(
        n4802) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_4/Q_reg  ( .D(n4940), .CK(n4969), .Q(
        n4800) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_5/Q_reg  ( .D(n4941), .CK(n4969), .Q(
        n4798) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_6/Q_reg  ( .D(n4942), .CK(n4969), .Q(
        n4796) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_7/Q_reg  ( .D(n4943), .CK(n4969), .Q(
        n4794) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_8/Q_reg  ( .D(n4944), .CK(n4969), .Q(
        n4792) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_9/Q_reg  ( .D(n4945), .CK(n4969), .Q(
        n4790) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_10/Q_reg  ( .D(n4946), .CK(n4969), .Q(
        n4850) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_11/Q_reg  ( .D(n4947), .CK(n4969), .Q(
        n4848) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_12/Q_reg  ( .D(n4948), .CK(n4969), .Q(
        n4846) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_13/Q_reg  ( .D(n4949), .CK(n4969), .Q(
        n4844) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_14/Q_reg  ( .D(n4950), .CK(n4969), .Q(
        n4842) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_15/Q_reg  ( .D(n4951), .CK(n4969), .Q(
        n4840) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_16/Q_reg  ( .D(n4952), .CK(n4969), .Q(
        n4838) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_17/Q_reg  ( .D(n4953), .CK(n4969), .Q(
        n4836) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_18/Q_reg  ( .D(n4954), .CK(n4969), .Q(
        n4834) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_19/Q_reg  ( .D(n4955), .CK(n4969), .Q(
        n4832) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_20/Q_reg  ( .D(n4956), .CK(n4969), .Q(
        n4828) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_21/Q_reg  ( .D(n4957), .CK(n4969), .Q(
        n4826) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_22/Q_reg  ( .D(n4958), .CK(n4969), .Q(
        n4824) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_23/Q_reg  ( .D(n4959), .CK(n4969), .Q(
        n4822) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_24/Q_reg  ( .D(n4960), .CK(n4969), .Q(
        n4820) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_25/Q_reg  ( .D(n4961), .CK(n4969), .Q(
        n4818) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_26/Q_reg  ( .D(n4962), .CK(n4969), .Q(
        n4816) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_27/Q_reg  ( .D(n4963), .CK(n4969), .Q(
        n4814) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_28/Q_reg  ( .D(n4964), .CK(n4969), .Q(
        n4812) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_29/Q_reg  ( .D(n4965), .CK(n4969), .Q(
        n4810) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_30/Q_reg  ( .D(n4966), .CK(n4969), .Q(
        n4806) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_31/Q_reg  ( .D(n4967), .CK(n4969), .Q(
        n4804) );
  DFF_X1 \unit_decode/RD1reg/ffi_0/Q_reg  ( .D(n4971), .CK(n5064), .QN(
        \unit_decode/RD1reg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_1/Q_reg  ( .D(n4972), .CK(n5064), .QN(
        \unit_decode/RD1reg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_2/Q_reg  ( .D(n4973), .CK(n5064), .QN(
        \unit_decode/RD1reg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_3/Q_reg  ( .D(n4974), .CK(n5064), .QN(
        \unit_decode/RD1reg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_4/Q_reg  ( .D(n4975), .CK(n5064), .QN(
        \unit_decode/RD1reg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_0/Q_reg  ( .D(n4976), .CK(n5064), .Q(n3786), 
        .QN(\unit_decode/IMMreg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_1/Q_reg  ( .D(n4977), .CK(n5064), .Q(n3781), 
        .QN(\unit_decode/IMMreg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_2/Q_reg  ( .D(n4978), .CK(n5064), .Q(n3790), 
        .QN(\unit_decode/IMMreg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_3/Q_reg  ( .D(n4979), .CK(n5064), .Q(n3778), 
        .QN(\unit_decode/IMMreg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_4/Q_reg  ( .D(n4981), .CK(n5064), .Q(n3787), 
        .QN(\unit_decode/IMMreg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_5/Q_reg  ( .D(n4980), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_6/Q_reg  ( .D(n4981), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_7/Q_reg  ( .D(n4982), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_8/Q_reg  ( .D(n4983), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_8/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_9/Q_reg  ( .D(n4984), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_10/Q_reg  ( .D(n4985), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_10/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_11/Q_reg  ( .D(n4986), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_12/Q_reg  ( .D(n4988), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_12/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_13/Q_reg  ( .D(n4987), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_14/Q_reg  ( .D(n4988), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_15/Q_reg  ( .D(n4989), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_16/Q_reg  ( .D(n4990), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_17/Q_reg  ( .D(n4991), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_18/Q_reg  ( .D(n4992), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_19/Q_reg  ( .D(n4993), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_19/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_20/Q_reg  ( .D(n4994), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_21/Q_reg  ( .D(n4995), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_22/Q_reg  ( .D(n4994), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_23/Q_reg  ( .D(n4996), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_24/Q_reg  ( .D(n4997), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_25/Q_reg  ( .D(n4998), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_25/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_26/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_26/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_27/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_27/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_28/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_28/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_29/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_29/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_30/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_30/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_31/Q_reg  ( .D(n4999), .CK(n5064), .QN(
        \unit_decode/IMMreg/ffi_31/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_0/Q_reg  ( .D(n5000), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_1/Q_reg  ( .D(n5001), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_2/Q_reg  ( .D(n5002), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_3/Q_reg  ( .D(n5003), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_4/Q_reg  ( .D(n5004), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_5/Q_reg  ( .D(n5005), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_6/Q_reg  ( .D(n5006), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_7/Q_reg  ( .D(n5007), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_8/Q_reg  ( .D(n5008), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_8/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_9/Q_reg  ( .D(n5009), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_10/Q_reg  ( .D(n5010), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_10/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_11/Q_reg  ( .D(n5011), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_12/Q_reg  ( .D(n5012), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_12/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_13/Q_reg  ( .D(n5013), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_14/Q_reg  ( .D(n5014), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_15/Q_reg  ( .D(n5015), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_16/Q_reg  ( .D(n5016), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_17/Q_reg  ( .D(n5017), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_18/Q_reg  ( .D(n5018), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_19/Q_reg  ( .D(n5019), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_19/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_20/Q_reg  ( .D(n5020), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_21/Q_reg  ( .D(n5021), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_22/Q_reg  ( .D(n5022), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_23/Q_reg  ( .D(n5023), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_24/Q_reg  ( .D(n5024), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_25/Q_reg  ( .D(n5025), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_25/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_26/Q_reg  ( .D(n5026), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_26/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_27/Q_reg  ( .D(n5027), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_27/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_28/Q_reg  ( .D(n5028), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_28/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_29/Q_reg  ( .D(n5029), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_29/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_30/Q_reg  ( .D(n5030), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_30/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_31/Q_reg  ( .D(n5031), .CK(n5064), .QN(
        \unit_decode/Areg/ffi_31/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_0/Q_reg  ( .D(n5032), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_1/Q_reg  ( .D(n5033), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_2/Q_reg  ( .D(n5034), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_3/Q_reg  ( .D(n5035), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_4/Q_reg  ( .D(n5036), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_5/Q_reg  ( .D(n5037), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_6/Q_reg  ( .D(n5038), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_7/Q_reg  ( .D(n5039), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_8/Q_reg  ( .D(n5040), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_8/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_9/Q_reg  ( .D(n5041), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_10/Q_reg  ( .D(n5042), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_10/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_11/Q_reg  ( .D(n5043), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_12/Q_reg  ( .D(n5044), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_12/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_13/Q_reg  ( .D(n5045), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_14/Q_reg  ( .D(n5046), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_15/Q_reg  ( .D(n5047), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_16/Q_reg  ( .D(n5048), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_17/Q_reg  ( .D(n5049), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_18/Q_reg  ( .D(n5050), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_19/Q_reg  ( .D(n5051), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_19/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_20/Q_reg  ( .D(n5052), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_21/Q_reg  ( .D(n5053), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_22/Q_reg  ( .D(n5054), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_23/Q_reg  ( .D(n5055), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_24/Q_reg  ( .D(n5056), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_25/Q_reg  ( .D(n5057), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_25/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_26/Q_reg  ( .D(n5058), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_26/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_27/Q_reg  ( .D(n5059), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_27/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_28/Q_reg  ( .D(n5060), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_28/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_29/Q_reg  ( .D(n5061), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_29/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_30/Q_reg  ( .D(n5062), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_30/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_31/Q_reg  ( .D(n5063), .CK(n5064), .QN(
        \unit_decode/NPC1reg/ffi_31/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_0/Q_reg  ( .D(n4865), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_0/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_1/Q_reg  ( .D(n4866), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_1/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_2/Q_reg  ( .D(n4867), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_2/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_3/Q_reg  ( .D(n4868), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_3/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_4/Q_reg  ( .D(n4869), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_4/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_5/Q_reg  ( .D(n4870), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_5/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_6/Q_reg  ( .D(n4871), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_6/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_7/Q_reg  ( .D(n4872), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_7/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_8/Q_reg  ( .D(n4873), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_8/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_9/Q_reg  ( .D(n4874), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_9/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_10/Q_reg  ( .D(n4875), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_10/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_11/Q_reg  ( .D(n4876), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_11/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_12/Q_reg  ( .D(n4877), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_12/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_13/Q_reg  ( .D(n4878), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_13/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_14/Q_reg  ( .D(n4879), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_14/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_15/Q_reg  ( .D(n4880), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_15/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_16/Q_reg  ( .D(n4881), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_16/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_17/Q_reg  ( .D(n4882), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_17/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_18/Q_reg  ( .D(n4883), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_18/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_19/Q_reg  ( .D(n4884), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_19/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_20/Q_reg  ( .D(n4885), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_20/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_21/Q_reg  ( .D(n4886), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_21/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_22/Q_reg  ( .D(n4887), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_22/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_23/Q_reg  ( .D(n4888), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_23/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_24/Q_reg  ( .D(n4889), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_24/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_25/Q_reg  ( .D(n4890), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_25/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_26/Q_reg  ( .D(n4891), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_26/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_27/Q_reg  ( .D(n4892), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_27/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_28/Q_reg  ( .D(n4893), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_28/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_29/Q_reg  ( .D(n4894), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_29/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_30/Q_reg  ( .D(n4895), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_30/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_31/Q_reg  ( .D(n4896), .CK(n4897), 
        .QN(\unit_fetch/unit_npcregister/ffi_31/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_0/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_0/n5 ), .CK(n4897), .Q(n3779), 
        .QN(\unit_fetch/unit_programCounter/ffi_0/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_1/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_1/n5 ), .CK(n4897), .Q(n3788), 
        .QN(\unit_fetch/unit_programCounter/ffi_1/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_2/Q_reg  ( .D(n4867), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[2] ), .QN(n3771) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_3/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_3/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[3] ), .QN(n3773) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_4/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_4/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[4] ), .QN(n3789) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_5/Q_reg  ( .D(n4870), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[5] ), .QN(n3780) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_6/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_6/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[6] ), .QN(n3797) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_7/Q_reg  ( .D(n4872), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[7] ), .QN(n3784) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_8/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_8/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[8] ), .QN(n3772) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_9/Q_reg  ( .D(n4874), .CK(n4897), 
        .QN(n3777) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_10/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_10/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[10] ), .QN(n3791) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_11/Q_reg  ( .D(n4876), .CK(n4897), 
        .QN(n4854) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_12/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_12/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[12] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_13/Q_reg  ( .D(n4878), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[13] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_14/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_14/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[14] ), .QN(n3783) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_15/Q_reg  ( .D(n4880), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[15] ), .QN(n3796) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_16/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_16/n5 ), .CK(n4897), .QN(n3774) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_17/Q_reg  ( .D(n4882), .CK(n4897), 
        .QN(n4855) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_18/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_18/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[18] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_19/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_19/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[19] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_20/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_20/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[20] ), .QN(n3792) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_21/Q_reg  ( .D(n4886), .CK(n4897), 
        .QN(n4856) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_22/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_22/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[22] ), .QN(n3775) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_23/Q_reg  ( .D(n4888), .CK(n4897), 
        .QN(n3794) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_24/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_24/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[24] ), .QN(n3782) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_25/Q_reg  ( .D(n4890), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[25] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_26/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_26/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[26] ), .QN(n3793) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_27/Q_reg  ( .D(n4892), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[27] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_28/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_28/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[28] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_29/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_29/n5 ), .CK(n4897), .Q(
        \unit_fetch/pc_regout[29] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_30/Q_reg  ( .D(n4895), .CK(n4897), 
        .Q(\unit_fetch/pc_regout[30] ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_31/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_31/n5 ), .CK(n4897), .QN(n4857) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_4/n5 ), .CK(CLK), .Q(\cw_mem[4] )
         );
  DFF_X1 \unit_control/uut_third_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_3/n5 ), .CK(CLK), .QN(n3752) );
  DFF_X1 \unit_control/uut_third_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_4/n5 ), .CK(CLK), .QN(n3753) );
  DFF_X1 \unit_control/uut_third_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_13/n5 ), .CK(CLK), .Q(n3795), .QN(
        n4860) );
  DFF_X1 \unit_control/uut_third_stage/ffi_14/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_14/n5 ), .CK(CLK), .QN(n4859) );
  DFF_X1 \unit_control/uut_third_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_17/n6 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_17/n5 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_19/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_15/n5 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_19/n5 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_3/Q_reg  ( .D(n2598), .CK(CLK), 
        .QN(n3759) );
  DFF_X1 \unit_control/uut_second_stage/ffi_4/Q_reg  ( .D(n3768), .CK(CLK), 
        .QN(n3760) );
  DFF_X1 \unit_control/uut_second_stage/ffi_9/Q_reg  ( .D(n2620), .CK(CLK), 
        .Q(\unit_control/cw1delay[9] ), .QN(n3761) );
  DFF_X1 \unit_control/uut_second_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_10/n5 ), .CK(CLK), .QN(n3754) );
  DFF_X1 \unit_control/uut_second_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_12/n5 ), .CK(CLK), .QN(n3755) );
  DFF_X1 \unit_control/uut_second_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_13/n5 ), .CK(CLK), .QN(n3756) );
  DFF_X1 \unit_control/uut_second_stage/ffi_14/Q_reg  ( .D(n3769), .CK(CLK), 
        .QN(n3757) );
  DFF_X1 \unit_control/uut_second_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_17/n5 ), .CK(CLK), .QN(n3758) );
  DFF_X1 \unit_control/uut_second_stage/ffi_20/Q_reg  ( .D(n2599), .CK(CLK), 
        .QN(n3776) );
  DFF_X1 \unit_control/uut_second_stage/ffi_21/Q_reg  ( .D(n2600), .CK(CLK), 
        .QN(n4864) );
  DFF_X1 \unit_control/uut_second_stage/ffi_22/Q_reg  ( .D(n2912), .CK(CLK), 
        .Q(\cw_dec[2] ), .QN(n1337) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[17]  ( .D(
        \unit_fetch/unit_instructionRegister/n81 ), .CK(CLK), .Q(n3800), .QN(
        \unit_fetch/unit_instructionRegister/n55 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_1/Q_reg  ( .D(n4968), .CK(n4969), 
        .Q(n4829) );
  DFF_X1 \unit_control/uut_third_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_10/n5 ), .CK(CLK), .QN(n4861) );
  DFF_X1 \unit_control/uut_third_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_12/n5 ), .CK(CLK), .QN(n4853) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[22]  ( .D(
        \unit_fetch/unit_instructionRegister/n78 ), .CK(CLK), .Q(
        \unit_decode/RS1s[1] ), .QN(\unit_fetch/unit_instructionRegister/n60 )
         );
  SNPS_CLOCK_GATE_HIGH_dlx_0 \clk_gate_unit_decode/NPC1reg/ffi_31/Q_reg  ( 
        .CLK(CLK), .EN(n3676), .ENCLK(n5064), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dlx_1 \clk_gate_unit_execution/COMP_REGN_ALUOUT/ffi_1/Q_reg  ( 
        .CLK(CLK), .EN(n3095), .ENCLK(n4969), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dlx_2 \clk_gate_unit_fetch/unit_programCounter/ffi_30/Q_reg  ( 
        .CLK(CLK), .EN(n4899), .ENCLK(n4897), .TE(1'b0) );
  DFF_X2 \unit_control/uut_third_stage/ffi_9/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_9/n6 ), .CK(CLK), .Q(n3785), .QN(
        n4862) );
  DFF_X2 \unit_control/uut_fourth_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_3/n6 ), .CK(CLK), .QN(n4858) );
  AOI221_X1 U3194 ( .B1(n4121), .B2(n4505), .C1(n4106), .C2(n4051), .A(n4628), 
        .ZN(n4613) );
  NAND3_X2 U3195 ( .A1(\unit_decode/IMMreg/ffi_3/n4 ), .A2(
        \unit_decode/IMMreg/ffi_4/n4 ), .A3(n4693), .ZN(n4272) );
  INV_X2 U3196 ( .A(n4193), .ZN(n4106) );
  AOI222_X1 U3197 ( .A1(n4030), .A2(n4119), .B1(n4107), .B2(n4028), .C1(n4033), 
        .C2(n4120), .ZN(n4111) );
  NOR2_X2 U3198 ( .A1(n4153), .A2(n4201), .ZN(n4030) );
  NOR2_X2 U3199 ( .A1(n4149), .A2(n4201), .ZN(n4121) );
  NOR2_X4 U3200 ( .A1(n4154), .A2(n4201), .ZN(n4177) );
  NOR2_X4 U3201 ( .A1(n4139), .A2(n4201), .ZN(n4120) );
  INV_X2 U3202 ( .A(n4134), .ZN(n4024) );
  NOR2_X4 U3203 ( .A1(n4201), .A2(n4147), .ZN(n4118) );
  NOR2_X2 U3204 ( .A1(n4012), .A2(n3829), .ZN(n3921) );
  NOR3_X2 U3205 ( .A1(n4862), .A2(n4861), .A3(n4097), .ZN(n4624) );
  NAND2_X2 U3206 ( .A1(n3825), .A2(n4012), .ZN(n3913) );
  NOR2_X2 U3207 ( .A1(n4165), .A2(n4853), .ZN(n4126) );
  NOR2_X4 U3208 ( .A1(n4151), .A2(n4201), .ZN(n4017) );
  NOR2_X2 U3209 ( .A1(n4013), .A2(RST), .ZN(n3825) );
  INV_X2 U3210 ( .A(RST), .ZN(n2912) );
  INV_X2 U3211 ( .A(\unit_control/uut_third_stage/ffi_19/n5 ), .ZN(n4012) );
  NOR2_X2 U3212 ( .A1(n4165), .A2(n4861), .ZN(n4036) );
  NOR2_X4 U3213 ( .A1(n4143), .A2(n4201), .ZN(n4028) );
  MUX2_X1 U3214 ( .A(n4790), .B(n4789), .S(n4858), .Z(wr_data[9]) );
  MUX2_X1 U3215 ( .A(n4792), .B(n4791), .S(n4858), .Z(wr_data[8]) );
  MUX2_X1 U3216 ( .A(n4794), .B(n4793), .S(n4858), .Z(wr_data[7]) );
  MUX2_X1 U3217 ( .A(n4796), .B(n4795), .S(n4858), .Z(wr_data[6]) );
  MUX2_X1 U3218 ( .A(n4798), .B(n4797), .S(n4858), .Z(wr_data[5]) );
  MUX2_X1 U3219 ( .A(n4800), .B(n4799), .S(n4858), .Z(wr_data[4]) );
  MUX2_X1 U3220 ( .A(n4802), .B(n4801), .S(n4858), .Z(wr_data[3]) );
  MUX2_X1 U3221 ( .A(n4804), .B(n4803), .S(n4858), .Z(wr_data[31]) );
  MUX2_X1 U3222 ( .A(n4806), .B(n4805), .S(n4858), .Z(wr_data[30]) );
  MUX2_X1 U3223 ( .A(n4808), .B(n4807), .S(n4858), .Z(wr_data[2]) );
  MUX2_X1 U3224 ( .A(n4810), .B(n4809), .S(n4858), .Z(wr_data[29]) );
  MUX2_X1 U3225 ( .A(n4812), .B(n4811), .S(n4858), .Z(wr_data[28]) );
  MUX2_X1 U3226 ( .A(n4814), .B(n4813), .S(n4858), .Z(wr_data[27]) );
  MUX2_X1 U3227 ( .A(n4816), .B(n4815), .S(n4858), .Z(wr_data[26]) );
  MUX2_X1 U3228 ( .A(n4818), .B(n4817), .S(n4858), .Z(wr_data[25]) );
  MUX2_X1 U3229 ( .A(n4820), .B(n4819), .S(n4858), .Z(wr_data[24]) );
  MUX2_X1 U3230 ( .A(n4822), .B(n4821), .S(n4858), .Z(wr_data[23]) );
  MUX2_X1 U3231 ( .A(n4824), .B(n4823), .S(n4858), .Z(wr_data[22]) );
  MUX2_X1 U3232 ( .A(n4826), .B(n4825), .S(n4858), .Z(wr_data[21]) );
  MUX2_X1 U3233 ( .A(n4828), .B(n4827), .S(n4858), .Z(wr_data[20]) );
  MUX2_X1 U3234 ( .A(n4830), .B(n4829), .S(n4858), .Z(wr_data[1]) );
  MUX2_X1 U3235 ( .A(n4832), .B(n4831), .S(n4858), .Z(wr_data[19]) );
  MUX2_X1 U3236 ( .A(n4834), .B(n4833), .S(n4858), .Z(wr_data[18]) );
  MUX2_X1 U3237 ( .A(n4836), .B(n4835), .S(n4858), .Z(wr_data[17]) );
  MUX2_X1 U3238 ( .A(n4838), .B(n4837), .S(n4858), .Z(wr_data[16]) );
  MUX2_X1 U3239 ( .A(n4840), .B(n4839), .S(n4858), .Z(wr_data[15]) );
  MUX2_X1 U3240 ( .A(n4842), .B(n4841), .S(n4858), .Z(wr_data[14]) );
  MUX2_X1 U3241 ( .A(n4844), .B(n4843), .S(n4858), .Z(wr_data[13]) );
  MUX2_X1 U3242 ( .A(n4846), .B(n4845), .S(n4858), .Z(wr_data[12]) );
  MUX2_X1 U3243 ( .A(n4848), .B(n4847), .S(n4858), .Z(wr_data[11]) );
  MUX2_X1 U3244 ( .A(n4850), .B(n4849), .S(n4858), .Z(wr_data[10]) );
  MUX2_X1 U3245 ( .A(n4852), .B(n4851), .S(n4858), .Z(wr_data[0]) );
  INV_X1 U3246 ( .A(n3802), .ZN(\unit_fetch/unit_programCounter/ffi_8/n5 ) );
  AOI21_X1 U3247 ( .B1(\unit_fetch/pc_regout[8] ), .B2(n3803), .A(n4873), .ZN(
        n3802) );
  INV_X1 U3248 ( .A(n3804), .ZN(\unit_fetch/unit_programCounter/ffi_6/n5 ) );
  AOI21_X1 U3249 ( .B1(\unit_fetch/pc_regout[6] ), .B2(n3803), .A(n4871), .ZN(
        n3804) );
  INV_X1 U3250 ( .A(n3805), .ZN(\unit_fetch/unit_programCounter/ffi_4/n5 ) );
  AOI21_X1 U3251 ( .B1(\unit_fetch/pc_regout[4] ), .B2(n3803), .A(n4869), .ZN(
        n3805) );
  OAI21_X1 U3252 ( .B1(n4857), .B2(n4899), .A(n3806), .ZN(
        \unit_fetch/unit_programCounter/ffi_31/n5 ) );
  INV_X1 U3253 ( .A(n4896), .ZN(n3806) );
  INV_X1 U3254 ( .A(n3807), .ZN(\unit_fetch/unit_programCounter/ffi_3/n5 ) );
  AOI21_X1 U3255 ( .B1(\unit_fetch/pc_regout[3] ), .B2(n3803), .A(n4868), .ZN(
        n3807) );
  INV_X1 U3256 ( .A(n3808), .ZN(\unit_fetch/unit_programCounter/ffi_29/n5 ) );
  AOI21_X1 U3257 ( .B1(n3803), .B2(\unit_fetch/pc_regout[29] ), .A(n4894), 
        .ZN(n3808) );
  INV_X1 U3258 ( .A(n3809), .ZN(\unit_fetch/unit_programCounter/ffi_28/n5 ) );
  AOI21_X1 U3259 ( .B1(n3803), .B2(\unit_fetch/pc_regout[28] ), .A(n4893), 
        .ZN(n3809) );
  OAI21_X1 U3260 ( .B1(n4899), .B2(n3793), .A(n3810), .ZN(
        \unit_fetch/unit_programCounter/ffi_26/n5 ) );
  INV_X1 U3261 ( .A(n4891), .ZN(n3810) );
  OAI21_X1 U3262 ( .B1(n4899), .B2(n3782), .A(n3811), .ZN(
        \unit_fetch/unit_programCounter/ffi_24/n5 ) );
  INV_X1 U3263 ( .A(n4889), .ZN(n3811) );
  OAI21_X1 U3264 ( .B1(n4899), .B2(n3775), .A(n3812), .ZN(
        \unit_fetch/unit_programCounter/ffi_22/n5 ) );
  INV_X1 U3265 ( .A(n4887), .ZN(n3812) );
  OAI21_X1 U3266 ( .B1(n4899), .B2(n3792), .A(n3813), .ZN(
        \unit_fetch/unit_programCounter/ffi_20/n5 ) );
  INV_X1 U3267 ( .A(n4885), .ZN(n3813) );
  INV_X1 U3268 ( .A(n3814), .ZN(\unit_fetch/unit_programCounter/ffi_19/n5 ) );
  AOI21_X1 U3269 ( .B1(n3803), .B2(\unit_fetch/pc_regout[19] ), .A(n4884), 
        .ZN(n3814) );
  INV_X1 U3270 ( .A(n3815), .ZN(\unit_fetch/unit_programCounter/ffi_18/n5 ) );
  AOI21_X1 U3271 ( .B1(n3803), .B2(\unit_fetch/pc_regout[18] ), .A(n4883), 
        .ZN(n3815) );
  OAI21_X1 U3272 ( .B1(n4899), .B2(n3774), .A(n3816), .ZN(
        \unit_fetch/unit_programCounter/ffi_16/n5 ) );
  INV_X1 U3273 ( .A(n4881), .ZN(n3816) );
  OAI21_X1 U3274 ( .B1(n4899), .B2(n3783), .A(n3817), .ZN(
        \unit_fetch/unit_programCounter/ffi_14/n5 ) );
  INV_X1 U3275 ( .A(n4879), .ZN(n3817) );
  INV_X1 U3276 ( .A(n3818), .ZN(\unit_fetch/unit_programCounter/ffi_12/n5 ) );
  AOI21_X1 U3277 ( .B1(n3803), .B2(\unit_fetch/pc_regout[12] ), .A(n4877), 
        .ZN(n3818) );
  INV_X1 U3278 ( .A(n4899), .ZN(n3803) );
  OAI21_X1 U3279 ( .B1(n4899), .B2(n3791), .A(n3819), .ZN(
        \unit_fetch/unit_programCounter/ffi_10/n5 ) );
  INV_X1 U3280 ( .A(n4875), .ZN(n3819) );
  OAI21_X1 U3281 ( .B1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .B2(n4899), 
        .A(n3820), .ZN(\unit_fetch/unit_programCounter/ffi_1/n5 ) );
  INV_X1 U3282 ( .A(n4866), .ZN(n3820) );
  OAI21_X1 U3283 ( .B1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n4899), 
        .A(n3821), .ZN(\unit_fetch/unit_programCounter/ffi_0/n5 ) );
  INV_X1 U3284 ( .A(n4865), .ZN(n3821) );
  OAI211_X1 U3285 ( .C1(n3779), .C2(n3822), .A(n3823), .B(n3824), .ZN(
        \unit_fetch/unit_instructionRegister/n98 ) );
  NAND3_X1 U3286 ( .A1(n3825), .A2(n3826), .A3(n3827), .ZN(n3823) );
  OAI221_X1 U3287 ( .B1(n3828), .B2(n3829), .C1(n3830), .C2(n3822), .A(n3824), 
        .ZN(\unit_fetch/unit_instructionRegister/n97 ) );
  OAI221_X1 U3288 ( .B1(n3831), .B2(n3829), .C1(n3832), .C2(n3822), .A(n3824), 
        .ZN(\unit_fetch/unit_instructionRegister/n96 ) );
  OR2_X1 U3289 ( .A1(n3829), .A2(n3833), .ZN(n3824) );
  AOI21_X1 U3290 ( .B1(n3834), .B2(n3835), .A(n3836), .ZN(n3833) );
  INV_X1 U3291 ( .A(n3837), .ZN(n3834) );
  NOR3_X1 U3292 ( .A1(n3838), .A2(n3839), .A3(n3840), .ZN(n3831) );
  OAI21_X1 U3293 ( .B1(\unit_fetch/pc_regout[3] ), .B2(n3841), .A(n3842), .ZN(
        \unit_fetch/unit_instructionRegister/n95 ) );
  OAI21_X1 U3294 ( .B1(n3836), .B2(n3843), .A(n3825), .ZN(n3842) );
  INV_X1 U3295 ( .A(n3844), .ZN(n3843) );
  OAI21_X1 U3296 ( .B1(n3845), .B2(n3830), .A(n3846), .ZN(n3836) );
  INV_X1 U3297 ( .A(n3847), .ZN(\unit_fetch/unit_instructionRegister/n94 ) );
  AOI21_X1 U3298 ( .B1(n3838), .B2(n3825), .A(n2619), .ZN(n3847) );
  OAI22_X1 U3299 ( .A1(n3848), .A2(n3830), .B1(n3849), .B2(n3850), .ZN(n3838)
         );
  AOI21_X1 U3300 ( .B1(n3851), .B2(n3852), .A(n3853), .ZN(n3849) );
  OAI21_X1 U3301 ( .B1(n3822), .B2(n3854), .A(n3855), .ZN(
        \unit_fetch/unit_instructionRegister/n93 ) );
  NAND2_X1 U3302 ( .A1(n3835), .A2(\unit_fetch/pc_regout[3] ), .ZN(n3854) );
  OAI21_X1 U3303 ( .B1(n3828), .B2(n3829), .A(n3856), .ZN(
        \unit_fetch/unit_instructionRegister/n90 ) );
  AOI211_X1 U3304 ( .C1(n3857), .C2(n3827), .A(n3858), .B(n3840), .ZN(n3828)
         );
  INV_X1 U3305 ( .A(n3859), .ZN(n3858) );
  OAI21_X1 U3306 ( .B1(n3860), .B2(n3822), .A(n3856), .ZN(
        \unit_fetch/unit_instructionRegister/n89 ) );
  AOI22_X1 U3307 ( .A1(n3861), .A2(n3862), .B1(n3863), .B2(n3825), .ZN(n3856)
         );
  INV_X1 U3308 ( .A(n3864), .ZN(n3862) );
  OAI22_X1 U3309 ( .A1(n3865), .A2(n3829), .B1(n3866), .B2(n3822), .ZN(
        \unit_fetch/unit_instructionRegister/n88 ) );
  AND2_X1 U3310 ( .A1(n3850), .A2(n3867), .ZN(n3866) );
  NOR4_X1 U3311 ( .A1(n3840), .A2(n3868), .A3(n3869), .A4(n3863), .ZN(n3865)
         );
  OAI21_X1 U3312 ( .B1(n3837), .B2(n3870), .A(n3871), .ZN(n3863) );
  AOI21_X1 U3313 ( .B1(n3871), .B2(n3844), .A(n3829), .ZN(
        \unit_fetch/unit_instructionRegister/n87 ) );
  NOR2_X1 U3314 ( .A1(n3872), .A2(n3873), .ZN(n3844) );
  AOI211_X1 U3315 ( .C1(n3771), .C2(n3853), .A(n3874), .B(n3839), .ZN(n3871)
         );
  INV_X1 U3316 ( .A(n3875), .ZN(\unit_fetch/unit_instructionRegister/n82 ) );
  AOI22_X1 U3317 ( .A1(n3876), .A2(n3825), .B1(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n3861), .ZN(n3875) );
  OAI221_X1 U3318 ( .B1(n3877), .B2(n3829), .C1(n3832), .C2(n3822), .A(n3841), 
        .ZN(\unit_fetch/unit_instructionRegister/n81 ) );
  INV_X1 U3319 ( .A(n3861), .ZN(n3822) );
  INV_X1 U3320 ( .A(n3878), .ZN(n3832) );
  OAI21_X1 U3321 ( .B1(n3879), .B2(n3829), .A(n3841), .ZN(
        \unit_fetch/unit_instructionRegister/n80 ) );
  NAND2_X1 U3322 ( .A1(n3880), .A2(n3861), .ZN(n3841) );
  NOR2_X1 U3323 ( .A1(n3837), .A2(n3829), .ZN(n3861) );
  NOR4_X1 U3324 ( .A1(n3840), .A2(n3874), .A3(n3881), .A4(n3876), .ZN(n3879)
         );
  OAI21_X1 U3325 ( .B1(n3837), .B2(n3850), .A(n3877), .ZN(n3876) );
  NOR2_X1 U3326 ( .A1(n3882), .A2(n3873), .ZN(n3877) );
  AND3_X1 U3327 ( .A1(n3883), .A2(n3773), .A3(n3884), .ZN(n3873) );
  INV_X1 U3328 ( .A(n3835), .ZN(n3850) );
  NOR2_X1 U3329 ( .A1(n3860), .A2(n3771), .ZN(n3835) );
  NOR2_X1 U3330 ( .A1(n3837), .A2(n3885), .ZN(n3840) );
  NOR2_X1 U3331 ( .A1(n3886), .A2(n3829), .ZN(
        \unit_fetch/unit_instructionRegister/n79 ) );
  NOR3_X1 U3332 ( .A1(n3882), .A2(n3839), .A3(n3872), .ZN(n3886) );
  NAND2_X1 U3333 ( .A1(n3859), .A2(n3887), .ZN(n3872) );
  OR3_X1 U3334 ( .A1(n3773), .A2(n3888), .A3(n3837), .ZN(n3887) );
  NAND2_X1 U3335 ( .A1(n3889), .A2(n3773), .ZN(n3859) );
  OAI21_X1 U3336 ( .B1(n3888), .B2(n3845), .A(n3890), .ZN(n3882) );
  NOR2_X1 U3337 ( .A1(n3771), .A2(n3891), .ZN(n3888) );
  NOR2_X1 U3338 ( .A1(n3892), .A2(n3829), .ZN(
        \unit_fetch/unit_instructionRegister/n78 ) );
  OAI21_X1 U3339 ( .B1(n3829), .B2(n3890), .A(n3893), .ZN(
        \unit_fetch/unit_instructionRegister/n77 ) );
  AND2_X1 U3340 ( .A1(n3894), .A2(n3825), .ZN(
        \unit_fetch/unit_instructionRegister/n75 ) );
  AND2_X1 U3341 ( .A1(n3895), .A2(n3825), .ZN(
        \unit_fetch/unit_instructionRegister/n74 ) );
  AND4_X1 U3342 ( .A1(n3896), .A2(n3830), .A3(n3897), .A4(n3825), .ZN(
        \unit_fetch/unit_instructionRegister/n71 ) );
  NAND2_X1 U3343 ( .A1(n3898), .A2(n3825), .ZN(
        \unit_fetch/unit_instructionRegister/n70 ) );
  NOR2_X1 U3344 ( .A1(RST), .A2(n3761), .ZN(
        \unit_control/uut_third_stage/ffi_9/n6 ) );
  NOR2_X1 U3345 ( .A1(RST), .A2(n3760), .ZN(
        \unit_control/uut_third_stage/ffi_4/n5 ) );
  NOR2_X1 U3346 ( .A1(RST), .A2(n3759), .ZN(
        \unit_control/uut_third_stage/ffi_3/n5 ) );
  NOR2_X1 U3347 ( .A1(RST), .A2(n3758), .ZN(
        \unit_control/uut_third_stage/ffi_17/n6 ) );
  NOR2_X1 U3348 ( .A1(RST), .A2(n3757), .ZN(
        \unit_control/uut_third_stage/ffi_14/n5 ) );
  NOR2_X1 U3349 ( .A1(RST), .A2(n3756), .ZN(
        \unit_control/uut_third_stage/ffi_13/n5 ) );
  NOR2_X1 U3350 ( .A1(RST), .A2(n3755), .ZN(
        \unit_control/uut_third_stage/ffi_12/n5 ) );
  NOR2_X1 U3351 ( .A1(RST), .A2(n3754), .ZN(
        \unit_control/uut_third_stage/ffi_10/n5 ) );
  NAND2_X1 U3352 ( .A1(n3899), .A2(n3900), .ZN(
        \unit_control/uut_second_stage/ffi_17/n5 ) );
  OAI21_X1 U3353 ( .B1(n3901), .B2(n3902), .A(n3900), .ZN(
        \unit_control/uut_second_stage/ffi_13/n5 ) );
  OAI21_X1 U3354 ( .B1(n3903), .B2(n3904), .A(n3905), .ZN(
        \unit_control/uut_second_stage/ffi_10/n5 ) );
  INV_X1 U3355 ( .A(\unit_control/uut_second_stage/ffi_12/n5 ), .ZN(n3905) );
  NOR2_X1 U3356 ( .A1(n3898), .A2(\unit_fetch/unit_instructionRegister/n68 ), 
        .ZN(\unit_control/uut_second_stage/ffi_12/n5 ) );
  OR2_X1 U3357 ( .A1(n3906), .A2(n3829), .ZN(
        \unit_fetch/unit_instructionRegister/n68 ) );
  NAND2_X1 U3358 ( .A1(n3907), .A2(n3901), .ZN(n3904) );
  NOR2_X1 U3359 ( .A1(RST), .A2(n3753), .ZN(
        \unit_control/uut_fourth_stage/ffi_4/n5 ) );
  NOR2_X1 U3360 ( .A1(RST), .A2(n3752), .ZN(
        \unit_control/uut_fourth_stage/ffi_3/n6 ) );
  NOR4_X1 U3361 ( .A1(\unit_control/n153 ), .A2(\unit_control/n152 ), .A3(
        n3908), .A4(n3909), .ZN(\unit_control/next_state[1] ) );
  NOR4_X1 U3362 ( .A1(\unit_control/n153 ), .A2(\unit_control/n152 ), .A3(
        n3910), .A4(n3911), .ZN(\unit_control/next_state[0] ) );
  OAI22_X1 U3363 ( .A1(n3912), .A2(n3913), .B1(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n3914), .ZN(n4865) );
  OAI22_X1 U3364 ( .A1(n3915), .A2(n3913), .B1(
        \unit_fetch/unit_programCounter/ffi_1/n4 ), .B2(n3914), .ZN(n4866) );
  OAI22_X1 U3365 ( .A1(n3916), .A2(n3913), .B1(n3917), .B2(n3914), .ZN(n4868)
         );
  XNOR2_X1 U3366 ( .A(\unit_fetch/pc_regout[3] ), .B(\unit_fetch/pc_regout[2] ), .ZN(n3917) );
  OAI21_X1 U3367 ( .B1(n3918), .B2(n3913), .A(n3919), .ZN(n4869) );
  OAI21_X1 U3368 ( .B1(n3897), .B2(n3920), .A(n3921), .ZN(n3919) );
  MUX2_X1 U3369 ( .A(n3922), .B(\unit_fetch/pc_regout[4] ), .S(n3771), .Z(
        n3920) );
  OAI22_X1 U3370 ( .A1(n3923), .A2(n3913), .B1(n3924), .B2(n3914), .ZN(n4871)
         );
  XNOR2_X1 U3371 ( .A(n3925), .B(\unit_fetch/pc_regout[6] ), .ZN(n3924) );
  OAI22_X1 U3372 ( .A1(n3926), .A2(n3913), .B1(n3927), .B2(n3914), .ZN(n4873)
         );
  XNOR2_X1 U3373 ( .A(n3772), .B(n3928), .ZN(n3927) );
  OAI22_X1 U3374 ( .A1(n3929), .A2(n3913), .B1(n3930), .B2(n3914), .ZN(n4875)
         );
  XNOR2_X1 U3375 ( .A(n3931), .B(n3791), .ZN(n3930) );
  OAI22_X1 U3376 ( .A1(n3932), .A2(n3913), .B1(n3933), .B2(n3914), .ZN(n4877)
         );
  XNOR2_X1 U3377 ( .A(\unit_fetch/pc_regout[12] ), .B(n3934), .ZN(n3933) );
  OAI22_X1 U3378 ( .A1(n3935), .A2(n3913), .B1(n3936), .B2(n3914), .ZN(n4879)
         );
  XNOR2_X1 U3379 ( .A(n3937), .B(\unit_fetch/pc_regout[14] ), .ZN(n3936) );
  OAI22_X1 U3380 ( .A1(n3938), .A2(n3913), .B1(n3939), .B2(n3914), .ZN(n4881)
         );
  XNOR2_X1 U3381 ( .A(n3774), .B(n3940), .ZN(n3939) );
  OAI22_X1 U3382 ( .A1(n3941), .A2(n3913), .B1(n3942), .B2(n3914), .ZN(n4883)
         );
  XNOR2_X1 U3383 ( .A(n3943), .B(\unit_fetch/pc_regout[18] ), .ZN(n3942) );
  OAI21_X1 U3384 ( .B1(n3944), .B2(n3913), .A(n3945), .ZN(n4884) );
  NAND3_X1 U3385 ( .A1(n3946), .A2(n3947), .A3(n3921), .ZN(n3945) );
  INV_X1 U3386 ( .A(n3948), .ZN(n3946) );
  AOI21_X1 U3387 ( .B1(n3943), .B2(\unit_fetch/pc_regout[18] ), .A(
        \unit_fetch/pc_regout[19] ), .ZN(n3948) );
  OAI22_X1 U3388 ( .A1(n3949), .A2(n3913), .B1(n3950), .B2(n3914), .ZN(n4885)
         );
  XNOR2_X1 U3389 ( .A(n3792), .B(n3947), .ZN(n3950) );
  OAI22_X1 U3390 ( .A1(n3951), .A2(n3913), .B1(n3952), .B2(n3914), .ZN(n4887)
         );
  XNOR2_X1 U3391 ( .A(n3953), .B(\unit_fetch/pc_regout[22] ), .ZN(n3952) );
  OAI22_X1 U3392 ( .A1(n3954), .A2(n3913), .B1(n3955), .B2(n3914), .ZN(n4889)
         );
  XNOR2_X1 U3393 ( .A(\unit_fetch/pc_regout[24] ), .B(n3956), .ZN(n3955) );
  OAI22_X1 U3394 ( .A1(n3957), .A2(n3913), .B1(n3958), .B2(n3914), .ZN(n4891)
         );
  XNOR2_X1 U3395 ( .A(n3959), .B(n3793), .ZN(n3958) );
  OAI21_X1 U3396 ( .B1(n3960), .B2(n3913), .A(n3961), .ZN(n4893) );
  OAI211_X1 U3397 ( .C1(n3962), .C2(\unit_fetch/pc_regout[28] ), .A(n3963), 
        .B(n3921), .ZN(n3961) );
  AND2_X1 U3398 ( .A1(n3964), .A2(\unit_fetch/pc_regout[27] ), .ZN(n3962) );
  OAI22_X1 U3399 ( .A1(n3965), .A2(n3913), .B1(n3966), .B2(n3914), .ZN(n4894)
         );
  XNOR2_X1 U3400 ( .A(n3967), .B(\unit_fetch/pc_regout[29] ), .ZN(n3966) );
  OAI22_X1 U3401 ( .A1(n3968), .A2(n3913), .B1(n3914), .B2(n3969), .ZN(n4896)
         );
  XOR2_X1 U3402 ( .A(n4857), .B(n3827), .Z(n3969) );
  OAI22_X1 U3403 ( .A1(n3970), .A2(n3913), .B1(\unit_fetch/pc_regout[2] ), 
        .B2(n3914), .ZN(n4867) );
  OAI21_X1 U3404 ( .B1(n3971), .B2(n3913), .A(n3972), .ZN(n4870) );
  OAI211_X1 U3405 ( .C1(n3973), .C2(\unit_fetch/pc_regout[5] ), .A(n3974), .B(
        n3921), .ZN(n3972) );
  NOR3_X1 U3406 ( .A1(n3773), .A2(n3771), .A3(n3789), .ZN(n3973) );
  OAI21_X1 U3407 ( .B1(n3975), .B2(n3913), .A(n3976), .ZN(n4872) );
  NAND3_X1 U3408 ( .A1(n3977), .A2(n3928), .A3(n3921), .ZN(n3976) );
  OAI21_X1 U3409 ( .B1(n3974), .B2(n3797), .A(n3784), .ZN(n3977) );
  INV_X1 U3410 ( .A(n3925), .ZN(n3974) );
  OAI21_X1 U3411 ( .B1(n3978), .B2(n3913), .A(n3979), .ZN(n4874) );
  NAND3_X1 U3412 ( .A1(n3980), .A2(n3931), .A3(n3921), .ZN(n3979) );
  OAI21_X1 U3413 ( .B1(n3772), .B2(n3928), .A(n3777), .ZN(n3980) );
  OAI21_X1 U3414 ( .B1(n3981), .B2(n3913), .A(n3982), .ZN(n4876) );
  NAND3_X1 U3415 ( .A1(n3983), .A2(n3984), .A3(n3921), .ZN(n3982) );
  INV_X1 U3416 ( .A(n3934), .ZN(n3984) );
  OAI21_X1 U3417 ( .B1(n3931), .B2(n3791), .A(n4854), .ZN(n3983) );
  OAI21_X1 U3418 ( .B1(n3985), .B2(n3913), .A(n3986), .ZN(n4878) );
  OR3_X1 U3419 ( .A1(n3987), .A2(n3937), .A3(n3914), .ZN(n3986) );
  AOI21_X1 U3420 ( .B1(n3934), .B2(\unit_fetch/pc_regout[12] ), .A(
        \unit_fetch/pc_regout[13] ), .ZN(n3987) );
  OAI21_X1 U3421 ( .B1(n3988), .B2(n3913), .A(n3989), .ZN(n4880) );
  NAND3_X1 U3422 ( .A1(n3990), .A2(n3940), .A3(n3921), .ZN(n3989) );
  OAI21_X1 U3423 ( .B1(n3991), .B2(n3783), .A(n3796), .ZN(n3990) );
  OAI21_X1 U3424 ( .B1(n3992), .B2(n3913), .A(n3993), .ZN(n4882) );
  NAND3_X1 U3425 ( .A1(n3994), .A2(n3995), .A3(n3921), .ZN(n3993) );
  INV_X1 U3426 ( .A(n3943), .ZN(n3995) );
  OAI21_X1 U3427 ( .B1(n3940), .B2(n3774), .A(n4855), .ZN(n3994) );
  OAI21_X1 U3428 ( .B1(n3996), .B2(n3913), .A(n3997), .ZN(n4886) );
  NAND3_X1 U3429 ( .A1(n3998), .A2(n3999), .A3(n3921), .ZN(n3997) );
  OAI21_X1 U3430 ( .B1(n3947), .B2(n3792), .A(n4856), .ZN(n3998) );
  OAI21_X1 U3431 ( .B1(n4000), .B2(n3913), .A(n4001), .ZN(n4888) );
  NAND3_X1 U3432 ( .A1(n4002), .A2(n4003), .A3(n3921), .ZN(n4001) );
  OAI21_X1 U3433 ( .B1(n3999), .B2(n3775), .A(n3794), .ZN(n4002) );
  OAI21_X1 U3434 ( .B1(n4004), .B2(n3913), .A(n4005), .ZN(n4890) );
  OAI211_X1 U3435 ( .C1(n4006), .C2(\unit_fetch/pc_regout[25] ), .A(n3959), 
        .B(n3921), .ZN(n4005) );
  NOR2_X1 U3436 ( .A1(n4003), .A2(n3782), .ZN(n4006) );
  INV_X1 U3437 ( .A(n3956), .ZN(n4003) );
  OAI22_X1 U3438 ( .A1(n4007), .A2(n3913), .B1(n4008), .B2(n3914), .ZN(n4892)
         );
  XNOR2_X1 U3439 ( .A(\unit_fetch/pc_regout[27] ), .B(n3964), .ZN(n4008) );
  OAI21_X1 U3440 ( .B1(n4009), .B2(n3913), .A(n4010), .ZN(n4895) );
  OR3_X1 U3441 ( .A1(n4011), .A2(n3827), .A3(n3914), .ZN(n4010) );
  INV_X1 U3442 ( .A(n3921), .ZN(n3914) );
  AND3_X1 U3443 ( .A1(\unit_fetch/pc_regout[29] ), .A2(n3967), .A3(
        \unit_fetch/pc_regout[30] ), .ZN(n3827) );
  AOI21_X1 U3444 ( .B1(n3967), .B2(\unit_fetch/pc_regout[29] ), .A(
        \unit_fetch/pc_regout[30] ), .ZN(n4011) );
  INV_X1 U3445 ( .A(n3963), .ZN(n3967) );
  NAND3_X1 U3446 ( .A1(\unit_fetch/pc_regout[27] ), .A2(n3964), .A3(
        \unit_fetch/pc_regout[28] ), .ZN(n3963) );
  NOR2_X1 U3447 ( .A1(n3793), .A2(n3959), .ZN(n3964) );
  NAND3_X1 U3448 ( .A1(\unit_fetch/pc_regout[24] ), .A2(n3956), .A3(
        \unit_fetch/pc_regout[25] ), .ZN(n3959) );
  NOR3_X1 U3449 ( .A1(n3775), .A2(n3999), .A3(n3794), .ZN(n3956) );
  INV_X1 U3450 ( .A(n3953), .ZN(n3999) );
  NOR3_X1 U3451 ( .A1(n3947), .A2(n4856), .A3(n3792), .ZN(n3953) );
  NAND3_X1 U3452 ( .A1(\unit_fetch/pc_regout[18] ), .A2(n3943), .A3(
        \unit_fetch/pc_regout[19] ), .ZN(n3947) );
  NOR3_X1 U3453 ( .A1(n3940), .A2(n4855), .A3(n3774), .ZN(n3943) );
  NAND3_X1 U3454 ( .A1(\unit_fetch/pc_regout[14] ), .A2(n3937), .A3(
        \unit_fetch/pc_regout[15] ), .ZN(n3940) );
  INV_X1 U3455 ( .A(n3991), .ZN(n3937) );
  NAND3_X1 U3456 ( .A1(\unit_fetch/pc_regout[12] ), .A2(n3934), .A3(
        \unit_fetch/pc_regout[13] ), .ZN(n3991) );
  NOR3_X1 U3457 ( .A1(n3931), .A2(n4854), .A3(n3791), .ZN(n3934) );
  OR3_X1 U3458 ( .A1(n3928), .A2(n3772), .A3(n3777), .ZN(n3931) );
  NAND3_X1 U3459 ( .A1(\unit_fetch/pc_regout[6] ), .A2(n3925), .A3(
        \unit_fetch/pc_regout[7] ), .ZN(n3928) );
  NOR4_X1 U3460 ( .A1(n3780), .A2(n3773), .A3(n3789), .A4(n3771), .ZN(n3925)
         );
  NAND2_X1 U3461 ( .A1(n4013), .A2(n2912), .ZN(n4899) );
  NOR2_X1 U3462 ( .A1(\unit_decode/RD1reg/ffi_0/n4 ), .A2(RST), .ZN(n4900) );
  NOR2_X1 U3463 ( .A1(\unit_decode/RD1reg/ffi_1/n4 ), .A2(RST), .ZN(n4901) );
  NOR2_X1 U3464 ( .A1(\unit_decode/RD1reg/ffi_2/n4 ), .A2(RST), .ZN(n4902) );
  NOR2_X1 U3465 ( .A1(\unit_decode/RD1reg/ffi_3/n4 ), .A2(RST), .ZN(n4903) );
  NOR2_X1 U3466 ( .A1(\unit_decode/RD1reg/ffi_4/n4 ), .A2(RST), .ZN(n4904) );
  NOR2_X1 U3467 ( .A1(RST), .A2(n3912), .ZN(n4905) );
  AND3_X1 U3468 ( .A1(n4014), .A2(n4015), .A3(n4016), .ZN(n3912) );
  AOI211_X1 U3469 ( .C1(n4017), .C2(n4018), .A(n4019), .B(n4020), .ZN(n4016)
         );
  MUX2_X1 U3470 ( .A(n4021), .B(n4022), .S(n4023), .Z(n4020) );
  NOR2_X1 U3471 ( .A1(n3786), .A2(n4024), .ZN(n4022) );
  OAI21_X1 U3472 ( .B1(\unit_decode/IMMreg/ffi_0/n4 ), .B2(n4025), .A(n4026), 
        .ZN(n4021) );
  INV_X1 U3473 ( .A(n4027), .ZN(n4019) );
  AOI222_X1 U3474 ( .A1(n4028), .A2(n4029), .B1(n4030), .B2(n4031), .C1(n4032), 
        .C2(n4033), .ZN(n4027) );
  AOI221_X1 U3475 ( .B1(n4034), .B2(n3785), .C1(n4035), .C2(n4036), .A(n4037), 
        .ZN(n4015) );
  AOI211_X1 U3476 ( .C1(n4038), .C2(n4039), .A(n3795), .B(n4859), .ZN(n4037)
         );
  OR2_X1 U3477 ( .A1(n4040), .A2(n4861), .ZN(n4039) );
  MUX2_X1 U3478 ( .A(n4041), .B(n4042), .S(n4853), .Z(n4038) );
  NAND2_X1 U3479 ( .A1(n4861), .A2(n4040), .ZN(n4042) );
  NAND4_X1 U3480 ( .A1(n4043), .A2(n4044), .A3(n4045), .A4(n4046), .ZN(n4040)
         );
  NOR4_X1 U3481 ( .A1(n4047), .A2(n4048), .A3(n4049), .A4(n4050), .ZN(n4046)
         );
  OR4_X1 U3482 ( .A1(n4051), .A2(n4052), .A3(n4053), .A4(n4054), .ZN(n4050) );
  OR4_X1 U3483 ( .A1(n4055), .A2(n4056), .A3(n4057), .A4(n4058), .ZN(n4049) );
  OR4_X1 U3484 ( .A1(n4059), .A2(n4060), .A3(n4061), .A4(n4062), .ZN(n4048) );
  OR4_X1 U3485 ( .A1(n4063), .A2(n4064), .A3(n4065), .A4(n4066), .ZN(n4047) );
  NOR4_X1 U3486 ( .A1(n4067), .A2(n4068), .A3(n4069), .A4(n4070), .ZN(n4045)
         );
  NAND3_X1 U3487 ( .A1(n4071), .A2(n4072), .A3(n4073), .ZN(n4068) );
  NAND4_X1 U3488 ( .A1(n4074), .A2(n4075), .A3(n4076), .A4(n4077), .ZN(n4067)
         );
  INV_X1 U3489 ( .A(n4078), .ZN(n4074) );
  NOR4_X1 U3490 ( .A1(n4079), .A2(n4080), .A3(n4081), .A4(n4082), .ZN(n4044)
         );
  NOR4_X1 U3491 ( .A1(n4083), .A2(n4084), .A3(n4085), .A4(n4086), .ZN(n4043)
         );
  XOR2_X1 U3492 ( .A(n4087), .B(\unit_decode/IMMreg/ffi_31/n4 ), .Z(n4041) );
  MUX2_X1 U3493 ( .A(n4088), .B(n4089), .S(n4090), .Z(n4087) );
  NOR2_X1 U3494 ( .A1(n4091), .A2(n4092), .ZN(n4090) );
  NOR4_X1 U3495 ( .A1(n4093), .A2(n4094), .A3(n4095), .A4(n4096), .ZN(n4091)
         );
  OR2_X1 U3496 ( .A1(n4097), .A2(n4098), .ZN(n4089) );
  NAND2_X1 U3497 ( .A1(n4097), .A2(n4099), .ZN(n4088) );
  OAI222_X1 U3498 ( .A1(n4100), .A2(n4101), .B1(n4102), .B2(n4103), .C1(n4104), 
        .C2(n4105), .ZN(n4034) );
  AOI22_X1 U3499 ( .A1(n4106), .A2(n4052), .B1(n4107), .B2(n4108), .ZN(n4014)
         );
  OAI21_X1 U3500 ( .B1(n4023), .B2(n3786), .A(n4109), .ZN(n4052) );
  NOR2_X1 U3501 ( .A1(RST), .A2(n3970), .ZN(n4906) );
  AND4_X1 U3502 ( .A1(n4110), .A2(n4111), .A3(n4112), .A4(n4113), .ZN(n3970)
         );
  AOI221_X1 U3503 ( .B1(n4017), .B2(n4114), .C1(n4058), .C2(n4106), .A(n4115), 
        .ZN(n4113) );
  NOR3_X1 U3504 ( .A1(n4101), .A2(n4862), .A3(n4104), .ZN(n4115) );
  XOR2_X1 U3505 ( .A(n4116), .B(n4117), .Z(n4058) );
  AOI222_X1 U3506 ( .A1(n4031), .A2(n4032), .B1(n4029), .B2(n4118), .C1(n4108), 
        .C2(n4018), .ZN(n4112) );
  AOI21_X1 U3507 ( .B1(n4121), .B2(n4122), .A(n4123), .ZN(n4110) );
  MUX2_X1 U3508 ( .A(n4124), .B(n4125), .S(n3790), .Z(n4123) );
  MUX2_X1 U3509 ( .A(n4126), .B(n4036), .S(n4102), .Z(n4125) );
  NOR2_X1 U3510 ( .A1(n4122), .A2(n4024), .ZN(n4124) );
  NOR2_X1 U3511 ( .A1(RST), .A2(n3916), .ZN(n4907) );
  AOI221_X1 U3512 ( .B1(n4106), .B2(n4082), .C1(n4127), .C2(n4128), .A(n4129), 
        .ZN(n3916) );
  INV_X1 U3513 ( .A(n4130), .ZN(n4129) );
  MUX2_X1 U3514 ( .A(n4131), .B(n4132), .S(n3778), .Z(n4130) );
  MUX2_X1 U3515 ( .A(n4025), .B(n4133), .S(n4104), .Z(n4132) );
  NAND2_X1 U3516 ( .A1(n4134), .A2(n4104), .ZN(n4131) );
  OR4_X1 U3517 ( .A1(n4135), .A2(n4136), .A3(n4137), .A4(n4138), .ZN(n4127) );
  OAI22_X1 U3518 ( .A1(n4139), .A2(n4140), .B1(n4141), .B2(n4142), .ZN(n4138)
         );
  OAI22_X1 U3519 ( .A1(n4143), .A2(n4144), .B1(n4145), .B2(n4146), .ZN(n4137)
         );
  OAI22_X1 U3520 ( .A1(n4147), .A2(n4148), .B1(n4104), .B2(n4149), .ZN(n4136)
         );
  OAI222_X1 U3521 ( .A1(n4150), .A2(n4151), .B1(n4152), .B2(n4153), .C1(n4154), 
        .C2(n4155), .ZN(n4135) );
  XNOR2_X1 U3522 ( .A(n4156), .B(n4104), .ZN(n4082) );
  XOR2_X1 U3523 ( .A(n4157), .B(n4158), .Z(n4156) );
  NOR2_X1 U3524 ( .A1(RST), .A2(n3918), .ZN(n4908) );
  AND4_X1 U3525 ( .A1(n4159), .A2(n4160), .A3(n4161), .A4(n4162), .ZN(n3918)
         );
  AOI221_X1 U3526 ( .B1(n4080), .B2(n4106), .C1(n4163), .C2(n3787), .A(n4164), 
        .ZN(n4162) );
  NOR3_X1 U3527 ( .A1(n4165), .A2(n4166), .A3(n4167), .ZN(n4164) );
  MUX2_X1 U3528 ( .A(n4126), .B(n4036), .S(n4168), .Z(n4163) );
  MUX2_X1 U3529 ( .A(n4169), .B(n4170), .S(n4171), .Z(n4080) );
  NOR2_X1 U3530 ( .A1(n4172), .A2(n4173), .ZN(n4170) );
  XNOR2_X1 U3531 ( .A(n4174), .B(n4168), .ZN(n4169) );
  AOI222_X1 U3532 ( .A1(n4017), .A2(n4175), .B1(n4108), .B2(n4114), .C1(n4030), 
        .C2(n4176), .ZN(n4161) );
  AOI222_X1 U3533 ( .A1(n4107), .A2(n4118), .B1(n4033), .B2(n4177), .C1(n4029), 
        .C2(n4121), .ZN(n4160) );
  AOI222_X1 U3534 ( .A1(n4032), .A2(n4119), .B1(n4031), .B2(n4120), .C1(n4028), 
        .C2(n4018), .ZN(n4159) );
  NOR2_X1 U3535 ( .A1(RST), .A2(n3971), .ZN(n4909) );
  AOI221_X1 U3536 ( .B1(n4056), .B2(n4106), .C1(n4178), .C2(n4128), .A(n4179), 
        .ZN(n3971) );
  INV_X1 U3537 ( .A(n4180), .ZN(n4179) );
  MUX2_X1 U3538 ( .A(n4181), .B(n4182), .S(\unit_decode/IMMreg/ffi_5/n4 ), .Z(
        n4180) );
  NAND2_X1 U3539 ( .A1(n4134), .A2(n4183), .ZN(n4182) );
  MUX2_X1 U3540 ( .A(n4025), .B(n4133), .S(n4183), .Z(n4181) );
  OR4_X1 U3541 ( .A1(n4184), .A2(n4185), .A3(n4186), .A4(n4187), .ZN(n4178) );
  OAI22_X1 U3542 ( .A1(n4141), .A2(n4139), .B1(n4145), .B2(n4143), .ZN(n4187)
         );
  OAI22_X1 U3543 ( .A1(n4147), .A2(n4144), .B1(n4149), .B2(n4148), .ZN(n4186)
         );
  INV_X1 U3544 ( .A(n4033), .ZN(n4148) );
  OAI22_X1 U3545 ( .A1(n4154), .A2(n4140), .B1(n4188), .B2(n4151), .ZN(n4185)
         );
  OAI222_X1 U3546 ( .A1(n4150), .A2(n4146), .B1(n4152), .B2(n4142), .C1(n4189), 
        .C2(n4153), .ZN(n4184) );
  XOR2_X1 U3547 ( .A(n4190), .B(n4191), .Z(n4056) );
  NOR2_X1 U3548 ( .A1(RST), .A2(n3923), .ZN(n4910) );
  INV_X1 U3549 ( .A(n4192), .ZN(n3923) );
  OAI211_X1 U3550 ( .C1(n4193), .C2(n4073), .A(n4194), .B(n4195), .ZN(n4192)
         );
  MUX2_X1 U3551 ( .A(n4196), .B(n4197), .S(\unit_decode/IMMreg/ffi_6/n4 ), .Z(
        n4195) );
  NAND2_X1 U3552 ( .A1(n4134), .A2(n4198), .ZN(n4197) );
  MUX2_X1 U3553 ( .A(n4025), .B(n4133), .S(n4198), .Z(n4196) );
  OAI21_X1 U3554 ( .B1(n4199), .B2(n4200), .A(n4128), .ZN(n4194) );
  INV_X1 U3555 ( .A(n4201), .ZN(n4128) );
  OAI221_X1 U3556 ( .B1(n4154), .B2(n4144), .C1(n4149), .C2(n4140), .A(n4202), 
        .ZN(n4200) );
  INV_X1 U3557 ( .A(n4203), .ZN(n4202) );
  OAI22_X1 U3558 ( .A1(n4147), .A2(n4141), .B1(n4139), .B2(n4145), .ZN(n4203)
         );
  INV_X1 U3559 ( .A(n4107), .ZN(n4140) );
  OAI221_X1 U3560 ( .B1(n4188), .B2(n4153), .C1(n4204), .C2(n4151), .A(n4205), 
        .ZN(n4199) );
  INV_X1 U3561 ( .A(n4206), .ZN(n4205) );
  OAI222_X1 U3562 ( .A1(n4146), .A2(n4189), .B1(n4143), .B2(n4152), .C1(n4142), 
        .C2(n4150), .ZN(n4206) );
  INV_X1 U3563 ( .A(n4175), .ZN(n4189) );
  NAND2_X1 U3564 ( .A1(n4207), .A2(n4208), .ZN(n4073) );
  NAND3_X1 U3565 ( .A1(n4209), .A2(n4210), .A3(n4211), .ZN(n4208) );
  INV_X1 U3566 ( .A(n4212), .ZN(n4207) );
  NOR2_X1 U3567 ( .A1(RST), .A2(n3975), .ZN(n4911) );
  AND3_X1 U3568 ( .A1(n4213), .A2(n4214), .A3(n4215), .ZN(n3975) );
  AOI211_X1 U3569 ( .C1(n4118), .C2(n4119), .A(n4216), .B(n4217), .ZN(n4215)
         );
  MUX2_X1 U3570 ( .A(n4218), .B(n4219), .S(\unit_decode/IMMreg/ffi_7/n4 ), .Z(
        n4217) );
  NOR2_X1 U3571 ( .A1(n4220), .A2(n4024), .ZN(n4219) );
  MUX2_X1 U3572 ( .A(n4126), .B(n4036), .S(n4221), .Z(n4218) );
  OAI222_X1 U3573 ( .A1(n4141), .A2(n4101), .B1(n4222), .B2(n4223), .C1(n4026), 
        .C2(n4144), .ZN(n4216) );
  INV_X1 U3574 ( .A(n4031), .ZN(n4144) );
  INV_X1 U3575 ( .A(n4018), .ZN(n4141) );
  AOI222_X1 U3576 ( .A1(n4028), .A2(n4176), .B1(n4057), .B2(n4106), .C1(n4120), 
        .C2(n4114), .ZN(n4214) );
  XNOR2_X1 U3577 ( .A(n4220), .B(n4224), .ZN(n4057) );
  XNOR2_X1 U3578 ( .A(n4225), .B(n4226), .ZN(n4224) );
  AOI222_X1 U3579 ( .A1(n4030), .A2(n4227), .B1(n4032), .B2(n4175), .C1(n4108), 
        .C2(n4228), .ZN(n4213) );
  NOR2_X1 U3580 ( .A1(RST), .A2(n3926), .ZN(n4912) );
  AND3_X1 U3581 ( .A1(n4229), .A2(n4230), .A3(n4231), .ZN(n3926) );
  AOI211_X1 U3582 ( .C1(n4121), .C2(n4018), .A(n4232), .B(n4233), .ZN(n4231)
         );
  MUX2_X1 U3583 ( .A(n4234), .B(n4235), .S(\unit_decode/IMMreg/ffi_8/n4 ), .Z(
        n4233) );
  NOR2_X1 U3584 ( .A1(n4236), .A2(n4024), .ZN(n4235) );
  MUX2_X1 U3585 ( .A(n4126), .B(n4036), .S(n4237), .Z(n4234) );
  OAI222_X1 U3586 ( .A1(n4238), .A2(n4223), .B1(n4222), .B2(n4239), .C1(n4145), 
        .C2(n4101), .ZN(n4232) );
  INV_X1 U3587 ( .A(n4017), .ZN(n4223) );
  INV_X1 U3588 ( .A(n4240), .ZN(n4230) );
  OAI222_X1 U3589 ( .A1(n4105), .A2(n4150), .B1(n4193), .B2(n4071), .C1(n4103), 
        .C2(n4152), .ZN(n4240) );
  INV_X1 U3590 ( .A(n4114), .ZN(n4152) );
  OAI21_X1 U3591 ( .B1(n4241), .B2(n4242), .A(n4243), .ZN(n4071) );
  INV_X1 U3592 ( .A(n4176), .ZN(n4150) );
  AOI222_X1 U3593 ( .A1(n4108), .A2(n4227), .B1(n4028), .B2(n4175), .C1(n4032), 
        .C2(n4228), .ZN(n4229) );
  NOR2_X1 U3594 ( .A1(RST), .A2(n3978), .ZN(n4913) );
  AND3_X1 U3595 ( .A1(n4244), .A2(n4245), .A3(n4246), .ZN(n3978) );
  AOI211_X1 U3596 ( .C1(n4028), .C2(n4228), .A(n4247), .B(n4248), .ZN(n4246)
         );
  MUX2_X1 U3597 ( .A(n4249), .B(n4250), .S(\unit_decode/IMMreg/ffi_9/n4 ), .Z(
        n4248) );
  NOR2_X1 U3598 ( .A1(n4251), .A2(n4024), .ZN(n4250) );
  MUX2_X1 U3599 ( .A(n4126), .B(n4036), .S(n4252), .Z(n4249) );
  OAI222_X1 U3600 ( .A1(n4204), .A2(n4253), .B1(n4145), .B2(n4026), .C1(n4222), 
        .C2(n4254), .ZN(n4247) );
  INV_X1 U3601 ( .A(n4119), .ZN(n4145) );
  INV_X1 U3602 ( .A(n4227), .ZN(n4204) );
  AOI222_X1 U3603 ( .A1(n4118), .A2(n4176), .B1(n4120), .B2(n4175), .C1(n4062), 
        .C2(n4106), .ZN(n4245) );
  XOR2_X1 U3604 ( .A(n4255), .B(n4256), .Z(n4062) );
  AOI222_X1 U3605 ( .A1(n4177), .A2(n4114), .B1(n4017), .B2(n4257), .C1(n4030), 
        .C2(n4258), .ZN(n4244) );
  NOR2_X1 U3606 ( .A1(RST), .A2(n3929), .ZN(n4914) );
  AND3_X1 U3607 ( .A1(n4259), .A2(n4260), .A3(n4261), .ZN(n3929) );
  AOI211_X1 U3608 ( .C1(n4017), .C2(n4262), .A(n4263), .B(n4264), .ZN(n4261)
         );
  MUX2_X1 U3609 ( .A(n4265), .B(n4266), .S(\unit_decode/IMMreg/ffi_10/n4 ), 
        .Z(n4264) );
  NOR2_X1 U3610 ( .A1(n4267), .A2(n4024), .ZN(n4266) );
  MUX2_X1 U3611 ( .A(n4126), .B(n4036), .S(n4268), .Z(n4265) );
  OAI222_X1 U3612 ( .A1(n4238), .A2(n4254), .B1(n4222), .B2(n4253), .C1(n4269), 
        .C2(n4239), .ZN(n4263) );
  INV_X1 U3613 ( .A(n4270), .ZN(n4222) );
  AOI222_X1 U3614 ( .A1(n4177), .A2(n4176), .B1(n4086), .B2(n4106), .C1(n4121), 
        .C2(n4114), .ZN(n4260) );
  OAI221_X1 U3615 ( .B1(n4271), .B2(n4268), .C1(n4102), .C2(n4272), .A(n4273), 
        .ZN(n4114) );
  XOR2_X1 U3616 ( .A(n4274), .B(n4275), .Z(n4086) );
  AOI222_X1 U3617 ( .A1(n4028), .A2(n4227), .B1(n4118), .B2(n4175), .C1(n4120), 
        .C2(n4228), .ZN(n4259) );
  NOR2_X1 U3618 ( .A1(RST), .A2(n3981), .ZN(n4915) );
  AND3_X1 U3619 ( .A1(n4276), .A2(n4277), .A3(n4278), .ZN(n3981) );
  AOI211_X1 U3620 ( .C1(n4017), .C2(n4279), .A(n4280), .B(n4281), .ZN(n4278)
         );
  MUX2_X1 U3621 ( .A(n4282), .B(n4283), .S(\unit_decode/IMMreg/ffi_11/n4 ), 
        .Z(n4281) );
  NOR2_X1 U3622 ( .A1(n4284), .A2(n4024), .ZN(n4283) );
  MUX2_X1 U3623 ( .A(n4126), .B(n4036), .S(n4285), .Z(n4282) );
  OAI222_X1 U3624 ( .A1(n4269), .A2(n4254), .B1(n4238), .B2(n4253), .C1(n4286), 
        .C2(n4239), .ZN(n4280) );
  AOI222_X1 U3625 ( .A1(n4177), .A2(n4175), .B1(n4121), .B2(n4176), .C1(n4059), 
        .C2(n4106), .ZN(n4277) );
  XOR2_X1 U3626 ( .A(n4287), .B(n4288), .Z(n4059) );
  AOI21_X1 U3627 ( .B1(n4275), .B2(n4274), .A(n4289), .ZN(n4288) );
  OAI211_X1 U3628 ( .C1(n4256), .C2(n4290), .A(n4291), .B(n4292), .ZN(n4274)
         );
  OAI211_X1 U3629 ( .C1(n4293), .C2(n4236), .A(n4242), .B(n4294), .ZN(n4291)
         );
  INV_X1 U3630 ( .A(n4256), .ZN(n4294) );
  OAI221_X1 U3631 ( .B1(n4271), .B2(n4285), .C1(n4104), .C2(n4272), .A(n4273), 
        .ZN(n4176) );
  AOI222_X1 U3632 ( .A1(n4028), .A2(n4270), .B1(n4118), .B2(n4228), .C1(n4120), 
        .C2(n4227), .ZN(n4276) );
  NOR2_X1 U3633 ( .A1(RST), .A2(n3932), .ZN(n4916) );
  AND3_X1 U3634 ( .A1(n4295), .A2(n4296), .A3(n4297), .ZN(n3932) );
  AOI211_X1 U3635 ( .C1(n4017), .C2(n4298), .A(n4299), .B(n4300), .ZN(n4297)
         );
  MUX2_X1 U3636 ( .A(n4301), .B(n4302), .S(\unit_decode/IMMreg/ffi_12/n4 ), 
        .Z(n4300) );
  NOR2_X1 U3637 ( .A1(n4303), .A2(n4024), .ZN(n4302) );
  MUX2_X1 U3638 ( .A(n4126), .B(n4036), .S(n4304), .Z(n4301) );
  OAI222_X1 U3639 ( .A1(n4286), .A2(n4254), .B1(n4269), .B2(n4253), .C1(n4305), 
        .C2(n4239), .ZN(n4299) );
  AOI222_X1 U3640 ( .A1(n4177), .A2(n4228), .B1(n4085), .B2(n4106), .C1(n4121), 
        .C2(n4175), .ZN(n4296) );
  OAI221_X1 U3641 ( .B1(n4271), .B2(n4304), .C1(n4168), .C2(n4272), .A(n4273), 
        .ZN(n4175) );
  XNOR2_X1 U3642 ( .A(n4306), .B(n4307), .ZN(n4085) );
  AOI222_X1 U3643 ( .A1(n4028), .A2(n4258), .B1(n4118), .B2(n4227), .C1(n4120), 
        .C2(n4270), .ZN(n4295) );
  NOR2_X1 U3644 ( .A1(RST), .A2(n3985), .ZN(n4917) );
  AND3_X1 U3645 ( .A1(n4308), .A2(n4309), .A3(n4310), .ZN(n3985) );
  AOI211_X1 U3646 ( .C1(n4028), .C2(n4257), .A(n4311), .B(n4312), .ZN(n4310)
         );
  MUX2_X1 U3647 ( .A(n4313), .B(n4314), .S(\unit_decode/IMMreg/ffi_13/n4 ), 
        .Z(n4312) );
  NOR2_X1 U3648 ( .A1(n4315), .A2(n4024), .ZN(n4314) );
  MUX2_X1 U3649 ( .A(n4126), .B(n4036), .S(n4316), .Z(n4313) );
  OAI222_X1 U3650 ( .A1(n4305), .A2(n4254), .B1(n4286), .B2(n4253), .C1(n4188), 
        .C2(n4026), .ZN(n4311) );
  INV_X1 U3651 ( .A(n4228), .ZN(n4188) );
  OAI221_X1 U3652 ( .B1(n4271), .B2(n4316), .C1(n4183), .C2(n4272), .A(n4273), 
        .ZN(n4228) );
  AOI222_X1 U3653 ( .A1(n4118), .A2(n4270), .B1(n4120), .B2(n4258), .C1(n4060), 
        .C2(n4106), .ZN(n4309) );
  XNOR2_X1 U3654 ( .A(n4317), .B(n4318), .ZN(n4060) );
  OAI21_X1 U3655 ( .B1(n4319), .B2(n4306), .A(n4320), .ZN(n4317) );
  AOI222_X1 U3656 ( .A1(n4177), .A2(n4227), .B1(n4017), .B2(n4321), .C1(n4030), 
        .C2(n4298), .ZN(n4308) );
  NOR2_X1 U3657 ( .A1(RST), .A2(n3935), .ZN(n4918) );
  AND3_X1 U3658 ( .A1(n4322), .A2(n4323), .A3(n4324), .ZN(n3935) );
  AOI211_X1 U3659 ( .C1(n4017), .C2(n4325), .A(n4326), .B(n4327), .ZN(n4324)
         );
  MUX2_X1 U3660 ( .A(n4328), .B(n4329), .S(\unit_decode/IMMreg/ffi_14/n4 ), 
        .Z(n4327) );
  NOR2_X1 U3661 ( .A1(n4330), .A2(n4024), .ZN(n4329) );
  MUX2_X1 U3662 ( .A(n4126), .B(n4036), .S(n4331), .Z(n4328) );
  OAI222_X1 U3663 ( .A1(n4332), .A2(n4254), .B1(n4305), .B2(n4253), .C1(n4333), 
        .C2(n4239), .ZN(n4326) );
  INV_X1 U3664 ( .A(n4279), .ZN(n4305) );
  AOI222_X1 U3665 ( .A1(n4177), .A2(n4270), .B1(n4121), .B2(n4227), .C1(n4106), 
        .C2(n4055), .ZN(n4323) );
  INV_X1 U3666 ( .A(n4334), .ZN(n4055) );
  MUX2_X1 U3667 ( .A(n4335), .B(n4336), .S(n4337), .Z(n4334) );
  OAI21_X1 U3668 ( .B1(n4338), .B2(n4307), .A(n4339), .ZN(n4336) );
  NAND2_X1 U3669 ( .A1(n4340), .A2(n4341), .ZN(n4335) );
  OAI221_X1 U3670 ( .B1(n4271), .B2(n4331), .C1(n4198), .C2(n4272), .A(n4273), 
        .ZN(n4227) );
  AOI222_X1 U3671 ( .A1(n4028), .A2(n4262), .B1(n4118), .B2(n4258), .C1(n4120), 
        .C2(n4257), .ZN(n4322) );
  NOR2_X1 U3672 ( .A1(RST), .A2(n3988), .ZN(n4919) );
  AND3_X1 U3673 ( .A1(n4342), .A2(n4343), .A3(n4344), .ZN(n3988) );
  AOI211_X1 U3674 ( .C1(n4017), .C2(n4345), .A(n4346), .B(n4347), .ZN(n4344)
         );
  MUX2_X1 U3675 ( .A(n4348), .B(n4349), .S(\unit_decode/IMMreg/ffi_15/n4 ), 
        .Z(n4347) );
  NOR2_X1 U3676 ( .A1(n4350), .A2(n4024), .ZN(n4349) );
  MUX2_X1 U3677 ( .A(n4126), .B(n4036), .S(n4351), .Z(n4348) );
  OAI222_X1 U3678 ( .A1(n4333), .A2(n4254), .B1(n4332), .B2(n4253), .C1(n4352), 
        .C2(n4239), .ZN(n4346) );
  INV_X1 U3679 ( .A(n4298), .ZN(n4332) );
  AOI222_X1 U3680 ( .A1(n4177), .A2(n4258), .B1(n4061), .B2(n4106), .C1(n4121), 
        .C2(n4270), .ZN(n4343) );
  OAI221_X1 U3681 ( .B1(n4271), .B2(n4351), .C1(n4221), .C2(n4272), .A(n4273), 
        .ZN(n4270) );
  XOR2_X1 U3682 ( .A(n4353), .B(n4354), .Z(n4061) );
  OAI21_X1 U3683 ( .B1(n4341), .B2(n4337), .A(n4355), .ZN(n4354) );
  INV_X1 U3684 ( .A(n4356), .ZN(n4355) );
  NAND2_X1 U3685 ( .A1(n4307), .A2(n4339), .ZN(n4341) );
  OAI21_X1 U3686 ( .B1(n4357), .B2(n4318), .A(n4358), .ZN(n4339) );
  NOR2_X1 U3687 ( .A1(n4359), .A2(n4303), .ZN(n4357) );
  AOI222_X1 U3688 ( .A1(n4028), .A2(n4279), .B1(n4118), .B2(n4257), .C1(n4120), 
        .C2(n4262), .ZN(n4342) );
  NOR2_X1 U3689 ( .A1(RST), .A2(n3938), .ZN(n4920) );
  AND3_X1 U3690 ( .A1(n4360), .A2(n4361), .A3(n4362), .ZN(n3938) );
  AOI211_X1 U3691 ( .C1(n4017), .C2(n4363), .A(n4364), .B(n4365), .ZN(n4362)
         );
  MUX2_X1 U3692 ( .A(n4366), .B(n4367), .S(\unit_decode/IMMreg/ffi_16/n4 ), 
        .Z(n4365) );
  NOR2_X1 U3693 ( .A1(n4368), .A2(n4024), .ZN(n4367) );
  MUX2_X1 U3694 ( .A(n4126), .B(n4036), .S(n4369), .Z(n4366) );
  OAI222_X1 U3695 ( .A1(n4352), .A2(n4254), .B1(n4333), .B2(n4253), .C1(n4370), 
        .C2(n4239), .ZN(n4364) );
  INV_X1 U3696 ( .A(n4321), .ZN(n4333) );
  INV_X1 U3697 ( .A(n4371), .ZN(n4361) );
  OAI222_X1 U3698 ( .A1(n4101), .A2(n4269), .B1(n4026), .B2(n4238), .C1(n4076), 
        .C2(n4193), .ZN(n4371) );
  OAI21_X1 U3699 ( .B1(n4372), .B2(n4373), .A(n4374), .ZN(n4076) );
  INV_X1 U3700 ( .A(n4258), .ZN(n4238) );
  OAI221_X1 U3701 ( .B1(n4369), .B2(n4166), .C1(n4237), .C2(n4272), .A(n4375), 
        .ZN(n4258) );
  AOI21_X1 U3702 ( .B1(n4376), .B2(n4377), .A(n4378), .ZN(n4375) );
  AOI222_X1 U3703 ( .A1(n4028), .A2(n4298), .B1(n4118), .B2(n4262), .C1(n4120), 
        .C2(n4279), .ZN(n4360) );
  NOR2_X1 U3704 ( .A1(RST), .A2(n3992), .ZN(n4921) );
  AND3_X1 U3705 ( .A1(n4379), .A2(n4380), .A3(n4381), .ZN(n3992) );
  AOI211_X1 U3706 ( .C1(n4028), .C2(n4321), .A(n4382), .B(n4383), .ZN(n4381)
         );
  MUX2_X1 U3707 ( .A(n4384), .B(n4385), .S(\unit_decode/IMMreg/ffi_17/n4 ), 
        .Z(n4383) );
  NOR2_X1 U3708 ( .A1(n4386), .A2(n4024), .ZN(n4385) );
  MUX2_X1 U3709 ( .A(n4126), .B(n4036), .S(n4387), .Z(n4384) );
  OAI222_X1 U3710 ( .A1(n4370), .A2(n4254), .B1(n4352), .B2(n4253), .C1(n4269), 
        .C2(n4026), .ZN(n4382) );
  INV_X1 U3711 ( .A(n4257), .ZN(n4269) );
  OAI221_X1 U3712 ( .B1(n4387), .B2(n4166), .C1(n4252), .C2(n4272), .A(n4388), 
        .ZN(n4257) );
  AOI21_X1 U3713 ( .B1(n4376), .B2(n4389), .A(n4378), .ZN(n4388) );
  INV_X1 U3714 ( .A(n4325), .ZN(n4352) );
  AOI222_X1 U3715 ( .A1(n4118), .A2(n4279), .B1(n4120), .B2(n4298), .C1(n4079), 
        .C2(n4106), .ZN(n4380) );
  AND2_X1 U3716 ( .A1(n4390), .A2(n4391), .ZN(n4079) );
  MUX2_X1 U3717 ( .A(n4374), .B(n4392), .S(n4393), .Z(n4390) );
  NAND2_X1 U3718 ( .A1(n4374), .A2(n4394), .ZN(n4392) );
  AOI222_X1 U3719 ( .A1(n4177), .A2(n4262), .B1(n4017), .B2(n4395), .C1(n4030), 
        .C2(n4363), .ZN(n4379) );
  NOR2_X1 U3720 ( .A1(RST), .A2(n3941), .ZN(n4922) );
  AND3_X1 U3721 ( .A1(n4396), .A2(n4397), .A3(n4398), .ZN(n3941) );
  AOI211_X1 U3722 ( .C1(n4028), .C2(n4325), .A(n4399), .B(n4400), .ZN(n4398)
         );
  MUX2_X1 U3723 ( .A(n4401), .B(n4402), .S(\unit_decode/IMMreg/ffi_18/n4 ), 
        .Z(n4400) );
  NOR2_X1 U3724 ( .A1(n4403), .A2(n4024), .ZN(n4402) );
  MUX2_X1 U3725 ( .A(n4126), .B(n4036), .S(n4404), .Z(n4401) );
  OAI222_X1 U3726 ( .A1(n4405), .A2(n4254), .B1(n4370), .B2(n4253), .C1(n4286), 
        .C2(n4026), .ZN(n4399) );
  INV_X1 U3727 ( .A(n4262), .ZN(n4286) );
  OAI221_X1 U3728 ( .B1(n4268), .B2(n4272), .C1(n4404), .C2(n4166), .A(n4406), 
        .ZN(n4262) );
  AOI21_X1 U3729 ( .B1(n4376), .B2(n4122), .A(n4378), .ZN(n4406) );
  AOI221_X1 U3730 ( .B1(n4118), .B2(n4298), .C1(n4120), .C2(n4321), .A(n4407), 
        .ZN(n4397) );
  AOI21_X1 U3731 ( .B1(n4077), .B2(n4072), .A(n4193), .ZN(n4407) );
  INV_X1 U3732 ( .A(n4408), .ZN(n4072) );
  AOI211_X1 U3733 ( .C1(n4409), .C2(n4373), .A(n4410), .B(n4411), .ZN(n4408)
         );
  OAI211_X1 U3734 ( .C1(n4373), .C2(n4411), .A(n4409), .B(n4410), .ZN(n4077)
         );
  AOI222_X1 U3735 ( .A1(n4177), .A2(n4279), .B1(n4017), .B2(n4412), .C1(n4030), 
        .C2(n4395), .ZN(n4396) );
  NOR2_X1 U3736 ( .A1(RST), .A2(n3944), .ZN(n4923) );
  AND3_X1 U3737 ( .A1(n4413), .A2(n4414), .A3(n4415), .ZN(n3944) );
  AOI211_X1 U3738 ( .C1(n4017), .C2(n4416), .A(n4417), .B(n4418), .ZN(n4415)
         );
  MUX2_X1 U3739 ( .A(n4419), .B(n4420), .S(\unit_decode/IMMreg/ffi_19/n4 ), 
        .Z(n4418) );
  NOR2_X1 U3740 ( .A1(n4421), .A2(n4024), .ZN(n4420) );
  MUX2_X1 U3741 ( .A(n4126), .B(n4036), .S(n4422), .Z(n4419) );
  OAI222_X1 U3742 ( .A1(n4423), .A2(n4254), .B1(n4405), .B2(n4253), .C1(n4424), 
        .C2(n4239), .ZN(n4417) );
  AOI222_X1 U3743 ( .A1(n4177), .A2(n4298), .B1(n4106), .B2(n4053), .C1(n4121), 
        .C2(n4279), .ZN(n4414) );
  OAI221_X1 U3744 ( .B1(n4285), .B2(n4272), .C1(n4422), .C2(n4166), .A(n4425), 
        .ZN(n4279) );
  AOI21_X1 U3745 ( .B1(n4376), .B2(n4426), .A(n4378), .ZN(n4425) );
  XNOR2_X1 U3746 ( .A(n4427), .B(n4428), .ZN(n4053) );
  OAI21_X1 U3747 ( .B1(n4429), .B2(n4373), .A(n4430), .ZN(n4427) );
  OAI21_X1 U3748 ( .B1(n4431), .B2(n4410), .A(n4432), .ZN(n4430) );
  INV_X1 U3749 ( .A(n4409), .ZN(n4431) );
  OAI21_X1 U3750 ( .B1(n4433), .B2(n4393), .A(n4434), .ZN(n4409) );
  AND2_X1 U3751 ( .A1(n4435), .A2(n4369), .ZN(n4433) );
  AOI222_X1 U3752 ( .A1(n4028), .A2(n4345), .B1(n4118), .B2(n4321), .C1(n4120), 
        .C2(n4325), .ZN(n4413) );
  NOR2_X1 U3753 ( .A1(RST), .A2(n3949), .ZN(n4924) );
  AND3_X1 U3754 ( .A1(n4436), .A2(n4437), .A3(n4438), .ZN(n3949) );
  AOI211_X1 U3755 ( .C1(n4017), .C2(n4439), .A(n4440), .B(n4441), .ZN(n4438)
         );
  MUX2_X1 U3756 ( .A(n4442), .B(n4443), .S(\unit_decode/IMMreg/ffi_20/n4 ), 
        .Z(n4441) );
  NOR2_X1 U3757 ( .A1(n4444), .A2(n4024), .ZN(n4443) );
  MUX2_X1 U3758 ( .A(n4126), .B(n4036), .S(n4445), .Z(n4442) );
  OAI222_X1 U3759 ( .A1(n4424), .A2(n4254), .B1(n4423), .B2(n4253), .C1(n4446), 
        .C2(n4239), .ZN(n4440) );
  AOI222_X1 U3760 ( .A1(n4177), .A2(n4321), .B1(n4121), .B2(n4298), .C1(n4070), 
        .C2(n4106), .ZN(n4437) );
  INV_X1 U3761 ( .A(n4447), .ZN(n4070) );
  OAI21_X1 U3762 ( .B1(n4448), .B2(n4449), .A(n4450), .ZN(n4447) );
  OAI221_X1 U3763 ( .B1(n4304), .B2(n4272), .C1(n4445), .C2(n4166), .A(n4451), 
        .ZN(n4298) );
  AOI21_X1 U3764 ( .B1(n4376), .B2(n4167), .A(n4378), .ZN(n4451) );
  AOI222_X1 U3765 ( .A1(n4028), .A2(n4363), .B1(n4118), .B2(n4325), .C1(n4120), 
        .C2(n4345), .ZN(n4436) );
  NOR2_X1 U3766 ( .A1(RST), .A2(n3996), .ZN(n4925) );
  AND3_X1 U3767 ( .A1(n4452), .A2(n4453), .A3(n4454), .ZN(n3996) );
  AOI211_X1 U3768 ( .C1(n4017), .C2(n4455), .A(n4456), .B(n4457), .ZN(n4454)
         );
  MUX2_X1 U3769 ( .A(n4458), .B(n4459), .S(\unit_decode/IMMreg/ffi_21/n4 ), 
        .Z(n4457) );
  NOR2_X1 U3770 ( .A1(n4460), .A2(n4024), .ZN(n4459) );
  MUX2_X1 U3771 ( .A(n4126), .B(n4036), .S(n4461), .Z(n4458) );
  OAI222_X1 U3772 ( .A1(n4446), .A2(n4254), .B1(n4424), .B2(n4253), .C1(n4462), 
        .C2(n4239), .ZN(n4456) );
  INV_X1 U3773 ( .A(n4412), .ZN(n4424) );
  AOI222_X1 U3774 ( .A1(n4177), .A2(n4325), .B1(n4121), .B2(n4321), .C1(n4078), 
        .C2(n4106), .ZN(n4453) );
  NOR2_X1 U3775 ( .A1(n4463), .A2(n4464), .ZN(n4078) );
  MUX2_X1 U3776 ( .A(n4465), .B(n4466), .S(n4450), .Z(n4463) );
  AND2_X1 U3777 ( .A1(n4467), .A2(n4468), .ZN(n4466) );
  OAI221_X1 U3778 ( .B1(n4316), .B2(n4272), .C1(n4461), .C2(n4166), .A(n4469), 
        .ZN(n4321) );
  AOI21_X1 U3779 ( .B1(n4376), .B2(n4470), .A(n4378), .ZN(n4469) );
  AOI222_X1 U3780 ( .A1(n4028), .A2(n4395), .B1(n4118), .B2(n4345), .C1(n4120), 
        .C2(n4363), .ZN(n4452) );
  NOR2_X1 U3781 ( .A1(RST), .A2(n3951), .ZN(n4926) );
  AND3_X1 U3782 ( .A1(n4471), .A2(n4472), .A3(n4473), .ZN(n3951) );
  AOI211_X1 U3783 ( .C1(n4017), .C2(n4474), .A(n4475), .B(n4476), .ZN(n4473)
         );
  MUX2_X1 U3784 ( .A(n4477), .B(n4478), .S(\unit_decode/IMMreg/ffi_22/n4 ), 
        .Z(n4476) );
  NOR2_X1 U3785 ( .A1(n4479), .A2(n4024), .ZN(n4478) );
  MUX2_X1 U3786 ( .A(n4126), .B(n4036), .S(n4480), .Z(n4477) );
  OAI222_X1 U3787 ( .A1(n4462), .A2(n4254), .B1(n4446), .B2(n4253), .C1(n4481), 
        .C2(n4239), .ZN(n4475) );
  AOI222_X1 U3788 ( .A1(n4177), .A2(n4345), .B1(n4069), .B2(n4106), .C1(n4121), 
        .C2(n4325), .ZN(n4472) );
  OAI221_X1 U3789 ( .B1(n4331), .B2(n4272), .C1(n4480), .C2(n4166), .A(n4482), 
        .ZN(n4325) );
  AOI21_X1 U3790 ( .B1(n4376), .B2(n4483), .A(n4378), .ZN(n4482) );
  INV_X1 U3791 ( .A(n4484), .ZN(n4069) );
  OAI21_X1 U3792 ( .B1(n4485), .B2(n4486), .A(n4487), .ZN(n4484) );
  AOI222_X1 U3793 ( .A1(n4028), .A2(n4412), .B1(n4118), .B2(n4363), .C1(n4120), 
        .C2(n4395), .ZN(n4471) );
  NOR2_X1 U3794 ( .A1(RST), .A2(n4000), .ZN(n4927) );
  AND3_X1 U3795 ( .A1(n4488), .A2(n4489), .A3(n4490), .ZN(n4000) );
  AOI211_X1 U3796 ( .C1(n4028), .C2(n4416), .A(n4491), .B(n4492), .ZN(n4490)
         );
  MUX2_X1 U3797 ( .A(n4493), .B(n4494), .S(\unit_decode/IMMreg/ffi_23/n4 ), 
        .Z(n4492) );
  NOR2_X1 U3798 ( .A1(n4495), .A2(n4024), .ZN(n4494) );
  MUX2_X1 U3799 ( .A(n4126), .B(n4036), .S(n4496), .Z(n4493) );
  OAI222_X1 U3800 ( .A1(n4481), .A2(n4254), .B1(n4462), .B2(n4253), .C1(n4370), 
        .C2(n4026), .ZN(n4491) );
  INV_X1 U3801 ( .A(n4345), .ZN(n4370) );
  OAI221_X1 U3802 ( .B1(n4351), .B2(n4272), .C1(n4496), .C2(n4166), .A(n4497), 
        .ZN(n4345) );
  AOI21_X1 U3803 ( .B1(n4376), .B2(n4220), .A(n4378), .ZN(n4497) );
  INV_X1 U3804 ( .A(n4439), .ZN(n4462) );
  AOI222_X1 U3805 ( .A1(n4118), .A2(n4395), .B1(n4120), .B2(n4412), .C1(n4063), 
        .C2(n4106), .ZN(n4489) );
  XNOR2_X1 U3806 ( .A(n4498), .B(n4499), .ZN(n4063) );
  NOR2_X1 U3807 ( .A1(n4500), .A2(n4501), .ZN(n4499) );
  INV_X1 U3808 ( .A(n4487), .ZN(n4500) );
  NAND2_X1 U3809 ( .A1(n4485), .A2(n4486), .ZN(n4487) );
  NAND2_X1 U3810 ( .A1(n4502), .A2(n4503), .ZN(n4486) );
  NAND3_X1 U3811 ( .A1(n4504), .A2(n4449), .A3(n4465), .ZN(n4503) );
  AOI222_X1 U3812 ( .A1(n4177), .A2(n4363), .B1(n4017), .B2(n4505), .C1(n4030), 
        .C2(n4474), .ZN(n4488) );
  NOR2_X1 U3813 ( .A1(RST), .A2(n3954), .ZN(n4928) );
  AND3_X1 U3814 ( .A1(n4506), .A2(n4507), .A3(n4508), .ZN(n3954) );
  AOI211_X1 U3815 ( .C1(n4028), .C2(n4439), .A(n4509), .B(n4510), .ZN(n4508)
         );
  MUX2_X1 U3816 ( .A(n4511), .B(n4512), .S(\unit_decode/IMMreg/ffi_24/n4 ), 
        .Z(n4510) );
  NOR2_X1 U3817 ( .A1(n4513), .A2(n4024), .ZN(n4512) );
  MUX2_X1 U3818 ( .A(n4126), .B(n4036), .S(n4514), .Z(n4511) );
  OAI222_X1 U3819 ( .A1(n4515), .A2(n4254), .B1(n4481), .B2(n4253), .C1(n4405), 
        .C2(n4026), .ZN(n4509) );
  INV_X1 U3820 ( .A(n4363), .ZN(n4405) );
  OAI211_X1 U3821 ( .C1(n4369), .C2(n4272), .A(n4516), .B(n4517), .ZN(n4363)
         );
  AOI222_X1 U3822 ( .A1(n4518), .A2(n4377), .B1(n4519), .B2(n4513), .C1(n4376), 
        .C2(n4236), .ZN(n4517) );
  AOI222_X1 U3823 ( .A1(n4118), .A2(n4412), .B1(n4120), .B2(n4416), .C1(n4083), 
        .C2(n4106), .ZN(n4507) );
  XOR2_X1 U3824 ( .A(n4520), .B(n4521), .Z(n4083) );
  NAND2_X1 U3825 ( .A1(n4522), .A2(n4523), .ZN(n4520) );
  INV_X1 U3826 ( .A(n4524), .ZN(n4522) );
  AOI222_X1 U3827 ( .A1(n4177), .A2(n4395), .B1(n4017), .B2(n4525), .C1(n4030), 
        .C2(n4505), .ZN(n4506) );
  NOR2_X1 U3828 ( .A1(RST), .A2(n4004), .ZN(n4929) );
  AND3_X1 U3829 ( .A1(n4526), .A2(n4527), .A3(n4528), .ZN(n4004) );
  AOI211_X1 U3830 ( .C1(n4028), .C2(n4455), .A(n4529), .B(n4530), .ZN(n4528)
         );
  MUX2_X1 U3831 ( .A(n4531), .B(n4532), .S(\unit_decode/IMMreg/ffi_25/n4 ), 
        .Z(n4530) );
  NOR2_X1 U3832 ( .A1(n4533), .A2(n4024), .ZN(n4532) );
  MUX2_X1 U3833 ( .A(n4126), .B(n4036), .S(n4534), .Z(n4531) );
  OAI222_X1 U3834 ( .A1(n4535), .A2(n4254), .B1(n4515), .B2(n4253), .C1(n4423), 
        .C2(n4026), .ZN(n4529) );
  INV_X1 U3835 ( .A(n4395), .ZN(n4423) );
  OAI211_X1 U3836 ( .C1(n4387), .C2(n4272), .A(n4516), .B(n4536), .ZN(n4395)
         );
  AOI222_X1 U3837 ( .A1(n4518), .A2(n4389), .B1(n4519), .B2(n4533), .C1(n4376), 
        .C2(n4251), .ZN(n4536) );
  INV_X1 U3838 ( .A(n4474), .ZN(n4515) );
  AOI222_X1 U3839 ( .A1(n4118), .A2(n4416), .B1(n4120), .B2(n4439), .C1(n4064), 
        .C2(n4106), .ZN(n4527) );
  XOR2_X1 U3840 ( .A(n4537), .B(n4538), .Z(n4064) );
  AOI222_X1 U3841 ( .A1(n4177), .A2(n4412), .B1(n4017), .B2(n4539), .C1(n4030), 
        .C2(n4525), .ZN(n4526) );
  NOR2_X1 U3842 ( .A1(RST), .A2(n3957), .ZN(n4930) );
  AND3_X1 U3843 ( .A1(n4540), .A2(n4541), .A3(n4542), .ZN(n3957) );
  AOI211_X1 U3844 ( .C1(n4017), .C2(n4543), .A(n4544), .B(n4545), .ZN(n4542)
         );
  MUX2_X1 U3845 ( .A(n4546), .B(n4547), .S(\unit_decode/IMMreg/ffi_26/n4 ), 
        .Z(n4545) );
  NOR2_X1 U3846 ( .A1(n4548), .A2(n4024), .ZN(n4547) );
  MUX2_X1 U3847 ( .A(n4126), .B(n4036), .S(n4549), .Z(n4546) );
  OAI222_X1 U3848 ( .A1(n4550), .A2(n4254), .B1(n4535), .B2(n4253), .C1(n4551), 
        .C2(n4239), .ZN(n4544) );
  INV_X1 U3849 ( .A(n4505), .ZN(n4535) );
  AOI222_X1 U3850 ( .A1(n4177), .A2(n4416), .B1(n4084), .B2(n4106), .C1(n4121), 
        .C2(n4412), .ZN(n4541) );
  OAI211_X1 U3851 ( .C1(n4404), .C2(n4272), .A(n4516), .B(n4552), .ZN(n4412)
         );
  AOI222_X1 U3852 ( .A1(n4518), .A2(n4122), .B1(n4519), .B2(n4548), .C1(n4376), 
        .C2(n4267), .ZN(n4552) );
  INV_X1 U3853 ( .A(n4268), .ZN(n4267) );
  INV_X1 U3854 ( .A(n4549), .ZN(n4548) );
  XOR2_X1 U3855 ( .A(n4553), .B(n4554), .Z(n4084) );
  AOI222_X1 U3856 ( .A1(n4028), .A2(n4474), .B1(n4118), .B2(n4439), .C1(n4120), 
        .C2(n4455), .ZN(n4540) );
  NOR2_X1 U3857 ( .A1(RST), .A2(n4007), .ZN(n4931) );
  AND3_X1 U3858 ( .A1(n4555), .A2(n4556), .A3(n4557), .ZN(n4007) );
  AOI211_X1 U3859 ( .C1(n4028), .C2(n4505), .A(n4558), .B(n4559), .ZN(n4557)
         );
  MUX2_X1 U3860 ( .A(n4560), .B(n4561), .S(\unit_decode/IMMreg/ffi_27/n4 ), 
        .Z(n4559) );
  NOR2_X1 U3861 ( .A1(n4562), .A2(n4024), .ZN(n4561) );
  MUX2_X1 U3862 ( .A(n4126), .B(n4036), .S(n4563), .Z(n4560) );
  OAI222_X1 U3863 ( .A1(n4551), .A2(n4254), .B1(n4550), .B2(n4253), .C1(n4446), 
        .C2(n4026), .ZN(n4558) );
  INV_X1 U3864 ( .A(n4416), .ZN(n4446) );
  OAI211_X1 U3865 ( .C1(n4422), .C2(n4272), .A(n4516), .B(n4564), .ZN(n4416)
         );
  AOI222_X1 U3866 ( .A1(n4518), .A2(n4426), .B1(n4519), .B2(n4562), .C1(n4376), 
        .C2(n4284), .ZN(n4564) );
  INV_X1 U3867 ( .A(n4285), .ZN(n4284) );
  INV_X1 U3868 ( .A(n4525), .ZN(n4550) );
  AOI222_X1 U3869 ( .A1(n4118), .A2(n4455), .B1(n4120), .B2(n4474), .C1(n4065), 
        .C2(n4106), .ZN(n4556) );
  XOR2_X1 U3870 ( .A(n4563), .B(n4565), .Z(n4065) );
  XNOR2_X1 U3871 ( .A(n4566), .B(n4567), .ZN(n4565) );
  AOI222_X1 U3872 ( .A1(n4177), .A2(n4439), .B1(n4017), .B2(n4568), .C1(n4030), 
        .C2(n4543), .ZN(n4555) );
  NOR2_X1 U3873 ( .A1(RST), .A2(n3960), .ZN(n4932) );
  AND3_X1 U3874 ( .A1(n4569), .A2(n4570), .A3(n4571), .ZN(n3960) );
  AOI211_X1 U3875 ( .C1(n4017), .C2(n4572), .A(n4573), .B(n4574), .ZN(n4571)
         );
  MUX2_X1 U3876 ( .A(n4575), .B(n4576), .S(\unit_decode/IMMreg/ffi_28/n4 ), 
        .Z(n4574) );
  NOR2_X1 U3877 ( .A1(n4577), .A2(n4024), .ZN(n4576) );
  MUX2_X1 U3878 ( .A(n4126), .B(n4036), .S(n4578), .Z(n4575) );
  OAI222_X1 U3879 ( .A1(n4579), .A2(n4254), .B1(n4551), .B2(n4253), .C1(n4580), 
        .C2(n4239), .ZN(n4573) );
  INV_X1 U3880 ( .A(n4030), .ZN(n4239) );
  INV_X1 U3881 ( .A(n4539), .ZN(n4551) );
  AOI222_X1 U3882 ( .A1(n4177), .A2(n4455), .B1(n4106), .B2(n4054), .C1(n4121), 
        .C2(n4439), .ZN(n4570) );
  OAI211_X1 U3883 ( .C1(n4445), .C2(n4272), .A(n4516), .B(n4581), .ZN(n4439)
         );
  AOI222_X1 U3884 ( .A1(n4518), .A2(n4167), .B1(n4519), .B2(n4577), .C1(n4376), 
        .C2(n4303), .ZN(n4581) );
  XNOR2_X1 U3885 ( .A(n4582), .B(n4095), .ZN(n4054) );
  AOI222_X1 U3886 ( .A1(n4028), .A2(n4525), .B1(n4118), .B2(n4474), .C1(n4120), 
        .C2(n4505), .ZN(n4569) );
  NOR2_X1 U3887 ( .A1(RST), .A2(n3965), .ZN(n4933) );
  AND3_X1 U3888 ( .A1(n4583), .A2(n4584), .A3(n4585), .ZN(n3965) );
  AOI211_X1 U3889 ( .C1(n4028), .C2(n4539), .A(n4586), .B(n4587), .ZN(n4585)
         );
  MUX2_X1 U3890 ( .A(n4588), .B(n4589), .S(\unit_decode/IMMreg/ffi_29/n4 ), 
        .Z(n4587) );
  NOR2_X1 U3891 ( .A1(n4590), .A2(n4024), .ZN(n4589) );
  MUX2_X1 U3892 ( .A(n4126), .B(n4036), .S(n4591), .Z(n4588) );
  OAI222_X1 U3893 ( .A1(n4580), .A2(n4254), .B1(n4579), .B2(n4253), .C1(n4481), 
        .C2(n4026), .ZN(n4586) );
  INV_X1 U3894 ( .A(n4455), .ZN(n4481) );
  OAI211_X1 U3895 ( .C1(n4461), .C2(n4272), .A(n4516), .B(n4592), .ZN(n4455)
         );
  AOI222_X1 U3896 ( .A1(n4518), .A2(n4470), .B1(n4519), .B2(n4590), .C1(n4376), 
        .C2(n4315), .ZN(n4592) );
  INV_X1 U3897 ( .A(n4032), .ZN(n4253) );
  INV_X1 U3898 ( .A(n4543), .ZN(n4579) );
  INV_X1 U3899 ( .A(n4108), .ZN(n4254) );
  INV_X1 U3900 ( .A(n4568), .ZN(n4580) );
  AOI222_X1 U3901 ( .A1(n4118), .A2(n4505), .B1(n4120), .B2(n4525), .C1(n4081), 
        .C2(n4106), .ZN(n4584) );
  XNOR2_X1 U3902 ( .A(n4093), .B(n4593), .ZN(n4081) );
  OAI21_X1 U3903 ( .B1(n4096), .B2(n4095), .A(n4594), .ZN(n4593) );
  OAI21_X1 U3904 ( .B1(n4595), .B2(n4577), .A(n4594), .ZN(n4095) );
  AOI222_X1 U3905 ( .A1(n4177), .A2(n4474), .B1(n4017), .B2(n4596), .C1(n4030), 
        .C2(n4572), .ZN(n4583) );
  NOR2_X1 U3906 ( .A1(RST), .A2(n4009), .ZN(n4934) );
  AND3_X1 U3907 ( .A1(n4597), .A2(n4598), .A3(n4599), .ZN(n4009) );
  AOI211_X1 U3908 ( .C1(n4028), .C2(n4543), .A(n4600), .B(n4601), .ZN(n4599)
         );
  MUX2_X1 U3909 ( .A(n4602), .B(n4603), .S(\unit_decode/IMMreg/ffi_30/n4 ), 
        .Z(n4601) );
  NOR2_X1 U3910 ( .A1(n4604), .A2(n4024), .ZN(n4603) );
  MUX2_X1 U3911 ( .A(n4126), .B(n4036), .S(n4605), .Z(n4602) );
  INV_X1 U3912 ( .A(n4606), .ZN(n4600) );
  AOI222_X1 U3913 ( .A1(n4572), .A2(n4108), .B1(n4568), .B2(n4032), .C1(n4474), 
        .C2(n4121), .ZN(n4606) );
  OAI211_X1 U3914 ( .C1(n4480), .C2(n4272), .A(n4516), .B(n4607), .ZN(n4474)
         );
  AOI222_X1 U3915 ( .A1(n4518), .A2(n4483), .B1(n4519), .B2(n4604), .C1(n4376), 
        .C2(n4330), .ZN(n4607) );
  AOI222_X1 U3916 ( .A1(n4118), .A2(n4525), .B1(n4120), .B2(n4539), .C1(n4066), 
        .C2(n4106), .ZN(n4598) );
  XOR2_X1 U3917 ( .A(n4094), .B(n4608), .Z(n4066) );
  AOI21_X1 U3918 ( .B1(n4582), .B2(n4609), .A(n4610), .ZN(n4608) );
  AOI222_X1 U3919 ( .A1(n4177), .A2(n4505), .B1(n4017), .B2(n4611), .C1(n4030), 
        .C2(n4596), .ZN(n4597) );
  NOR2_X1 U3920 ( .A1(RST), .A2(n3968), .ZN(n4935) );
  AND3_X1 U3921 ( .A1(n4612), .A2(n4613), .A3(n4614), .ZN(n3968) );
  AOI211_X1 U3922 ( .C1(n4032), .C2(n4572), .A(n4615), .B(n4616), .ZN(n4614)
         );
  MUX2_X1 U3923 ( .A(n4617), .B(n4618), .S(\unit_decode/IMMreg/ffi_31/n4 ), 
        .Z(n4616) );
  NOR2_X1 U3924 ( .A1(n4619), .A2(n4024), .ZN(n4618) );
  MUX2_X1 U3925 ( .A(n4126), .B(n4036), .S(n4097), .Z(n4617) );
  INV_X1 U3926 ( .A(n4620), .ZN(n4615) );
  AOI222_X1 U3927 ( .A1(n4596), .A2(n4108), .B1(n4611), .B2(n4030), .C1(n4568), 
        .C2(n4028), .ZN(n4620) );
  OAI221_X1 U3928 ( .B1(n4285), .B2(n4621), .C1(n4563), .C2(n4272), .A(n4622), 
        .ZN(n4568) );
  AOI221_X1 U3929 ( .B1(n4623), .B2(n4426), .C1(n4376), .C2(n4421), .A(n4624), 
        .ZN(n4622) );
  OAI221_X1 U3930 ( .B1(n4331), .B2(n4621), .C1(n4605), .C2(n4272), .A(n4625), 
        .ZN(n4611) );
  AOI221_X1 U3931 ( .B1(n4623), .B2(n4483), .C1(n4376), .C2(n4479), .A(n4624), 
        .ZN(n4625) );
  INV_X1 U3932 ( .A(n4480), .ZN(n4479) );
  OAI221_X1 U3933 ( .B1(n4316), .B2(n4621), .C1(n4591), .C2(n4272), .A(n4626), 
        .ZN(n4596) );
  AOI221_X1 U3934 ( .B1(n4623), .B2(n4470), .C1(n4376), .C2(n4460), .A(n4624), 
        .ZN(n4626) );
  INV_X1 U3935 ( .A(n4183), .ZN(n4470) );
  OAI221_X1 U3936 ( .B1(n4304), .B2(n4621), .C1(n4578), .C2(n4272), .A(n4627), 
        .ZN(n4572) );
  AOI221_X1 U3937 ( .B1(n4623), .B2(n4167), .C1(n4376), .C2(n4444), .A(n4624), 
        .ZN(n4627) );
  INV_X1 U3938 ( .A(n4168), .ZN(n4167) );
  NOR4_X1 U3939 ( .A1(n4629), .A2(n3786), .A3(n4201), .A4(n4630), .ZN(n4628)
         );
  AOI221_X1 U3940 ( .B1(n4518), .B2(n4350), .C1(n4631), .C2(n4619), .A(n4632), 
        .ZN(n4629) );
  OAI22_X1 U3941 ( .A1(n4221), .A2(n4633), .B1(n4496), .B2(n4634), .ZN(n4632)
         );
  INV_X1 U3942 ( .A(n4272), .ZN(n4631) );
  XNOR2_X1 U3943 ( .A(n4635), .B(n4099), .ZN(n4051) );
  XNOR2_X1 U3944 ( .A(n4097), .B(n4098), .ZN(n4099) );
  XNOR2_X1 U3945 ( .A(\unit_decode/IMMreg/ffi_31/n4 ), .B(n3785), .ZN(n4098)
         );
  OAI21_X1 U3946 ( .B1(n4582), .B2(n4092), .A(n4636), .ZN(n4635) );
  OAI21_X1 U3947 ( .B1(n4637), .B2(n4094), .A(n4638), .ZN(n4636) );
  INV_X1 U3948 ( .A(n4609), .ZN(n4637) );
  OAI21_X1 U3949 ( .B1(n4639), .B2(n4093), .A(n4640), .ZN(n4609) );
  NOR2_X1 U3950 ( .A1(n4595), .A2(n4577), .ZN(n4639) );
  OAI21_X1 U3951 ( .B1(n4641), .B2(n4094), .A(n4638), .ZN(n4092) );
  OAI21_X1 U3952 ( .B1(n4604), .B2(n4642), .A(n4638), .ZN(n4094) );
  NAND2_X1 U3953 ( .A1(n4604), .A2(n4642), .ZN(n4638) );
  XOR2_X1 U3954 ( .A(\unit_decode/IMMreg/ffi_30/n4 ), .B(n4862), .Z(n4642) );
  INV_X1 U3955 ( .A(n4605), .ZN(n4604) );
  MUX2_X1 U3956 ( .A(\unit_decode/Areg/ffi_30/n4 ), .B(
        \unit_decode/NPC1reg/ffi_30/n4 ), .S(n4012), .Z(n4605) );
  INV_X1 U3957 ( .A(n4610), .ZN(n4641) );
  OAI21_X1 U3958 ( .B1(n4093), .B2(n4594), .A(n4640), .ZN(n4610) );
  NAND2_X1 U3959 ( .A1(n4595), .A2(n4577), .ZN(n4594) );
  INV_X1 U3960 ( .A(n4578), .ZN(n4577) );
  MUX2_X1 U3961 ( .A(\unit_decode/Areg/ffi_28/n4 ), .B(
        \unit_decode/NPC1reg/ffi_28/n4 ), .S(n4012), .Z(n4578) );
  XOR2_X1 U3962 ( .A(\unit_decode/IMMreg/ffi_28/n4 ), .B(n4862), .Z(n4595) );
  OAI21_X1 U3963 ( .B1(n4643), .B2(n4590), .A(n4640), .ZN(n4093) );
  NAND2_X1 U3964 ( .A1(n4643), .A2(n4590), .ZN(n4640) );
  INV_X1 U3965 ( .A(n4591), .ZN(n4590) );
  MUX2_X1 U3966 ( .A(\unit_decode/Areg/ffi_29/n4 ), .B(
        \unit_decode/NPC1reg/ffi_29/n4 ), .S(n4012), .Z(n4591) );
  XOR2_X1 U3967 ( .A(\unit_decode/IMMreg/ffi_29/n4 ), .B(n4862), .Z(n4643) );
  INV_X1 U3968 ( .A(n4096), .ZN(n4582) );
  OAI22_X1 U3969 ( .A1(n4567), .A2(n4566), .B1(n4644), .B2(n4562), .ZN(n4096)
         );
  INV_X1 U3970 ( .A(n4563), .ZN(n4562) );
  MUX2_X1 U3971 ( .A(\unit_decode/Areg/ffi_27/n4 ), .B(
        \unit_decode/NPC1reg/ffi_27/n4 ), .S(n4012), .Z(n4563) );
  AND2_X1 U3972 ( .A1(n4566), .A2(n4567), .ZN(n4644) );
  OAI22_X1 U3973 ( .A1(n4549), .A2(n4645), .B1(n4554), .B2(n4553), .ZN(n4566)
         );
  XNOR2_X1 U3974 ( .A(n4549), .B(n4645), .ZN(n4553) );
  AOI21_X1 U3975 ( .B1(n4537), .B2(n4538), .A(n4646), .ZN(n4554) );
  INV_X1 U3976 ( .A(n4647), .ZN(n4646) );
  INV_X1 U3977 ( .A(n4648), .ZN(n4538) );
  OAI21_X1 U3978 ( .B1(n4649), .B2(n4533), .A(n4647), .ZN(n4648) );
  NAND2_X1 U3979 ( .A1(n4649), .A2(n4533), .ZN(n4647) );
  INV_X1 U3980 ( .A(n4534), .ZN(n4533) );
  XOR2_X1 U3981 ( .A(\unit_decode/IMMreg/ffi_25/n4 ), .B(n4862), .Z(n4649) );
  OAI21_X1 U3982 ( .B1(n4524), .B2(n4521), .A(n4523), .ZN(n4537) );
  NAND2_X1 U3983 ( .A1(n4513), .A2(n4650), .ZN(n4523) );
  AOI22_X1 U3984 ( .A1(n4495), .A2(n4651), .B1(n4652), .B2(n4498), .ZN(n4521)
         );
  XNOR2_X1 U3985 ( .A(n4496), .B(n4651), .ZN(n4498) );
  INV_X1 U3986 ( .A(n4653), .ZN(n4652) );
  AOI21_X1 U3987 ( .B1(n4485), .B2(n4654), .A(n4501), .ZN(n4653) );
  OAI21_X1 U3988 ( .B1(n4467), .B2(n4450), .A(n4502), .ZN(n4654) );
  AOI21_X1 U3989 ( .B1(n4655), .B2(n4460), .A(n4464), .ZN(n4502) );
  NOR2_X1 U3990 ( .A1(n4468), .A2(n4467), .ZN(n4464) );
  NAND2_X1 U3991 ( .A1(n4448), .A2(n4449), .ZN(n4450) );
  OAI21_X1 U3992 ( .B1(n4422), .B2(n4656), .A(n4657), .ZN(n4449) );
  OAI21_X1 U3993 ( .B1(n4658), .B2(n4429), .A(n4428), .ZN(n4657) );
  XNOR2_X1 U3994 ( .A(n4421), .B(n4656), .ZN(n4428) );
  INV_X1 U3995 ( .A(n4422), .ZN(n4421) );
  OAI21_X1 U3996 ( .B1(n4659), .B2(n4410), .A(n4432), .ZN(n4429) );
  INV_X1 U3997 ( .A(n4411), .ZN(n4659) );
  NAND2_X1 U3998 ( .A1(n4434), .A2(n4391), .ZN(n4411) );
  OR2_X1 U3999 ( .A1(n4393), .A2(n4394), .ZN(n4391) );
  INV_X1 U4000 ( .A(n4660), .ZN(n4394) );
  NOR3_X1 U4001 ( .A1(n4374), .A2(n4393), .A3(n4410), .ZN(n4658) );
  OAI21_X1 U4002 ( .B1(n4661), .B2(n4403), .A(n4432), .ZN(n4410) );
  NAND2_X1 U4003 ( .A1(n4661), .A2(n4403), .ZN(n4432) );
  XOR2_X1 U4004 ( .A(\unit_decode/IMMreg/ffi_18/n4 ), .B(n4862), .Z(n4661) );
  OAI21_X1 U4005 ( .B1(n4662), .B2(n4386), .A(n4434), .ZN(n4393) );
  NAND2_X1 U4006 ( .A1(n4662), .A2(n4386), .ZN(n4434) );
  XOR2_X1 U4007 ( .A(\unit_decode/IMMreg/ffi_17/n4 ), .B(n4862), .Z(n4662) );
  NAND2_X1 U4008 ( .A1(n4372), .A2(n4373), .ZN(n4374) );
  OAI21_X1 U4009 ( .B1(n4351), .B2(n4663), .A(n4664), .ZN(n4373) );
  OAI21_X1 U4010 ( .B1(n4665), .B2(n4356), .A(n4353), .ZN(n4664) );
  XNOR2_X1 U4011 ( .A(n4350), .B(n4663), .ZN(n4353) );
  OAI22_X1 U4012 ( .A1(n4331), .A2(n4666), .B1(n4340), .B2(n4337), .ZN(n4356)
         );
  INV_X1 U4013 ( .A(n4338), .ZN(n4340) );
  OAI21_X1 U4014 ( .B1(n4318), .B2(n4320), .A(n4358), .ZN(n4338) );
  NAND2_X1 U4015 ( .A1(n4667), .A2(n4315), .ZN(n4358) );
  INV_X1 U4016 ( .A(n4316), .ZN(n4315) );
  NOR4_X1 U4017 ( .A1(n4319), .A2(n4318), .A3(n4306), .A4(n4337), .ZN(n4665)
         );
  XOR2_X1 U4018 ( .A(n4330), .B(n4666), .Z(n4337) );
  XNOR2_X1 U4019 ( .A(\unit_decode/IMMreg/ffi_14/n4 ), .B(n4862), .ZN(n4666)
         );
  INV_X1 U4020 ( .A(n4331), .ZN(n4330) );
  MUX2_X1 U4021 ( .A(\unit_decode/Areg/ffi_14/n4 ), .B(
        \unit_decode/NPC1reg/ffi_14/n4 ), .S(n4012), .Z(n4331) );
  OAI21_X1 U4022 ( .B1(n4359), .B2(n4303), .A(n4320), .ZN(n4306) );
  NAND2_X1 U4023 ( .A1(n4359), .A2(n4303), .ZN(n4320) );
  INV_X1 U4024 ( .A(n4304), .ZN(n4303) );
  MUX2_X1 U4025 ( .A(\unit_decode/Areg/ffi_12/n4 ), .B(
        \unit_decode/NPC1reg/ffi_12/n4 ), .S(n4012), .Z(n4304) );
  XOR2_X1 U4026 ( .A(\unit_decode/IMMreg/ffi_12/n4 ), .B(n4862), .Z(n4359) );
  XOR2_X1 U4027 ( .A(n4316), .B(n4667), .Z(n4318) );
  XOR2_X1 U4028 ( .A(\unit_decode/IMMreg/ffi_13/n4 ), .B(n4862), .Z(n4667) );
  MUX2_X1 U4029 ( .A(\unit_decode/Areg/ffi_13/n4 ), .B(
        \unit_decode/NPC1reg/ffi_13/n4 ), .S(n4012), .Z(n4316) );
  INV_X1 U4030 ( .A(n4307), .ZN(n4319) );
  OAI22_X1 U4031 ( .A1(n4285), .A2(n4668), .B1(n4669), .B2(n4287), .ZN(n4307)
         );
  XNOR2_X1 U4032 ( .A(n4285), .B(n4668), .ZN(n4287) );
  AOI21_X1 U4033 ( .B1(n4275), .B2(n4670), .A(n4289), .ZN(n4669) );
  OAI21_X1 U4034 ( .B1(n4255), .B2(n4256), .A(n4292), .ZN(n4670) );
  OAI21_X1 U4035 ( .B1(n4671), .B2(n4251), .A(n4292), .ZN(n4256) );
  NAND2_X1 U4036 ( .A1(n4671), .A2(n4251), .ZN(n4292) );
  INV_X1 U4037 ( .A(n4252), .ZN(n4251) );
  XOR2_X1 U4038 ( .A(\unit_decode/IMMreg/ffi_9/n4 ), .B(n4862), .Z(n4671) );
  AND2_X1 U4039 ( .A1(n4243), .A2(n4290), .ZN(n4255) );
  NAND2_X1 U4040 ( .A1(n4241), .A2(n4242), .ZN(n4243) );
  OAI21_X1 U4041 ( .B1(n4225), .B2(n4226), .A(n4672), .ZN(n4242) );
  INV_X1 U4042 ( .A(n4673), .ZN(n4672) );
  AOI21_X1 U4043 ( .B1(n4226), .B2(n4225), .A(n4221), .ZN(n4673) );
  XOR2_X1 U4044 ( .A(\unit_decode/IMMreg/ffi_7/n4 ), .B(n3785), .Z(n4226) );
  AOI21_X1 U4045 ( .B1(n4483), .B2(n4674), .A(n4212), .ZN(n4225) );
  AOI21_X1 U4046 ( .B1(n4210), .B2(n4209), .A(n4211), .ZN(n4212) );
  XOR2_X1 U4047 ( .A(n4198), .B(n4674), .Z(n4211) );
  NAND2_X1 U4048 ( .A1(n4190), .A2(n4191), .ZN(n4209) );
  AOI21_X1 U4049 ( .B1(n4183), .B2(n4675), .A(n4676), .ZN(n4191) );
  AOI21_X1 U4050 ( .B1(n4677), .B2(n4171), .A(n4172), .ZN(n4190) );
  AND2_X1 U4051 ( .A1(n4174), .A2(n4168), .ZN(n4172) );
  AOI21_X1 U4052 ( .B1(n4157), .B2(n4158), .A(n4678), .ZN(n4171) );
  INV_X1 U4053 ( .A(n4679), .ZN(n4678) );
  OAI21_X1 U4054 ( .B1(n4158), .B2(n4157), .A(n4426), .ZN(n4679) );
  INV_X1 U4055 ( .A(n4104), .ZN(n4426) );
  XNOR2_X1 U4056 ( .A(\unit_decode/IMMreg/ffi_3/n4 ), .B(n3785), .ZN(n4158) );
  OAI21_X1 U4057 ( .B1(n4117), .B2(n4116), .A(n4680), .ZN(n4157) );
  OAI21_X1 U4058 ( .B1(n4122), .B2(n4681), .A(n4680), .ZN(n4116) );
  NAND2_X1 U4059 ( .A1(n4122), .A2(n4681), .ZN(n4680) );
  AND2_X1 U4060 ( .A1(n4682), .A2(n4683), .ZN(n4117) );
  INV_X1 U4061 ( .A(n4173), .ZN(n4677) );
  NOR2_X1 U4062 ( .A1(n4168), .A2(n4174), .ZN(n4173) );
  AOI21_X1 U4063 ( .B1(n3787), .B2(n4862), .A(n4684), .ZN(n4174) );
  INV_X1 U4064 ( .A(n4676), .ZN(n4210) );
  NOR2_X1 U4065 ( .A1(n4183), .A2(n4675), .ZN(n4676) );
  XNOR2_X1 U4066 ( .A(\unit_decode/IMMreg/ffi_5/n4 ), .B(n4862), .ZN(n4675) );
  XNOR2_X1 U4067 ( .A(\unit_decode/IMMreg/ffi_6/n4 ), .B(n3785), .ZN(n4674) );
  INV_X1 U4068 ( .A(n4198), .ZN(n4483) );
  INV_X1 U4069 ( .A(n4685), .ZN(n4241) );
  OAI21_X1 U4070 ( .B1(n4293), .B2(n4236), .A(n4290), .ZN(n4685) );
  NAND2_X1 U4071 ( .A1(n4293), .A2(n4236), .ZN(n4290) );
  INV_X1 U4072 ( .A(n4237), .ZN(n4236) );
  XOR2_X1 U4073 ( .A(\unit_decode/IMMreg/ffi_8/n4 ), .B(n4862), .Z(n4293) );
  AOI21_X1 U4074 ( .B1(n4686), .B2(n4268), .A(n4289), .ZN(n4275) );
  NOR2_X1 U4075 ( .A1(n4686), .A2(n4268), .ZN(n4289) );
  XNOR2_X1 U4076 ( .A(\unit_decode/IMMreg/ffi_10/n4 ), .B(n4862), .ZN(n4686)
         );
  XOR2_X1 U4077 ( .A(\unit_decode/IMMreg/ffi_11/n4 ), .B(n3785), .Z(n4668) );
  MUX2_X1 U4078 ( .A(\unit_decode/Areg/ffi_11/n4 ), .B(
        \unit_decode/NPC1reg/ffi_11/n4 ), .S(n4012), .Z(n4285) );
  XNOR2_X1 U4079 ( .A(\unit_decode/IMMreg/ffi_15/n4 ), .B(n4862), .ZN(n4663)
         );
  AOI21_X1 U4080 ( .B1(n4435), .B2(n4369), .A(n4660), .ZN(n4372) );
  NOR2_X1 U4081 ( .A1(n4435), .A2(n4369), .ZN(n4660) );
  XNOR2_X1 U4082 ( .A(\unit_decode/IMMreg/ffi_16/n4 ), .B(n4862), .ZN(n4435)
         );
  XOR2_X1 U4083 ( .A(\unit_decode/IMMreg/ffi_19/n4 ), .B(n3785), .Z(n4656) );
  MUX2_X1 U4084 ( .A(\unit_decode/Areg/ffi_19/n4 ), .B(
        \unit_decode/NPC1reg/ffi_19/n4 ), .S(n4012), .Z(n4422) );
  AND2_X1 U4085 ( .A1(n4504), .A2(n4468), .ZN(n4448) );
  NAND2_X1 U4086 ( .A1(n4444), .A2(n4687), .ZN(n4468) );
  OR2_X1 U4087 ( .A1(n4687), .A2(n4444), .ZN(n4504) );
  INV_X1 U4088 ( .A(n4445), .ZN(n4444) );
  MUX2_X1 U4089 ( .A(\unit_decode/Areg/ffi_20/n4 ), .B(
        \unit_decode/NPC1reg/ffi_20/n4 ), .S(n4012), .Z(n4445) );
  XNOR2_X1 U4090 ( .A(\unit_decode/IMMreg/ffi_20/n4 ), .B(n3785), .ZN(n4687)
         );
  INV_X1 U4091 ( .A(n4465), .ZN(n4467) );
  XOR2_X1 U4092 ( .A(n4460), .B(n4655), .Z(n4465) );
  XNOR2_X1 U4093 ( .A(\unit_decode/IMMreg/ffi_21/n4 ), .B(n3785), .ZN(n4655)
         );
  INV_X1 U4094 ( .A(n4461), .ZN(n4460) );
  MUX2_X1 U4095 ( .A(\unit_decode/Areg/ffi_21/n4 ), .B(
        \unit_decode/NPC1reg/ffi_21/n4 ), .S(n4012), .Z(n4461) );
  AOI21_X1 U4096 ( .B1(n4480), .B2(n4688), .A(n4501), .ZN(n4485) );
  NOR2_X1 U4097 ( .A1(n4480), .A2(n4688), .ZN(n4501) );
  XNOR2_X1 U4098 ( .A(\unit_decode/IMMreg/ffi_22/n4 ), .B(n4862), .ZN(n4688)
         );
  MUX2_X1 U4099 ( .A(\unit_decode/Areg/ffi_22/n4 ), .B(
        \unit_decode/NPC1reg/ffi_22/n4 ), .S(n4012), .Z(n4480) );
  XNOR2_X1 U4100 ( .A(\unit_decode/IMMreg/ffi_23/n4 ), .B(n3785), .ZN(n4651)
         );
  INV_X1 U4101 ( .A(n4496), .ZN(n4495) );
  NOR2_X1 U4102 ( .A1(n4650), .A2(n4513), .ZN(n4524) );
  INV_X1 U4103 ( .A(n4514), .ZN(n4513) );
  XNOR2_X1 U4104 ( .A(\unit_decode/IMMreg/ffi_24/n4 ), .B(n3785), .ZN(n4650)
         );
  XOR2_X1 U4105 ( .A(\unit_decode/IMMreg/ffi_26/n4 ), .B(n3785), .Z(n4645) );
  XNOR2_X1 U4106 ( .A(\unit_decode/IMMreg/ffi_27/n4 ), .B(n3785), .ZN(n4567)
         );
  OAI211_X1 U4107 ( .C1(n4496), .C2(n4272), .A(n4516), .B(n4689), .ZN(n4505)
         );
  AOI222_X1 U4108 ( .A1(n4518), .A2(n4220), .B1(n4519), .B2(n4619), .C1(n4376), 
        .C2(n4350), .ZN(n4689) );
  INV_X1 U4109 ( .A(n4351), .ZN(n4350) );
  MUX2_X1 U4110 ( .A(\unit_decode/Areg/ffi_15/n4 ), .B(
        \unit_decode/NPC1reg/ffi_15/n4 ), .S(n4012), .Z(n4351) );
  INV_X1 U4111 ( .A(n4097), .ZN(n4619) );
  NOR2_X1 U4112 ( .A1(n4166), .A2(n3778), .ZN(n4519) );
  INV_X1 U4113 ( .A(n4684), .ZN(n4166) );
  INV_X1 U4114 ( .A(n4221), .ZN(n4220) );
  INV_X1 U4115 ( .A(n4621), .ZN(n4518) );
  AOI21_X1 U4116 ( .B1(n3778), .B2(n4624), .A(n4378), .ZN(n4516) );
  MUX2_X1 U4117 ( .A(\unit_decode/Areg/ffi_23/n4 ), .B(
        \unit_decode/NPC1reg/ffi_23/n4 ), .S(n4012), .Z(n4496) );
  AOI222_X1 U4118 ( .A1(n4120), .A2(n4543), .B1(n4177), .B2(n4525), .C1(n4118), 
        .C2(n4539), .ZN(n4612) );
  OAI221_X1 U4119 ( .B1(n4252), .B2(n4621), .C1(n4534), .C2(n4272), .A(n4690), 
        .ZN(n4539) );
  AOI221_X1 U4120 ( .B1(n4623), .B2(n4389), .C1(n4376), .C2(n4386), .A(n4624), 
        .ZN(n4690) );
  INV_X1 U4121 ( .A(n4387), .ZN(n4386) );
  MUX2_X1 U4122 ( .A(\unit_decode/Areg/ffi_17/n4 ), .B(
        \unit_decode/NPC1reg/ffi_17/n4 ), .S(n4012), .Z(n4387) );
  MUX2_X1 U4123 ( .A(\unit_decode/Areg/ffi_25/n4 ), .B(
        \unit_decode/NPC1reg/ffi_25/n4 ), .S(n4012), .Z(n4534) );
  OAI221_X1 U4124 ( .B1(n4237), .B2(n4621), .C1(n4514), .C2(n4272), .A(n4691), 
        .ZN(n4525) );
  AOI221_X1 U4125 ( .B1(n4623), .B2(n4377), .C1(n4376), .C2(n4368), .A(n4624), 
        .ZN(n4691) );
  INV_X1 U4126 ( .A(n4369), .ZN(n4368) );
  MUX2_X1 U4127 ( .A(\unit_decode/Areg/ffi_16/n4 ), .B(
        \unit_decode/NPC1reg/ffi_16/n4 ), .S(n4012), .Z(n4369) );
  INV_X1 U4128 ( .A(n4023), .ZN(n4377) );
  MUX2_X1 U4129 ( .A(\unit_decode/Areg/ffi_24/n4 ), .B(
        \unit_decode/NPC1reg/ffi_24/n4 ), .S(n4012), .Z(n4514) );
  OAI221_X1 U4130 ( .B1(n4268), .B2(n4621), .C1(n4549), .C2(n4272), .A(n4692), 
        .ZN(n4543) );
  AOI221_X1 U4131 ( .B1(n4623), .B2(n4122), .C1(n4376), .C2(n4403), .A(n4624), 
        .ZN(n4692) );
  INV_X1 U4132 ( .A(n4404), .ZN(n4403) );
  MUX2_X1 U4133 ( .A(\unit_decode/Areg/ffi_18/n4 ), .B(
        \unit_decode/NPC1reg/ffi_18/n4 ), .S(n4012), .Z(n4404) );
  INV_X1 U4134 ( .A(n4634), .ZN(n4376) );
  NAND3_X1 U4135 ( .A1(\unit_decode/IMMreg/ffi_4/n4 ), .A2(n3778), .A3(n4693), 
        .ZN(n4634) );
  INV_X1 U4136 ( .A(n4102), .ZN(n4122) );
  INV_X1 U4137 ( .A(n4633), .ZN(n4623) );
  NAND3_X1 U4138 ( .A1(n3778), .A2(n3787), .A3(n4693), .ZN(n4633) );
  MUX2_X1 U4139 ( .A(\unit_decode/Areg/ffi_26/n4 ), .B(
        \unit_decode/NPC1reg/ffi_26/n4 ), .S(n4012), .Z(n4549) );
  NAND3_X1 U4140 ( .A1(\unit_decode/IMMreg/ffi_3/n4 ), .A2(n3787), .A3(n4693), 
        .ZN(n4621) );
  MUX2_X1 U4141 ( .A(\unit_decode/Areg/ffi_10/n4 ), .B(
        \unit_decode/NPC1reg/ffi_10/n4 ), .S(n4012), .Z(n4268) );
  NOR2_X1 U4142 ( .A1(\unit_decode/NPC1reg/ffi_0/n4 ), .A2(RST), .ZN(n4936) );
  NOR2_X1 U4143 ( .A1(\unit_decode/NPC1reg/ffi_1/n4 ), .A2(RST), .ZN(n4937) );
  NOR2_X1 U4144 ( .A1(\unit_decode/NPC1reg/ffi_2/n4 ), .A2(RST), .ZN(n4938) );
  NOR2_X1 U4145 ( .A1(\unit_decode/NPC1reg/ffi_3/n4 ), .A2(RST), .ZN(n4939) );
  NOR2_X1 U4146 ( .A1(\unit_decode/NPC1reg/ffi_4/n4 ), .A2(RST), .ZN(n4940) );
  NOR2_X1 U4147 ( .A1(\unit_decode/NPC1reg/ffi_5/n4 ), .A2(RST), .ZN(n4941) );
  NOR2_X1 U4148 ( .A1(\unit_decode/NPC1reg/ffi_6/n4 ), .A2(RST), .ZN(n4942) );
  NOR2_X1 U4149 ( .A1(\unit_decode/NPC1reg/ffi_7/n4 ), .A2(RST), .ZN(n4943) );
  NOR2_X1 U4150 ( .A1(\unit_decode/NPC1reg/ffi_8/n4 ), .A2(RST), .ZN(n4944) );
  NOR2_X1 U4151 ( .A1(\unit_decode/NPC1reg/ffi_9/n4 ), .A2(RST), .ZN(n4945) );
  NOR2_X1 U4152 ( .A1(\unit_decode/NPC1reg/ffi_10/n4 ), .A2(RST), .ZN(n4946)
         );
  NOR2_X1 U4153 ( .A1(\unit_decode/NPC1reg/ffi_11/n4 ), .A2(RST), .ZN(n4947)
         );
  NOR2_X1 U4154 ( .A1(\unit_decode/NPC1reg/ffi_12/n4 ), .A2(RST), .ZN(n4948)
         );
  NOR2_X1 U4155 ( .A1(\unit_decode/NPC1reg/ffi_13/n4 ), .A2(RST), .ZN(n4949)
         );
  NOR2_X1 U4156 ( .A1(\unit_decode/NPC1reg/ffi_14/n4 ), .A2(RST), .ZN(n4950)
         );
  NOR2_X1 U4157 ( .A1(\unit_decode/NPC1reg/ffi_15/n4 ), .A2(RST), .ZN(n4951)
         );
  NOR2_X1 U4158 ( .A1(\unit_decode/NPC1reg/ffi_16/n4 ), .A2(RST), .ZN(n4952)
         );
  NOR2_X1 U4159 ( .A1(\unit_decode/NPC1reg/ffi_17/n4 ), .A2(RST), .ZN(n4953)
         );
  NOR2_X1 U4160 ( .A1(\unit_decode/NPC1reg/ffi_18/n4 ), .A2(RST), .ZN(n4954)
         );
  NOR2_X1 U4161 ( .A1(\unit_decode/NPC1reg/ffi_19/n4 ), .A2(RST), .ZN(n4955)
         );
  NOR2_X1 U4162 ( .A1(\unit_decode/NPC1reg/ffi_20/n4 ), .A2(RST), .ZN(n4956)
         );
  NOR2_X1 U4163 ( .A1(\unit_decode/NPC1reg/ffi_21/n4 ), .A2(RST), .ZN(n4957)
         );
  NOR2_X1 U4164 ( .A1(\unit_decode/NPC1reg/ffi_22/n4 ), .A2(RST), .ZN(n4958)
         );
  NOR2_X1 U4165 ( .A1(\unit_decode/NPC1reg/ffi_23/n4 ), .A2(RST), .ZN(n4959)
         );
  NOR2_X1 U4166 ( .A1(\unit_decode/NPC1reg/ffi_24/n4 ), .A2(RST), .ZN(n4960)
         );
  NOR2_X1 U4167 ( .A1(\unit_decode/NPC1reg/ffi_25/n4 ), .A2(RST), .ZN(n4961)
         );
  NOR2_X1 U4168 ( .A1(\unit_decode/NPC1reg/ffi_26/n4 ), .A2(RST), .ZN(n4962)
         );
  NOR2_X1 U4169 ( .A1(\unit_decode/NPC1reg/ffi_27/n4 ), .A2(RST), .ZN(n4963)
         );
  NOR2_X1 U4170 ( .A1(\unit_decode/NPC1reg/ffi_28/n4 ), .A2(RST), .ZN(n4964)
         );
  NOR2_X1 U4171 ( .A1(\unit_decode/NPC1reg/ffi_29/n4 ), .A2(RST), .ZN(n4965)
         );
  NOR2_X1 U4172 ( .A1(\unit_decode/NPC1reg/ffi_30/n4 ), .A2(RST), .ZN(n4966)
         );
  NOR2_X1 U4173 ( .A1(\unit_decode/NPC1reg/ffi_31/n4 ), .A2(RST), .ZN(n4967)
         );
  NOR2_X1 U4174 ( .A1(RST), .A2(n3915), .ZN(n4968) );
  AND3_X1 U4175 ( .A1(n4694), .A2(n4695), .A3(n4696), .ZN(n3915) );
  AOI221_X1 U4176 ( .B1(n4017), .B2(n4119), .C1(n4697), .C2(n4106), .A(n4698), 
        .ZN(n4696) );
  OAI21_X1 U4177 ( .B1(n4105), .B2(n4155), .A(n4699), .ZN(n4698) );
  MUX2_X1 U4178 ( .A(n4700), .B(n4701), .S(n3781), .Z(n4699) );
  MUX2_X1 U4179 ( .A(n4025), .B(n4133), .S(n4100), .Z(n4701) );
  INV_X1 U4180 ( .A(n4036), .ZN(n4133) );
  INV_X1 U4181 ( .A(n4126), .ZN(n4025) );
  NAND2_X1 U4182 ( .A1(n4134), .A2(n4100), .ZN(n4700) );
  NOR2_X1 U4183 ( .A1(n4165), .A2(n4862), .ZN(n4134) );
  OR2_X1 U4184 ( .A1(n4860), .A2(n4859), .ZN(n4165) );
  INV_X1 U4185 ( .A(n4029), .ZN(n4155) );
  NOR2_X1 U4186 ( .A1(n4168), .A2(n4862), .ZN(n4029) );
  MUX2_X1 U4187 ( .A(\unit_decode/Areg/ffi_4/n4 ), .B(
        \unit_decode/NPC1reg/ffi_4/n4 ), .S(n4012), .Z(n4168) );
  INV_X1 U4188 ( .A(n4120), .ZN(n4105) );
  NAND2_X1 U4189 ( .A1(n4702), .A2(n4703), .ZN(n4139) );
  MUX2_X1 U4190 ( .A(n4862), .B(\unit_decode/IMMreg/ffi_2/n4 ), .S(n3781), .Z(
        n4702) );
  NAND2_X1 U4191 ( .A1(n4859), .A2(n3795), .ZN(n4193) );
  INV_X1 U4192 ( .A(n4075), .ZN(n4697) );
  OAI21_X1 U4193 ( .B1(n4704), .B2(n4705), .A(n4683), .ZN(n4075) );
  NAND2_X1 U4194 ( .A1(n4704), .A2(n4705), .ZN(n4683) );
  AOI21_X1 U4195 ( .B1(n4862), .B2(\unit_decode/IMMreg/ffi_0/n4 ), .A(n4035), 
        .ZN(n4705) );
  INV_X1 U4196 ( .A(n4109), .ZN(n4035) );
  NAND2_X1 U4197 ( .A1(n4023), .A2(n3786), .ZN(n4109) );
  INV_X1 U4198 ( .A(n4706), .ZN(n4704) );
  OAI21_X1 U4199 ( .B1(n4707), .B2(n4389), .A(n4682), .ZN(n4706) );
  NAND2_X1 U4200 ( .A1(n4707), .A2(n4389), .ZN(n4682) );
  INV_X1 U4201 ( .A(n4100), .ZN(n4389) );
  AOI21_X1 U4202 ( .B1(n4862), .B2(\unit_decode/IMMreg/ffi_1/n4 ), .A(n4708), 
        .ZN(n4707) );
  OAI221_X1 U4203 ( .B1(n4271), .B2(n4252), .C1(n4100), .C2(n4272), .A(n4273), 
        .ZN(n4119) );
  MUX2_X1 U4204 ( .A(\unit_decode/Areg/ffi_9/n4 ), .B(
        \unit_decode/NPC1reg/ffi_9/n4 ), .S(n4012), .Z(n4252) );
  NAND2_X1 U4205 ( .A1(n4709), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .ZN(n4151)
         );
  AOI222_X1 U4206 ( .A1(n4033), .A2(n4028), .B1(n4710), .B2(n3785), .C1(n4031), 
        .C2(n4108), .ZN(n4695) );
  NOR2_X1 U4207 ( .A1(n4146), .A2(n4201), .ZN(n4108) );
  OR3_X1 U4208 ( .A1(n4681), .A2(\unit_decode/IMMreg/ffi_1/n4 ), .A3(n3786), 
        .ZN(n4146) );
  NOR2_X1 U4209 ( .A1(n4221), .A2(n4862), .ZN(n4031) );
  MUX2_X1 U4210 ( .A(\unit_decode/Areg/ffi_7/n4 ), .B(
        \unit_decode/NPC1reg/ffi_7/n4 ), .S(n4012), .Z(n4221) );
  OAI222_X1 U4211 ( .A1(n4100), .A2(n4026), .B1(n4102), .B2(n4101), .C1(n4104), 
        .C2(n4103), .ZN(n4710) );
  INV_X1 U4212 ( .A(n4118), .ZN(n4103) );
  NAND3_X1 U4213 ( .A1(n4681), .A2(n3781), .A3(\unit_decode/IMMreg/ffi_0/n4 ), 
        .ZN(n4147) );
  XNOR2_X1 U4214 ( .A(\unit_decode/IMMreg/ffi_2/n4 ), .B(n3785), .ZN(n4681) );
  MUX2_X1 U4215 ( .A(\unit_decode/Areg/ffi_3/n4 ), .B(
        \unit_decode/NPC1reg/ffi_3/n4 ), .S(n4012), .Z(n4104) );
  INV_X1 U4216 ( .A(n4177), .ZN(n4101) );
  NAND2_X1 U4217 ( .A1(n4711), .A2(n4703), .ZN(n4154) );
  AOI21_X1 U4218 ( .B1(n4862), .B2(\unit_decode/IMMreg/ffi_2/n4 ), .A(
        \unit_decode/IMMreg/ffi_0/n4 ), .ZN(n4703) );
  MUX2_X1 U4219 ( .A(n3781), .B(n4712), .S(n3785), .Z(n4711) );
  MUX2_X1 U4220 ( .A(\unit_decode/Areg/ffi_2/n4 ), .B(
        \unit_decode/NPC1reg/ffi_2/n4 ), .S(n4012), .Z(n4102) );
  INV_X1 U4221 ( .A(n4121), .ZN(n4026) );
  NAND3_X1 U4222 ( .A1(\unit_decode/IMMreg/ffi_0/n4 ), .A2(n3785), .A3(n4712), 
        .ZN(n4149) );
  MUX2_X1 U4223 ( .A(\unit_decode/Areg/ffi_1/n4 ), .B(
        \unit_decode/NPC1reg/ffi_1/n4 ), .S(n4012), .Z(n4100) );
  NAND3_X1 U4224 ( .A1(\unit_decode/IMMreg/ffi_1/n4 ), .A2(n3790), .A3(
        \unit_decode/IMMreg/ffi_0/n4 ), .ZN(n4143) );
  NOR2_X1 U4225 ( .A1(n4183), .A2(n4862), .ZN(n4033) );
  MUX2_X1 U4226 ( .A(\unit_decode/Areg/ffi_5/n4 ), .B(
        \unit_decode/NPC1reg/ffi_5/n4 ), .S(n4012), .Z(n4183) );
  AOI22_X1 U4227 ( .A1(n4030), .A2(n4018), .B1(n4107), .B2(n4032), .ZN(n4694)
         );
  NOR2_X1 U4228 ( .A1(n4142), .A2(n4201), .ZN(n4032) );
  NAND3_X1 U4229 ( .A1(n4630), .A2(n3786), .A3(n4713), .ZN(n4142) );
  AOI21_X1 U4230 ( .B1(n4862), .B2(n3790), .A(n4708), .ZN(n4713) );
  NOR2_X1 U4231 ( .A1(n4198), .A2(n4862), .ZN(n4107) );
  MUX2_X1 U4232 ( .A(\unit_decode/Areg/ffi_6/n4 ), .B(
        \unit_decode/NPC1reg/ffi_6/n4 ), .S(n4012), .Z(n4198) );
  OAI221_X1 U4233 ( .B1(n4271), .B2(n4237), .C1(n4023), .C2(n4272), .A(n4273), 
        .ZN(n4018) );
  NAND2_X1 U4234 ( .A1(n4378), .A2(n3778), .ZN(n4273) );
  AND2_X1 U4235 ( .A1(n4624), .A2(n3787), .ZN(n4378) );
  MUX2_X1 U4236 ( .A(\unit_decode/Areg/ffi_31/n4 ), .B(
        \unit_decode/NPC1reg/ffi_31/n4 ), .S(n4012), .Z(n4097) );
  AND2_X1 U4237 ( .A1(n4861), .A2(n4862), .ZN(n4693) );
  MUX2_X1 U4238 ( .A(\unit_decode/Areg/ffi_0/n4 ), .B(
        \unit_decode/NPC1reg/ffi_0/n4 ), .S(n4012), .Z(n4023) );
  MUX2_X1 U4239 ( .A(\unit_decode/Areg/ffi_8/n4 ), .B(
        \unit_decode/NPC1reg/ffi_8/n4 ), .S(n4012), .Z(n4237) );
  AOI21_X1 U4240 ( .B1(n3785), .B2(\unit_decode/IMMreg/ffi_3/n4 ), .A(n4684), 
        .ZN(n4271) );
  NOR2_X1 U4241 ( .A1(n3787), .A2(n4862), .ZN(n4684) );
  NAND2_X1 U4242 ( .A1(n4860), .A2(n4859), .ZN(n4201) );
  OAI21_X1 U4243 ( .B1(n4709), .B2(n4714), .A(n3786), .ZN(n4153) );
  AND2_X1 U4244 ( .A1(n3790), .A2(n4708), .ZN(n4714) );
  NOR2_X1 U4245 ( .A1(\unit_decode/IMMreg/ffi_1/n4 ), .A2(n4862), .ZN(n4708)
         );
  NOR2_X1 U4246 ( .A1(n4630), .A2(n3785), .ZN(n4709) );
  INV_X1 U4247 ( .A(n4712), .ZN(n4630) );
  NOR2_X1 U4248 ( .A1(n3781), .A2(n3790), .ZN(n4712) );
  NOR2_X1 U4249 ( .A1(RST), .A2(n4715), .ZN(n4971) );
  NOR2_X1 U4250 ( .A1(RST), .A2(n4716), .ZN(n4972) );
  NOR2_X1 U4251 ( .A1(RST), .A2(n4717), .ZN(n4973) );
  NOR2_X1 U4252 ( .A1(RST), .A2(n4718), .ZN(n4974) );
  NOR2_X1 U4253 ( .A1(RST), .A2(n4719), .ZN(n4975) );
  NOR2_X1 U4254 ( .A1(\unit_fetch/unit_instructionRegister/n38 ), .A2(RST), 
        .ZN(n4976) );
  NOR2_X1 U4255 ( .A1(\unit_fetch/unit_instructionRegister/n39 ), .A2(RST), 
        .ZN(n4977) );
  NOR2_X1 U4256 ( .A1(\unit_fetch/unit_instructionRegister/n40 ), .A2(RST), 
        .ZN(n4978) );
  NOR2_X1 U4257 ( .A1(\unit_fetch/unit_instructionRegister/n41 ), .A2(RST), 
        .ZN(n4979) );
  NOR2_X1 U4258 ( .A1(\unit_fetch/unit_instructionRegister/n43 ), .A2(RST), 
        .ZN(n4980) );
  NOR2_X1 U4259 ( .A1(\unit_fetch/unit_instructionRegister/n44 ), .A2(RST), 
        .ZN(n4981) );
  NOR2_X1 U4260 ( .A1(\unit_fetch/unit_instructionRegister/n45 ), .A2(RST), 
        .ZN(n4982) );
  NOR2_X1 U4261 ( .A1(\unit_fetch/unit_instructionRegister/n46 ), .A2(RST), 
        .ZN(n4983) );
  NOR2_X1 U4262 ( .A1(\unit_fetch/unit_instructionRegister/n47 ), .A2(RST), 
        .ZN(n4984) );
  NOR2_X1 U4263 ( .A1(\unit_fetch/unit_instructionRegister/n48 ), .A2(RST), 
        .ZN(n4985) );
  NOR2_X1 U4264 ( .A1(\unit_fetch/unit_instructionRegister/n49 ), .A2(RST), 
        .ZN(n4986) );
  NOR2_X1 U4265 ( .A1(\unit_fetch/unit_instructionRegister/n51 ), .A2(RST), 
        .ZN(n4987) );
  NOR2_X1 U4266 ( .A1(\unit_fetch/unit_instructionRegister/n52 ), .A2(RST), 
        .ZN(n4988) );
  OAI21_X1 U4267 ( .B1(\unit_fetch/unit_instructionRegister/n54 ), .B2(n4720), 
        .A(n4721), .ZN(n4990) );
  OAI21_X1 U4268 ( .B1(\unit_fetch/unit_instructionRegister/n55 ), .B2(n4720), 
        .A(n4721), .ZN(n4991) );
  OAI21_X1 U4269 ( .B1(\unit_fetch/unit_instructionRegister/n56 ), .B2(n4720), 
        .A(n4721), .ZN(n4992) );
  OAI21_X1 U4270 ( .B1(\unit_fetch/unit_instructionRegister/n57 ), .B2(n4720), 
        .A(n4721), .ZN(n4993) );
  OAI21_X1 U4271 ( .B1(\unit_fetch/unit_instructionRegister/n59 ), .B2(n4720), 
        .A(n4721), .ZN(n4995) );
  NAND2_X1 U4272 ( .A1(n4722), .A2(n4723), .ZN(n4994) );
  OR3_X1 U4273 ( .A1(n1337), .A2(\unit_fetch/unit_instructionRegister/n60 ), 
        .A3(n4720), .ZN(n4723) );
  OAI21_X1 U4274 ( .B1(\unit_fetch/unit_instructionRegister/n61 ), .B2(n4720), 
        .A(n4721), .ZN(n4996) );
  OAI21_X1 U4275 ( .B1(\unit_fetch/unit_instructionRegister/n62 ), .B2(n4720), 
        .A(n4721), .ZN(n4997) );
  OAI21_X1 U4276 ( .B1(\unit_fetch/unit_instructionRegister/n63 ), .B2(n4720), 
        .A(n4721), .ZN(n4998) );
  NAND4_X1 U4277 ( .A1(n4864), .A2(n2912), .A3(n3776), .A4(n3799), .ZN(n4721)
         );
  INV_X1 U4278 ( .A(\unit_control/uut_third_stage/ffi_15/n5 ), .ZN(n4720) );
  NAND2_X1 U4279 ( .A1(n4722), .A2(n4724), .ZN(n4999) );
  NAND4_X1 U4280 ( .A1(n4864), .A2(\unit_control/uut_third_stage/ffi_15/n5 ), 
        .A3(\cw_dec[2] ), .A4(\unit_decode/RS1s[4] ), .ZN(n4724) );
  NOR2_X1 U4281 ( .A1(n3776), .A2(RST), .ZN(
        \unit_control/uut_third_stage/ffi_15/n5 ) );
  NAND4_X1 U4282 ( .A1(n4989), .A2(n4864), .A3(\cw_dec[2] ), .A4(n3776), .ZN(
        n4722) );
  NOR2_X1 U4283 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n53 ), 
        .ZN(n4989) );
  AND2_X1 U4284 ( .A1(\unit_decode/registerA[0] ), .A2(n2912), .ZN(n5000) );
  AND2_X1 U4285 ( .A1(\unit_decode/registerA[1] ), .A2(n2912), .ZN(n5001) );
  AND2_X1 U4286 ( .A1(\unit_decode/registerA[2] ), .A2(n2912), .ZN(n5002) );
  AND2_X1 U4287 ( .A1(\unit_decode/registerA[3] ), .A2(n2912), .ZN(n5003) );
  AND2_X1 U4288 ( .A1(\unit_decode/registerA[4] ), .A2(n2912), .ZN(n5004) );
  AND2_X1 U4289 ( .A1(\unit_decode/registerA[5] ), .A2(n2912), .ZN(n5005) );
  AND2_X1 U4290 ( .A1(\unit_decode/registerA[6] ), .A2(n2912), .ZN(n5006) );
  AND2_X1 U4291 ( .A1(\unit_decode/registerA[7] ), .A2(n2912), .ZN(n5007) );
  AND2_X1 U4292 ( .A1(\unit_decode/registerA[8] ), .A2(n2912), .ZN(n5008) );
  AND2_X1 U4293 ( .A1(\unit_decode/registerA[9] ), .A2(n2912), .ZN(n5009) );
  AND2_X1 U4294 ( .A1(\unit_decode/registerA[10] ), .A2(n2912), .ZN(n5010) );
  AND2_X1 U4295 ( .A1(\unit_decode/registerA[11] ), .A2(n2912), .ZN(n5011) );
  AND2_X1 U4296 ( .A1(\unit_decode/registerA[12] ), .A2(n2912), .ZN(n5012) );
  AND2_X1 U4297 ( .A1(\unit_decode/registerA[13] ), .A2(n2912), .ZN(n5013) );
  AND2_X1 U4298 ( .A1(\unit_decode/registerA[14] ), .A2(n2912), .ZN(n5014) );
  AND2_X1 U4299 ( .A1(\unit_decode/registerA[15] ), .A2(n2912), .ZN(n5015) );
  AND2_X1 U4300 ( .A1(\unit_decode/registerA[16] ), .A2(n2912), .ZN(n5016) );
  AND2_X1 U4301 ( .A1(\unit_decode/registerA[17] ), .A2(n2912), .ZN(n5017) );
  AND2_X1 U4302 ( .A1(\unit_decode/registerA[18] ), .A2(n2912), .ZN(n5018) );
  AND2_X1 U4303 ( .A1(\unit_decode/registerA[19] ), .A2(n2912), .ZN(n5019) );
  AND2_X1 U4304 ( .A1(\unit_decode/registerA[20] ), .A2(n2912), .ZN(n5020) );
  AND2_X1 U4305 ( .A1(\unit_decode/registerA[21] ), .A2(n2912), .ZN(n5021) );
  AND2_X1 U4306 ( .A1(\unit_decode/registerA[22] ), .A2(n2912), .ZN(n5022) );
  AND2_X1 U4307 ( .A1(\unit_decode/registerA[23] ), .A2(n2912), .ZN(n5023) );
  AND2_X1 U4308 ( .A1(\unit_decode/registerA[24] ), .A2(n2912), .ZN(n5024) );
  AND2_X1 U4309 ( .A1(\unit_decode/registerA[25] ), .A2(n2912), .ZN(n5025) );
  AND2_X1 U4310 ( .A1(\unit_decode/registerA[26] ), .A2(n2912), .ZN(n5026) );
  AND2_X1 U4311 ( .A1(\unit_decode/registerA[27] ), .A2(n2912), .ZN(n5027) );
  AND2_X1 U4312 ( .A1(\unit_decode/registerA[28] ), .A2(n2912), .ZN(n5028) );
  AND2_X1 U4313 ( .A1(\unit_decode/registerA[29] ), .A2(n2912), .ZN(n5029) );
  AND2_X1 U4314 ( .A1(\unit_decode/registerA[30] ), .A2(n2912), .ZN(n5030) );
  AND2_X1 U4315 ( .A1(\unit_decode/registerA[31] ), .A2(n2912), .ZN(n5031) );
  NOR2_X1 U4316 ( .A1(\unit_fetch/unit_npcregister/ffi_0/n4 ), .A2(RST), .ZN(
        n5032) );
  NOR2_X1 U4317 ( .A1(\unit_fetch/unit_npcregister/ffi_1/n4 ), .A2(RST), .ZN(
        n5033) );
  NOR2_X1 U4318 ( .A1(\unit_fetch/unit_npcregister/ffi_2/n4 ), .A2(RST), .ZN(
        n5034) );
  NOR2_X1 U4319 ( .A1(\unit_fetch/unit_npcregister/ffi_3/n4 ), .A2(RST), .ZN(
        n5035) );
  NOR2_X1 U4320 ( .A1(\unit_fetch/unit_npcregister/ffi_4/n4 ), .A2(RST), .ZN(
        n5036) );
  NOR2_X1 U4321 ( .A1(\unit_fetch/unit_npcregister/ffi_5/n4 ), .A2(RST), .ZN(
        n5037) );
  NOR2_X1 U4322 ( .A1(\unit_fetch/unit_npcregister/ffi_6/n4 ), .A2(RST), .ZN(
        n5038) );
  NOR2_X1 U4323 ( .A1(\unit_fetch/unit_npcregister/ffi_7/n4 ), .A2(RST), .ZN(
        n5039) );
  NOR2_X1 U4324 ( .A1(\unit_fetch/unit_npcregister/ffi_8/n4 ), .A2(RST), .ZN(
        n5040) );
  NOR2_X1 U4325 ( .A1(\unit_fetch/unit_npcregister/ffi_9/n4 ), .A2(RST), .ZN(
        n5041) );
  NOR2_X1 U4326 ( .A1(\unit_fetch/unit_npcregister/ffi_10/n4 ), .A2(RST), .ZN(
        n5042) );
  NOR2_X1 U4327 ( .A1(\unit_fetch/unit_npcregister/ffi_11/n4 ), .A2(RST), .ZN(
        n5043) );
  NOR2_X1 U4328 ( .A1(\unit_fetch/unit_npcregister/ffi_12/n4 ), .A2(RST), .ZN(
        n5044) );
  NOR2_X1 U4329 ( .A1(\unit_fetch/unit_npcregister/ffi_13/n4 ), .A2(RST), .ZN(
        n5045) );
  NOR2_X1 U4330 ( .A1(\unit_fetch/unit_npcregister/ffi_14/n4 ), .A2(RST), .ZN(
        n5046) );
  NOR2_X1 U4331 ( .A1(\unit_fetch/unit_npcregister/ffi_15/n4 ), .A2(RST), .ZN(
        n5047) );
  NOR2_X1 U4332 ( .A1(\unit_fetch/unit_npcregister/ffi_16/n4 ), .A2(RST), .ZN(
        n5048) );
  NOR2_X1 U4333 ( .A1(\unit_fetch/unit_npcregister/ffi_17/n4 ), .A2(RST), .ZN(
        n5049) );
  NOR2_X1 U4334 ( .A1(\unit_fetch/unit_npcregister/ffi_18/n4 ), .A2(RST), .ZN(
        n5050) );
  NOR2_X1 U4335 ( .A1(\unit_fetch/unit_npcregister/ffi_19/n4 ), .A2(RST), .ZN(
        n5051) );
  NOR2_X1 U4336 ( .A1(\unit_fetch/unit_npcregister/ffi_20/n4 ), .A2(RST), .ZN(
        n5052) );
  NOR2_X1 U4337 ( .A1(\unit_fetch/unit_npcregister/ffi_21/n4 ), .A2(RST), .ZN(
        n5053) );
  NOR2_X1 U4338 ( .A1(\unit_fetch/unit_npcregister/ffi_22/n4 ), .A2(RST), .ZN(
        n5054) );
  NOR2_X1 U4339 ( .A1(\unit_fetch/unit_npcregister/ffi_23/n4 ), .A2(RST), .ZN(
        n5055) );
  NOR2_X1 U4340 ( .A1(\unit_fetch/unit_npcregister/ffi_24/n4 ), .A2(RST), .ZN(
        n5056) );
  NOR2_X1 U4341 ( .A1(\unit_fetch/unit_npcregister/ffi_25/n4 ), .A2(RST), .ZN(
        n5057) );
  NOR2_X1 U4342 ( .A1(\unit_fetch/unit_npcregister/ffi_26/n4 ), .A2(RST), .ZN(
        n5058) );
  NOR2_X1 U4343 ( .A1(\unit_fetch/unit_npcregister/ffi_27/n4 ), .A2(RST), .ZN(
        n5059) );
  NOR2_X1 U4344 ( .A1(\unit_fetch/unit_npcregister/ffi_28/n4 ), .A2(RST), .ZN(
        n5060) );
  NOR2_X1 U4345 ( .A1(\unit_fetch/unit_npcregister/ffi_29/n4 ), .A2(RST), .ZN(
        n5061) );
  NOR2_X1 U4346 ( .A1(\unit_fetch/unit_npcregister/ffi_30/n4 ), .A2(RST), .ZN(
        n5062) );
  NOR2_X1 U4347 ( .A1(\unit_fetch/unit_npcregister/ffi_31/n4 ), .A2(RST), .ZN(
        n5063) );
  INV_X1 U4348 ( .A(n4725), .ZN(n3770) );
  AOI21_X1 U4349 ( .B1(n3825), .B2(n3839), .A(n2618), .ZN(n4725) );
  NOR3_X1 U4350 ( .A1(n3837), .A2(n3773), .A3(n3870), .ZN(n3839) );
  INV_X1 U4351 ( .A(n3880), .ZN(n3870) );
  NAND2_X1 U4352 ( .A1(n3899), .A2(n4726), .ZN(n3768) );
  NAND2_X1 U4353 ( .A1(n1337), .A2(n2912), .ZN(n3676) );
  NAND2_X1 U4354 ( .A1(\unit_control/uut_third_stage/ffi_17/n5 ), .A2(n2912), 
        .ZN(n3095) );
  INV_X1 U4355 ( .A(n3893), .ZN(n2621) );
  NAND2_X1 U4356 ( .A1(n4727), .A2(n3825), .ZN(n3893) );
  INV_X1 U4357 ( .A(n3899), .ZN(n2620) );
  NAND2_X1 U4358 ( .A1(n3825), .A2(n4728), .ZN(n3899) );
  INV_X1 U4359 ( .A(n3855), .ZN(n2619) );
  NAND2_X1 U4360 ( .A1(n3825), .A2(n4729), .ZN(n3855) );
  OAI21_X1 U4361 ( .B1(n3845), .B2(n3885), .A(n3846), .ZN(n4729) );
  AOI211_X1 U4362 ( .C1(n3878), .C2(n3853), .A(n3868), .B(n3874), .ZN(n3846)
         );
  INV_X1 U4363 ( .A(n4730), .ZN(n3874) );
  INV_X1 U4364 ( .A(n3890), .ZN(n3868) );
  NAND3_X1 U4365 ( .A1(\unit_fetch/pc_regout[3] ), .A2(n3883), .A3(n3884), 
        .ZN(n3890) );
  INV_X1 U4366 ( .A(n4731), .ZN(n3883) );
  INV_X1 U4367 ( .A(n3845), .ZN(n3853) );
  NAND2_X1 U4368 ( .A1(n3864), .A2(n3867), .ZN(n3878) );
  INV_X1 U4369 ( .A(n4732), .ZN(n2617) );
  AOI21_X1 U4370 ( .B1(n3869), .B2(n3825), .A(n2618), .ZN(n4732) );
  AND2_X1 U4371 ( .A1(n3825), .A2(n4733), .ZN(n2618) );
  OAI21_X1 U4372 ( .B1(n4734), .B2(n3845), .A(n4730), .ZN(n4733) );
  NAND2_X1 U4373 ( .A1(n3889), .A2(\unit_fetch/pc_regout[3] ), .ZN(n4730) );
  NOR3_X1 U4374 ( .A1(n3896), .A2(n3771), .A3(n3837), .ZN(n3889) );
  NAND2_X1 U4375 ( .A1(n3884), .A2(n3852), .ZN(n3837) );
  AND3_X1 U4376 ( .A1(n3860), .A2(n3885), .A3(n3867), .ZN(n4734) );
  INV_X1 U4377 ( .A(n3891), .ZN(n3860) );
  OAI21_X1 U4378 ( .B1(n3848), .B2(n3864), .A(n4735), .ZN(n3869) );
  NAND3_X1 U4379 ( .A1(n4736), .A2(n3852), .A3(n3880), .ZN(n4735) );
  NOR3_X1 U4380 ( .A1(n3771), .A2(\unit_fetch/unit_programCounter/ffi_0/n4 ), 
        .A3(n3788), .ZN(n3880) );
  NAND3_X1 U4381 ( .A1(n3771), .A2(n3779), .A3(
        \unit_fetch/unit_programCounter/ffi_1/n4 ), .ZN(n3864) );
  NAND2_X1 U4382 ( .A1(n4737), .A2(n4738), .ZN(n2600) );
  NAND3_X1 U4383 ( .A1(n3898), .A2(n3906), .A3(
        \unit_fetch/unit_instructionRegister/n72 ), .ZN(n4738) );
  INV_X1 U4384 ( .A(n3769), .ZN(n4737) );
  NOR2_X1 U4385 ( .A1(n4739), .A2(n3902), .ZN(n3769) );
  INV_X1 U4386 ( .A(\unit_fetch/unit_instructionRegister/n72 ), .ZN(n3902) );
  NOR2_X1 U4387 ( .A1(n3829), .A2(n3907), .ZN(
        \unit_fetch/unit_instructionRegister/n72 ) );
  INV_X1 U4388 ( .A(n3825), .ZN(n3829) );
  INV_X1 U4389 ( .A(n4726), .ZN(n2598) );
  NAND2_X1 U4390 ( .A1(n2599), .A2(n3906), .ZN(n4726) );
  OAI221_X1 U4391 ( .B1(n3780), .B2(n3885), .C1(n3789), .C2(n3896), .A(n4740), 
        .ZN(n3906) );
  AOI22_X1 U4392 ( .A1(n3897), .A2(n4741), .B1(n3884), .B2(
        \unit_fetch/pc_regout[2] ), .ZN(n4740) );
  NAND2_X1 U4393 ( .A1(\unit_fetch/pc_regout[2] ), .A2(n3788), .ZN(n4741) );
  INV_X1 U4394 ( .A(n3900), .ZN(n2599) );
  NAND3_X1 U4395 ( .A1(n3907), .A2(n3898), .A3(
        \unit_fetch/unit_instructionRegister/n73 ), .ZN(n3900) );
  INV_X1 U4396 ( .A(n3903), .ZN(\unit_fetch/unit_instructionRegister/n73 ) );
  NAND2_X1 U4397 ( .A1(n3825), .A2(n4739), .ZN(n3903) );
  NOR2_X1 U4398 ( .A1(n4742), .A2(\unit_control/n153 ), .ZN(n4013) );
  AOI211_X1 U4399 ( .C1(n3910), .C2(n4743), .A(n4744), .B(\unit_control/n152 ), 
        .ZN(n4742) );
  INV_X1 U4400 ( .A(n3911), .ZN(n4744) );
  NAND2_X1 U4401 ( .A1(n4743), .A2(n4745), .ZN(n3911) );
  NAND3_X1 U4402 ( .A1(\unit_decode/RD1reg/ffi_3/n4 ), .A2(
        \unit_decode/RD1reg/ffi_1/n4 ), .A3(\unit_decode/RD1reg/ffi_4/n4 ), 
        .ZN(n4745) );
  INV_X1 U4403 ( .A(n3909), .ZN(n4743) );
  NAND4_X1 U4404 ( .A1(n4728), .A2(n4746), .A3(n4747), .A4(n4748), .ZN(n3909)
         );
  AND4_X1 U4405 ( .A1(n4717), .A2(n4715), .A3(n4749), .A4(n4750), .ZN(n4748)
         );
  MUX2_X1 U4406 ( .A(n3894), .B(n4751), .S(n4718), .Z(n4750) );
  OAI21_X1 U4407 ( .B1(n3910), .B2(\unit_decode/RD1reg/ffi_3/n4 ), .A(n3894), 
        .ZN(n4751) );
  MUX2_X1 U4408 ( .A(n3895), .B(n4752), .S(n4719), .Z(n4749) );
  OAI21_X1 U4409 ( .B1(n3910), .B2(\unit_decode/RD1reg/ffi_4/n4 ), .A(n3895), 
        .ZN(n4752) );
  AND2_X1 U4410 ( .A1(n4753), .A2(n4754), .ZN(n4715) );
  MUX2_X1 U4411 ( .A(\unit_fetch/unit_instructionRegister/n49 ), .B(
        \unit_fetch/unit_instructionRegister/n54 ), .S(n4755), .Z(n4753) );
  AND2_X1 U4412 ( .A1(n4756), .A2(n4754), .ZN(n4717) );
  MUX2_X1 U4413 ( .A(\unit_fetch/unit_instructionRegister/n51 ), .B(
        \unit_fetch/unit_instructionRegister/n56 ), .S(n4755), .Z(n4756) );
  INV_X1 U4414 ( .A(n4757), .ZN(n4747) );
  OAI21_X1 U4415 ( .B1(n4758), .B2(n4716), .A(n2912), .ZN(n4757) );
  OAI21_X1 U4416 ( .B1(n4759), .B2(n4760), .A(n3908), .ZN(n4746) );
  INV_X1 U4417 ( .A(n3910), .ZN(n3908) );
  NAND2_X1 U4418 ( .A1(\unit_decode/RD1reg/ffi_2/n4 ), .A2(
        \unit_decode/RD1reg/ffi_0/n4 ), .ZN(n4760) );
  OAI222_X1 U4419 ( .A1(\unit_decode/RD1reg/ffi_4/n4 ), .A2(n3895), .B1(
        \unit_decode/RD1reg/ffi_3/n4 ), .B2(n3894), .C1(
        \unit_decode/RD1reg/ffi_1/n4 ), .C2(n4758), .ZN(n4759) );
  INV_X1 U4420 ( .A(n3892), .ZN(n4758) );
  NOR2_X1 U4421 ( .A1(n3881), .A2(n4727), .ZN(n3892) );
  AOI21_X1 U4422 ( .B1(n3788), .B2(n3885), .A(n3845), .ZN(n4727) );
  NAND3_X1 U4423 ( .A1(n3852), .A2(n3780), .A3(n3897), .ZN(n3845) );
  OAI22_X1 U4424 ( .A1(n3848), .A2(n3867), .B1(n4761), .B2(n4731), .ZN(n3881)
         );
  NAND3_X1 U4425 ( .A1(n3852), .A2(n3826), .A3(\unit_fetch/pc_regout[2] ), 
        .ZN(n4731) );
  NAND2_X1 U4426 ( .A1(n3826), .A2(n3771), .ZN(n3867) );
  OAI21_X1 U4427 ( .B1(n3851), .B2(n4762), .A(n3852), .ZN(n3848) );
  AND4_X1 U4428 ( .A1(n4763), .A2(n4764), .A3(n4765), .A4(n4766), .ZN(n3852)
         );
  NOR4_X1 U4429 ( .A1(n4767), .A2(\unit_fetch/pc_regout[28] ), .A3(
        \unit_fetch/pc_regout[30] ), .A4(\unit_fetch/pc_regout[29] ), .ZN(
        n4766) );
  NAND4_X1 U4430 ( .A1(n3797), .A2(n3784), .A3(n3772), .A4(n3777), .ZN(n4767)
         );
  NOR4_X1 U4431 ( .A1(n4768), .A2(\unit_fetch/pc_regout[25] ), .A3(
        \unit_fetch/pc_regout[27] ), .A4(\unit_fetch/pc_regout[26] ), .ZN(
        n4765) );
  NAND3_X1 U4432 ( .A1(n3794), .A2(n3782), .A3(n3775), .ZN(n4768) );
  NOR4_X1 U4433 ( .A1(n4769), .A2(\unit_fetch/pc_regout[18] ), .A3(
        \unit_fetch/pc_regout[20] ), .A4(\unit_fetch/pc_regout[19] ), .ZN(
        n4764) );
  NAND3_X1 U4434 ( .A1(n3796), .A2(n3774), .A3(n3783), .ZN(n4769) );
  NOR4_X1 U4435 ( .A1(n4770), .A2(\unit_fetch/pc_regout[10] ), .A3(
        \unit_fetch/pc_regout[13] ), .A4(\unit_fetch/pc_regout[12] ), .ZN(
        n4763) );
  NAND3_X1 U4436 ( .A1(n4855), .A2(n4856), .A3(n4854), .ZN(n4770) );
  NOR3_X1 U4437 ( .A1(n3780), .A2(\unit_fetch/pc_regout[4] ), .A3(
        \unit_fetch/pc_regout[3] ), .ZN(n4762) );
  NOR2_X1 U4438 ( .A1(n3773), .A2(n4761), .ZN(n3851) );
  INV_X1 U4439 ( .A(n4736), .ZN(n4761) );
  NOR2_X1 U4440 ( .A1(n3789), .A2(\unit_fetch/pc_regout[5] ), .ZN(n4736) );
  OAI21_X1 U4441 ( .B1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n4771), 
        .A(n4772), .ZN(n3894) );
  NAND2_X1 U4442 ( .A1(n4773), .A2(n4774), .ZN(n3895) );
  MUX2_X1 U4443 ( .A(n4775), .B(n4771), .S(n3788), .Z(n4773) );
  NOR2_X1 U4444 ( .A1(n3884), .A2(n4776), .ZN(n4771) );
  NOR3_X1 U4445 ( .A1(\unit_fetch/pc_regout[3] ), .A2(
        \unit_fetch/pc_regout[5] ), .A3(\unit_fetch/pc_regout[2] ), .ZN(n4776)
         );
  NOR2_X1 U4446 ( .A1(\unit_fetch/pc_regout[4] ), .A2(
        \unit_fetch/pc_regout[5] ), .ZN(n3884) );
  NAND2_X1 U4447 ( .A1(n3897), .A2(\unit_fetch/pc_regout[2] ), .ZN(n4775) );
  XOR2_X1 U4448 ( .A(n4777), .B(n3907), .Z(n4728) );
  NAND2_X1 U4449 ( .A1(n3901), .A2(n4739), .ZN(n4777) );
  NAND3_X1 U4450 ( .A1(n4778), .A2(n4774), .A3(n4772), .ZN(n4739) );
  NAND2_X1 U4451 ( .A1(n4779), .A2(n3897), .ZN(n4772) );
  XNOR2_X1 U4452 ( .A(\unit_fetch/unit_programCounter/ffi_1/n4 ), .B(
        \unit_fetch/pc_regout[2] ), .ZN(n4779) );
  NAND3_X1 U4453 ( .A1(n3771), .A2(n3779), .A3(n3897), .ZN(n4774) );
  INV_X1 U4454 ( .A(n3922), .ZN(n4778) );
  NAND3_X1 U4455 ( .A1(n4719), .A2(n4718), .A3(n4716), .ZN(n3910) );
  AOI21_X1 U4456 ( .B1(n3800), .B2(n4755), .A(n4780), .ZN(n4716) );
  AOI21_X1 U4457 ( .B1(n3801), .B2(n4755), .A(n4780), .ZN(n4718) );
  OAI21_X1 U4458 ( .B1(\unit_fetch/unit_instructionRegister/n52 ), .B2(n4755), 
        .A(n4754), .ZN(n4780) );
  AND2_X1 U4459 ( .A1(n4781), .A2(n4754), .ZN(n4719) );
  NAND4_X1 U4460 ( .A1(\unit_fetch/unit_instructionRegister/n66 ), .A2(
        \unit_fetch/unit_instructionRegister/n65 ), .A3(n4782), .A4(n3798), 
        .ZN(n4754) );
  NOR2_X1 U4461 ( .A1(\unit_fetch/unit_instructionRegister/n64 ), .A2(n4863), 
        .ZN(n4782) );
  MUX2_X1 U4462 ( .A(\unit_fetch/unit_instructionRegister/n53 ), .B(
        \unit_fetch/unit_instructionRegister/n60 ), .S(n4755), .Z(n4781) );
  NAND4_X1 U4463 ( .A1(\unit_fetch/unit_instructionRegister/n65 ), .A2(n3798), 
        .A3(\unit_fetch/unit_instructionRegister/n66 ), .A4(n4783), .ZN(n4755)
         );
  AND2_X1 U4464 ( .A1(n4863), .A2(\unit_fetch/unit_instructionRegister/n64 ), 
        .ZN(n4783) );
  INV_X1 U4465 ( .A(n3901), .ZN(n3898) );
  OAI221_X1 U4466 ( .B1(n4784), .B2(n4785), .C1(n3780), .C2(n3885), .A(n4786), 
        .ZN(n3901) );
  NAND3_X1 U4467 ( .A1(\unit_fetch/pc_regout[3] ), .A2(
        \unit_fetch/pc_regout[4] ), .A3(n3857), .ZN(n4786) );
  NAND2_X1 U4468 ( .A1(n3857), .A2(n3771), .ZN(n3885) );
  INV_X1 U4469 ( .A(n3897), .ZN(n4785) );
  AOI211_X1 U4470 ( .C1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .C2(n3779), 
        .A(\unit_fetch/pc_regout[2] ), .B(n3826), .ZN(n4784) );
  NOR2_X1 U4471 ( .A1(n3779), .A2(\unit_fetch/unit_programCounter/ffi_1/n4 ), 
        .ZN(n3826) );
  MUX2_X1 U4472 ( .A(n4787), .B(n4788), .S(n3896), .Z(n3907) );
  INV_X1 U4473 ( .A(n3857), .ZN(n3896) );
  NOR2_X1 U4474 ( .A1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_1/n4 ), .ZN(n3857) );
  NAND2_X1 U4475 ( .A1(n3897), .A2(n3830), .ZN(n4788) );
  NAND2_X1 U4476 ( .A1(n3891), .A2(n3771), .ZN(n3830) );
  NOR2_X1 U4477 ( .A1(n3788), .A2(n3779), .ZN(n3891) );
  NOR2_X1 U4478 ( .A1(n3789), .A2(\unit_fetch/pc_regout[3] ), .ZN(n3897) );
  NAND2_X1 U4479 ( .A1(n3922), .A2(\unit_fetch/pc_regout[2] ), .ZN(n4787) );
  NOR2_X1 U4480 ( .A1(n3773), .A2(\unit_fetch/pc_regout[4] ), .ZN(n3922) );
endmodule

