package CONSTANTS is
   constant NumBit : integer := 8;	
end CONSTANTS;
