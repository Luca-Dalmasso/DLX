
module ffd_0 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n3, n1, n2, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n3) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_351 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_350 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_349 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_348 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_347 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_346 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_345 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_344 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_343 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_342 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_341 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_340 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_339 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_338 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_337 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_336 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_335 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_334 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_333 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_332 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_331 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_330 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_329 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_328 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N25 ( regIn, Clk, Reset, Enable, regOut );
  input [24:0] regIn;
  output [24:0] regOut;
  input Clk, Reset, Enable;


  ffd_0 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_351 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_350 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_349 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_348 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_347 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_346 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_345 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_344 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_343 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_342 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_341 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_340 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_339 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_338 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_337 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_336 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_335 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_334 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_333 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_332 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_331 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_330 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_329 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_328 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_327 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_326 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_325 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X8 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_324 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_323 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_322 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_321 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_320 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X2 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_319 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X2 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_318 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X2 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_317 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_316 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_315 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_314 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_313 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_312 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_311 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_310 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_309 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_308 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N20 ( regIn, Clk, Reset, Enable, regOut );
  input [19:0] regIn;
  output [19:0] regOut;
  input Clk, Reset, Enable;


  ffd_327 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_326 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_325 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_324 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_323 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_322 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_321 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_320 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_319 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_318 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_317 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_316 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_315 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_314 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_313 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_312 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_311 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_310 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_309 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_308 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_307 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_306 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_305 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_304 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_303 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_302 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module ffd_301 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_300 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_299 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N9 ( regIn, Clk, Reset, Enable, regOut );
  input [8:0] regIn;
  output [8:0] regOut;
  input Clk, Reset, Enable;


  ffd_307 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_306 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_305 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_304 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_303 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_302 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_301 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_300 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_299 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module dlx_cu ( Clk, Rst, IR_IN, IR_OUT_OPCODE, RD1_IN, RD1_OUT, CW_FETCH, 
        CW_DECODE, CW_EXE, CW_MEMWB, FETCH_STALL );
  input [31:0] IR_IN;
  input [5:0] IR_OUT_OPCODE;
  input [4:0] RD1_IN;
  input [4:0] RD1_OUT;
  output [2:0] CW_FETCH;
  output [4:0] CW_DECODE;
  output [10:0] CW_EXE;
  output [8:0] CW_MEMWB;
  input Clk, Rst;
  output FETCH_STALL;
  wire   IR_IN_10, IR_IN_9, IR_IN_8, IR_IN_7, IR_IN_6, IR_IN_5, IR_IN_4,
         IR_IN_3, IR_IN_2, IR_IN_1, IR_IN_0, cw_selected_24, cw_selected_23,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n155, n156;
  wire   [1:0] next_state;
  wire   [21:0] cw_selected;
  wire   [19:0] cw1delay;
  wire   [8:0] cw2delay;
  assign CW_FETCH[0] = 1'b1;
  assign CW_FETCH[1] = 1'b1;
  assign CW_FETCH[2] = 1'b1;
  assign IR_IN_10 = IR_IN[10];
  assign IR_IN_9 = IR_IN[9];
  assign IR_IN_8 = IR_IN[8];
  assign IR_IN_7 = IR_IN[7];
  assign IR_IN_6 = IR_IN[6];
  assign IR_IN_5 = IR_IN[5];
  assign IR_IN_4 = IR_IN[4];
  assign IR_IN_3 = IR_IN[3];
  assign IR_IN_2 = IR_IN[2];
  assign IR_IN_1 = IR_IN[1];
  assign IR_IN_0 = IR_IN[0];

  DFFR_X1 \current_state_reg[0]  ( .D(next_state[0]), .CK(Clk), .RN(n156), .Q(
        n153) );
  DFFR_X1 \current_state_reg[1]  ( .D(next_state[1]), .CK(Clk), .RN(n156), .Q(
        n152), .QN(n1) );
  regN_N25 uut_second_stage ( .regIn({cw_selected_24, cw_selected_23, 1'b1, 
        cw_selected[21:19], n155, cw_selected[17:6], cw_selected[6], 
        cw_selected[4:0]}), .Clk(Clk), .Reset(Rst), .Enable(1'b1), .regOut({
        CW_DECODE, cw1delay}) );
  regN_N20 uut_third_stage ( .regIn(cw1delay), .Clk(Clk), .Reset(Rst), 
        .Enable(1'b1), .regOut({CW_EXE, cw2delay}) );
  regN_N9 uut_fourth_stage ( .regIn(cw2delay), .Clk(Clk), .Reset(Rst), 
        .Enable(1'b1), .regOut(CW_MEMWB) );
  NOR4_X2 U3 ( .A1(RD1_IN[3]), .A2(RD1_IN[4]), .A3(RD1_IN[2]), .A4(n151), .ZN(
        n102) );
  NOR3_X1 U4 ( .A1(n2), .A2(n152), .A3(n153), .ZN(next_state[1]) );
  NOR4_X1 U5 ( .A1(n152), .A2(n153), .A3(n3), .A4(n4), .ZN(next_state[0]) );
  INV_X1 U6 ( .A(n5), .ZN(n155) );
  INV_X1 U7 ( .A(Rst), .ZN(n156) );
  NOR2_X1 U8 ( .A1(n6), .A2(n7), .ZN(cw_selected_24) );
  NAND2_X1 U9 ( .A1(n5), .A2(n8), .ZN(cw_selected_23) );
  NOR2_X1 U10 ( .A1(n9), .A2(n7), .ZN(cw_selected[9]) );
  NOR4_X1 U11 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n9) );
  OAI211_X1 U12 ( .C1(n14), .C2(n15), .A(n16), .B(n17), .ZN(n10) );
  NAND2_X1 U13 ( .A1(n18), .A2(n8), .ZN(cw_selected[6]) );
  INV_X1 U14 ( .A(cw_selected[7]), .ZN(n8) );
  NOR2_X1 U15 ( .A1(n7), .A2(n19), .ZN(cw_selected[7]) );
  NAND4_X1 U16 ( .A1(n18), .A2(n5), .A3(n20), .A4(n21), .ZN(cw_selected[4]) );
  AOI21_X1 U17 ( .B1(n22), .B2(n23), .A(cw_selected[21]), .ZN(n21) );
  INV_X1 U18 ( .A(cw_selected[3]), .ZN(n20) );
  INV_X1 U19 ( .A(cw_selected[8]), .ZN(n18) );
  NOR2_X1 U20 ( .A1(n7), .A2(n24), .ZN(cw_selected[8]) );
  AOI21_X1 U21 ( .B1(n25), .B2(n26), .A(n27), .ZN(cw_selected[3]) );
  NOR3_X1 U22 ( .A1(n28), .A2(n29), .A3(n30), .ZN(cw_selected[2]) );
  AOI21_X1 U23 ( .B1(n17), .B2(n31), .A(n7), .ZN(cw_selected[21]) );
  OAI22_X1 U24 ( .A1(n7), .A2(n32), .B1(n33), .B2(n28), .ZN(cw_selected[1]) );
  XNOR2_X1 U25 ( .A(IR_IN[26]), .B(IR_IN[28]), .ZN(n33) );
  INV_X1 U26 ( .A(n34), .ZN(cw_selected[19]) );
  AOI21_X1 U27 ( .B1(n35), .B2(cw_selected[20]), .A(cw_selected[16]), .ZN(n34)
         );
  OAI21_X1 U28 ( .B1(n36), .B2(n7), .A(n5), .ZN(cw_selected[17]) );
  NAND2_X1 U29 ( .A1(n22), .A2(n37), .ZN(n5) );
  OAI21_X1 U30 ( .B1(IR_IN[26]), .B2(n38), .A(n27), .ZN(cw_selected[15]) );
  NOR2_X1 U31 ( .A1(n39), .A2(n7), .ZN(cw_selected[14]) );
  NOR4_X1 U32 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n39) );
  INV_X1 U33 ( .A(n44), .ZN(n42) );
  NAND3_X1 U34 ( .A1(n45), .A2(n17), .A3(n46), .ZN(n41) );
  OAI211_X1 U35 ( .C1(n47), .C2(n25), .A(n48), .B(n49), .ZN(n40) );
  AND3_X1 U36 ( .A1(n50), .A2(n51), .A3(n15), .ZN(n49) );
  OAI211_X1 U37 ( .C1(n52), .C2(n7), .A(n38), .B(n27), .ZN(cw_selected[13]) );
  INV_X1 U38 ( .A(cw_selected[20]), .ZN(n27) );
  NOR2_X1 U39 ( .A1(n7), .A2(n53), .ZN(cw_selected[20]) );
  INV_X1 U40 ( .A(cw_selected[16]), .ZN(n38) );
  NOR3_X1 U41 ( .A1(n54), .A2(n55), .A3(n7), .ZN(cw_selected[16]) );
  NOR3_X1 U42 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n52) );
  OAI211_X1 U43 ( .C1(n59), .C2(n60), .A(n61), .B(n45), .ZN(n56) );
  NOR3_X1 U44 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n59) );
  NOR2_X1 U45 ( .A1(n65), .A2(n7), .ZN(cw_selected[12]) );
  AOI211_X1 U46 ( .C1(n64), .C2(n35), .A(n66), .B(n67), .ZN(n65) );
  OAI211_X1 U47 ( .C1(n68), .C2(n69), .A(n70), .B(n45), .ZN(n66) );
  NAND3_X1 U48 ( .A1(IR_IN_1), .A2(n71), .A3(n72), .ZN(n70) );
  INV_X1 U49 ( .A(n73), .ZN(n68) );
  NOR2_X1 U50 ( .A1(n74), .A2(n7), .ZN(cw_selected[11]) );
  NOR3_X1 U51 ( .A1(n75), .A2(n43), .A3(n76), .ZN(n74) );
  NOR4_X1 U52 ( .A1(IR_IN[27]), .A2(n77), .A3(n30), .A4(n25), .ZN(n76) );
  INV_X1 U53 ( .A(n78), .ZN(n43) );
  NOR2_X1 U54 ( .A1(n79), .A2(n7), .ZN(cw_selected[10]) );
  AOI211_X1 U55 ( .C1(n80), .C2(n81), .A(n82), .B(n83), .ZN(n79) );
  OAI33_X1 U56 ( .A1(n51), .A2(IR_IN_1), .A3(IR_IN_0), .B1(n84), .B2(n29), 
        .B3(n85), .ZN(n83) );
  INV_X1 U57 ( .A(n86), .ZN(n82) );
  AOI211_X1 U58 ( .C1(n87), .C2(n63), .A(n67), .B(n75), .ZN(n86) );
  OAI211_X1 U59 ( .C1(n71), .C2(n45), .A(n88), .B(n89), .ZN(n75) );
  AOI22_X1 U60 ( .A1(n80), .A2(n72), .B1(n90), .B2(n73), .ZN(n89) );
  NAND2_X1 U61 ( .A1(n91), .A2(n16), .ZN(n73) );
  INV_X1 U62 ( .A(n58), .ZN(n88) );
  OAI211_X1 U63 ( .C1(n26), .C2(n15), .A(n50), .B(n46), .ZN(n58) );
  OAI21_X1 U64 ( .B1(n92), .B2(n69), .A(n44), .ZN(n67) );
  INV_X1 U65 ( .A(n87), .ZN(n69) );
  AOI21_X1 U66 ( .B1(IR_IN[28]), .B2(n93), .A(n64), .ZN(n92) );
  INV_X1 U67 ( .A(n15), .ZN(n64) );
  NOR2_X1 U68 ( .A1(n71), .A2(n94), .ZN(n80) );
  OAI22_X1 U69 ( .A1(n7), .A2(n95), .B1(IR_IN[26]), .B2(n28), .ZN(
        cw_selected[0]) );
  NAND2_X1 U70 ( .A1(n96), .A2(n22), .ZN(n28) );
  INV_X1 U71 ( .A(n22), .ZN(n7) );
  NOR2_X1 U72 ( .A1(FETCH_STALL), .A2(Rst), .ZN(n22) );
  NOR2_X1 U73 ( .A1(n97), .A2(n153), .ZN(FETCH_STALL) );
  AND3_X1 U74 ( .A1(n2), .A2(n1), .A3(n4), .ZN(n97) );
  OAI21_X1 U75 ( .B1(n98), .B2(n99), .A(n100), .ZN(n4) );
  OR4_X1 U76 ( .A1(RD1_OUT[3]), .A2(RD1_OUT[4]), .A3(RD1_OUT[2]), .A4(n101), 
        .ZN(n100) );
  OR2_X1 U77 ( .A1(RD1_OUT[1]), .A2(RD1_OUT[0]), .ZN(n101) );
  OAI21_X1 U78 ( .B1(n98), .B2(n99), .A(n3), .ZN(n2) );
  INV_X1 U79 ( .A(n102), .ZN(n3) );
  AND4_X1 U80 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(n99) );
  NOR4_X1 U81 ( .A1(Rst), .A2(n6), .A3(n107), .A4(n108), .ZN(n106) );
  XNOR2_X1 U82 ( .A(n109), .B(IR_IN[21]), .ZN(n108) );
  XNOR2_X1 U83 ( .A(n110), .B(IR_IN[22]), .ZN(n107) );
  NOR2_X1 U84 ( .A1(n37), .A2(n111), .ZN(n6) );
  AOI21_X1 U85 ( .B1(n35), .B2(n112), .A(n36), .ZN(n111) );
  NOR3_X1 U86 ( .A1(n23), .A2(n57), .A3(n113), .ZN(n36) );
  OAI211_X1 U87 ( .C1(n54), .C2(n55), .A(n17), .B(n53), .ZN(n113) );
  NAND2_X1 U88 ( .A1(n114), .A2(n115), .ZN(n17) );
  OAI21_X1 U89 ( .B1(n116), .B2(n30), .A(n91), .ZN(n114) );
  NAND3_X1 U90 ( .A1(n85), .A2(n117), .A3(IR_IN[28]), .ZN(n54) );
  NAND3_X1 U91 ( .A1(n19), .A2(n31), .A3(n24), .ZN(n57) );
  NOR2_X1 U92 ( .A1(n96), .A2(n118), .ZN(n24) );
  AND4_X1 U93 ( .A1(n119), .A2(IR_IN[31]), .A3(n30), .A4(n77), .ZN(n118) );
  AND4_X1 U94 ( .A1(IR_IN[31]), .A2(n85), .A3(n77), .A4(n117), .ZN(n96) );
  OAI21_X1 U95 ( .B1(n62), .B2(n63), .A(n119), .ZN(n31) );
  OR4_X1 U96 ( .A1(n13), .A2(n120), .A3(n11), .A4(n121), .ZN(n23) );
  OAI211_X1 U97 ( .C1(n84), .C2(IR_IN[26]), .A(n15), .B(n50), .ZN(n121) );
  NAND4_X1 U98 ( .A1(n122), .A2(IR_IN[28]), .A3(IR_IN[27]), .A4(n123), .ZN(n50) );
  NAND3_X1 U99 ( .A1(IR_IN[28]), .A2(n85), .A3(n122), .ZN(n15) );
  INV_X1 U100 ( .A(n48), .ZN(n11) );
  AOI22_X1 U101 ( .A1(n87), .A2(n63), .B1(n115), .B2(n62), .ZN(n48) );
  INV_X1 U102 ( .A(n16), .ZN(n62) );
  INV_X1 U103 ( .A(n14), .ZN(n115) );
  NOR2_X1 U104 ( .A1(n90), .A2(n87), .ZN(n14) );
  INV_X1 U105 ( .A(n47), .ZN(n63) );
  NOR2_X1 U106 ( .A1(n117), .A2(IR_IN[26]), .ZN(n87) );
  NOR2_X1 U107 ( .A1(n47), .A2(n60), .ZN(n120) );
  OAI222_X1 U108 ( .A1(n85), .A2(n84), .B1(n47), .B2(n25), .C1(n60), .C2(n16), 
        .ZN(n13) );
  NAND2_X1 U109 ( .A1(n122), .A2(n124), .ZN(n16) );
  INV_X1 U110 ( .A(n90), .ZN(n25) );
  NOR2_X1 U111 ( .A1(n117), .A2(n29), .ZN(n90) );
  INV_X1 U112 ( .A(IR_IN[30]), .ZN(n117) );
  NAND3_X1 U113 ( .A1(n85), .A2(n30), .A3(n122), .ZN(n47) );
  NOR2_X1 U114 ( .A1(n77), .A2(IR_IN[31]), .ZN(n122) );
  INV_X1 U115 ( .A(IR_IN[29]), .ZN(n77) );
  NAND3_X1 U116 ( .A1(IR_IN[30]), .A2(n125), .A3(IR_IN[28]), .ZN(n84) );
  INV_X1 U117 ( .A(n53), .ZN(n112) );
  NAND2_X1 U118 ( .A1(n124), .A2(n125), .ZN(n53) );
  NAND2_X1 U119 ( .A1(n60), .A2(n26), .ZN(n35) );
  XOR2_X1 U120 ( .A(IR_IN[25]), .B(n126), .Z(n105) );
  XOR2_X1 U121 ( .A(IR_IN[24]), .B(n127), .Z(n104) );
  XOR2_X1 U122 ( .A(IR_IN[23]), .B(n128), .Z(n103) );
  AND4_X1 U123 ( .A1(n129), .A2(n130), .A3(n131), .A4(n132), .ZN(n98) );
  NOR3_X1 U124 ( .A1(n133), .A2(n134), .A3(n135), .ZN(n132) );
  XNOR2_X1 U125 ( .A(n128), .B(IR_IN[18]), .ZN(n135) );
  AOI21_X1 U126 ( .B1(n102), .B2(RD1_OUT[2]), .A(RD1_IN[2]), .ZN(n128) );
  XNOR2_X1 U127 ( .A(n127), .B(IR_IN[19]), .ZN(n134) );
  AOI21_X1 U128 ( .B1(n102), .B2(RD1_OUT[3]), .A(RD1_IN[3]), .ZN(n127) );
  XNOR2_X1 U129 ( .A(n126), .B(IR_IN[20]), .ZN(n133) );
  AOI21_X1 U130 ( .B1(n102), .B2(RD1_OUT[4]), .A(RD1_IN[4]), .ZN(n126) );
  AOI21_X1 U131 ( .B1(n136), .B2(n19), .A(Rst), .ZN(n131) );
  INV_X1 U132 ( .A(n137), .ZN(n19) );
  OAI211_X1 U133 ( .C1(n26), .C2(n91), .A(n32), .B(n95), .ZN(n137) );
  NAND3_X1 U134 ( .A1(n123), .A2(n30), .A3(n93), .ZN(n95) );
  NAND3_X1 U135 ( .A1(n93), .A2(n30), .A3(n119), .ZN(n32) );
  INV_X1 U136 ( .A(IR_IN[28]), .ZN(n30) );
  INV_X1 U137 ( .A(n116), .ZN(n93) );
  NAND3_X1 U138 ( .A1(IR_IN[29]), .A2(n85), .A3(IR_IN[31]), .ZN(n116) );
  NAND3_X1 U139 ( .A1(IR_IN[31]), .A2(IR_IN[29]), .A3(n124), .ZN(n91) );
  NOR2_X1 U140 ( .A1(n85), .A2(IR_IN[28]), .ZN(n124) );
  INV_X1 U141 ( .A(IR_IN[27]), .ZN(n85) );
  INV_X1 U142 ( .A(n119), .ZN(n26) );
  NOR2_X1 U143 ( .A1(n29), .A2(IR_IN[30]), .ZN(n119) );
  INV_X1 U144 ( .A(IR_IN[26]), .ZN(n29) );
  INV_X1 U145 ( .A(n37), .ZN(n136) );
  NAND4_X1 U146 ( .A1(n46), .A2(n45), .A3(n61), .A4(n138), .ZN(n37) );
  AOI21_X1 U147 ( .B1(n81), .B2(n71), .A(n12), .ZN(n138) );
  NAND4_X1 U148 ( .A1(n139), .A2(n51), .A3(n78), .A4(n44), .ZN(n12) );
  NAND3_X1 U149 ( .A1(n140), .A2(n71), .A3(IR_IN_3), .ZN(n44) );
  NAND3_X1 U150 ( .A1(IR_IN_3), .A2(n140), .A3(IR_IN_0), .ZN(n78) );
  INV_X1 U151 ( .A(n72), .ZN(n51) );
  NOR3_X1 U152 ( .A1(n141), .A2(n142), .A3(n143), .ZN(n72) );
  OAI21_X1 U153 ( .B1(n144), .B2(n81), .A(IR_IN_1), .ZN(n139) );
  NOR4_X1 U154 ( .A1(n145), .A2(n146), .A3(IR_IN_3), .A4(IR_IN_5), .ZN(n81) );
  INV_X1 U155 ( .A(n147), .ZN(n146) );
  INV_X1 U156 ( .A(n144), .ZN(n61) );
  NOR3_X1 U157 ( .A1(n142), .A2(IR_IN_3), .A3(n141), .ZN(n144) );
  NAND2_X1 U158 ( .A1(n140), .A2(n143), .ZN(n45) );
  NOR3_X1 U159 ( .A1(n145), .A2(IR_IN_1), .A3(n141), .ZN(n140) );
  NAND4_X1 U160 ( .A1(n71), .A2(n143), .A3(n142), .A4(n148), .ZN(n46) );
  NOR2_X1 U161 ( .A1(n141), .A2(n94), .ZN(n148) );
  INV_X1 U162 ( .A(IR_IN_1), .ZN(n94) );
  NAND3_X1 U163 ( .A1(n149), .A2(n147), .A3(IR_IN_5), .ZN(n141) );
  NOR4_X1 U164 ( .A1(IR_IN_6), .A2(IR_IN_4), .A3(IR_IN_10), .A4(n150), .ZN(
        n147) );
  OR3_X1 U165 ( .A1(IR_IN_9), .A2(IR_IN_8), .A3(IR_IN_7), .ZN(n150) );
  INV_X1 U166 ( .A(n145), .ZN(n142) );
  NAND2_X1 U167 ( .A1(IR_IN_2), .A2(n149), .ZN(n145) );
  NOR4_X1 U168 ( .A1(n60), .A2(n55), .A3(IR_IN[27]), .A4(IR_IN[28]), .ZN(n149)
         );
  INV_X1 U169 ( .A(n125), .ZN(n55) );
  NOR2_X1 U170 ( .A1(IR_IN[31]), .A2(IR_IN[29]), .ZN(n125) );
  INV_X1 U171 ( .A(n123), .ZN(n60) );
  NOR2_X1 U172 ( .A1(IR_IN[26]), .A2(IR_IN[30]), .ZN(n123) );
  INV_X1 U173 ( .A(IR_IN_3), .ZN(n143) );
  INV_X1 U174 ( .A(IR_IN_0), .ZN(n71) );
  XOR2_X1 U175 ( .A(IR_IN[17]), .B(n110), .Z(n130) );
  AOI21_X1 U176 ( .B1(n102), .B2(RD1_OUT[1]), .A(RD1_IN[1]), .ZN(n110) );
  XOR2_X1 U177 ( .A(IR_IN[16]), .B(n109), .Z(n129) );
  AOI21_X1 U178 ( .B1(n102), .B2(RD1_OUT[0]), .A(RD1_IN[0]), .ZN(n109) );
  OR2_X1 U179 ( .A1(RD1_IN[1]), .A2(RD1_IN[0]), .ZN(n151) );
endmodule


module ffd_298 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_297 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_296 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_295 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_294 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_293 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_292 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_291 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_290 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_289 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_288 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_287 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_286 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_285 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_284 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_283 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_282 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_281 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_280 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_279 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_278 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_277 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_276 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_275 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_274 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_273 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_272 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_271 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_270 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_269 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_268 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_267 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_0 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_298 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_297 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_296 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_295 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_294 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_293 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_292 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_291 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_290 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_289 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_288 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_287 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_286 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_285 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_284 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_283 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_282 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_281 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_280 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_279 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_278 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_277 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_276 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_275 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_274 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_273 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_272 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_271 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_270 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_269 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_268 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_267 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module IMemory_RAM_DEPTH40_I_SIZE8_NBIT32 ( Addr, Dout );
  input [31:0] Addr;
  output [31:0] Dout;
  wire   Dout_19, Dout_18, Dout_17, Dout_16, Dout_15, Dout_14, Dout_13,
         Dout_11, Dout_10, Dout_9, Dout_8, Dout_7, Dout_6, Dout_5, Dout_3,
         Dout_2, Dout_1, Dout_0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125;
  assign Dout[28] = Dout[30];
  assign Dout[20] = Dout[22];
  assign Dout[19] = Dout_19;
  assign Dout[18] = Dout_18;
  assign Dout[17] = Dout_17;
  assign Dout[16] = Dout_16;
  assign Dout[15] = Dout_15;
  assign Dout[12] = Dout_14;
  assign Dout[14] = Dout_14;
  assign Dout[13] = Dout_13;
  assign Dout[11] = Dout_11;
  assign Dout[10] = Dout_10;
  assign Dout[9] = Dout_9;
  assign Dout[8] = Dout_8;
  assign Dout[7] = Dout_7;
  assign Dout[4] = Dout_6;
  assign Dout[6] = Dout_6;
  assign Dout[5] = Dout_5;
  assign Dout[3] = Dout_3;
  assign Dout[2] = Dout_2;
  assign Dout[1] = Dout_1;
  assign Dout[0] = Dout_0;

  OAI211_X2 U1 ( .C1(n92), .C2(n93), .A(n94), .B(n95), .ZN(Dout[30]) );
  INV_X1 U2 ( .A(n1), .ZN(Dout[31]) );
  NAND3_X1 U3 ( .A1(n2), .A2(n3), .A3(n4), .ZN(Dout_9) );
  NAND2_X1 U4 ( .A1(n5), .A2(n4), .ZN(Dout_8) );
  AOI21_X1 U5 ( .B1(n6), .B2(n7), .A(n8), .ZN(n4) );
  NAND2_X1 U6 ( .A1(n9), .A2(n10), .ZN(Dout_6) );
  NAND2_X1 U7 ( .A1(n11), .A2(n10), .ZN(Dout_5) );
  INV_X1 U8 ( .A(Dout_7), .ZN(n10) );
  NAND2_X1 U9 ( .A1(n12), .A2(n13), .ZN(Dout_7) );
  INV_X1 U10 ( .A(n14), .ZN(n12) );
  NAND4_X1 U11 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Dout_3) );
  NOR2_X1 U12 ( .A1(n14), .A2(n19), .ZN(n18) );
  NAND3_X1 U13 ( .A1(n20), .A2(n9), .A3(n21), .ZN(Dout_2) );
  INV_X1 U14 ( .A(n22), .ZN(n21) );
  OAI211_X1 U15 ( .C1(n23), .C2(n24), .A(n25), .B(n26), .ZN(n22) );
  AOI221_X1 U16 ( .B1(n27), .B2(n28), .C1(n29), .C2(n30), .A(n31), .ZN(n9) );
  INV_X1 U17 ( .A(n32), .ZN(n28) );
  NAND4_X1 U18 ( .A1(n33), .A2(n34), .A3(n35), .A4(n26), .ZN(Dout_19) );
  INV_X1 U19 ( .A(n19), .ZN(n34) );
  NAND3_X1 U20 ( .A1(n36), .A2(n37), .A3(n38), .ZN(Dout_18) );
  AND3_X1 U21 ( .A1(n39), .A2(n25), .A3(n2), .ZN(n38) );
  OAI21_X1 U22 ( .B1(n24), .B2(n23), .A(n37), .ZN(Dout_17) );
  AND4_X1 U23 ( .A1(n33), .A2(n40), .A3(n17), .A4(n35), .ZN(n37) );
  NAND2_X1 U24 ( .A1(n41), .A2(n6), .ZN(n40) );
  NAND4_X1 U25 ( .A1(n42), .A2(n33), .A3(n17), .A4(n3), .ZN(Dout_16) );
  AOI211_X1 U26 ( .C1(n43), .C2(n44), .A(n31), .B(n45), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n46), .A2(n47), .ZN(Dout_14) );
  NAND2_X1 U28 ( .A1(n26), .A2(n47), .ZN(Dout_13) );
  INV_X1 U29 ( .A(Dout_15), .ZN(n47) );
  NAND4_X1 U30 ( .A1(n48), .A2(n16), .A3(n13), .A4(n49), .ZN(Dout_15) );
  NAND4_X1 U31 ( .A1(n17), .A2(n26), .A3(n48), .A4(n50), .ZN(Dout_11) );
  NOR2_X1 U32 ( .A1(n45), .A2(n19), .ZN(n50) );
  OAI21_X1 U33 ( .B1(n51), .B2(n52), .A(n11), .ZN(n19) );
  AOI22_X1 U34 ( .A1(n53), .A2(n54), .B1(n55), .B2(n56), .ZN(n51) );
  NAND3_X1 U35 ( .A1(n57), .A2(n58), .A3(n24), .ZN(n54) );
  NOR2_X1 U36 ( .A1(n7), .A2(n44), .ZN(n24) );
  NAND4_X1 U37 ( .A1(n46), .A2(n42), .A3(n59), .A4(n25), .ZN(Dout_10) );
  INV_X1 U38 ( .A(n8), .ZN(n59) );
  NAND4_X1 U39 ( .A1(n60), .A2(n48), .A3(n15), .A4(n26), .ZN(n8) );
  NAND2_X1 U40 ( .A1(n61), .A2(n53), .ZN(n26) );
  NAND2_X1 U41 ( .A1(n55), .A2(n61), .ZN(n15) );
  INV_X1 U42 ( .A(n45), .ZN(n60) );
  INV_X1 U43 ( .A(n62), .ZN(n42) );
  OAI211_X1 U44 ( .C1(n23), .C2(n63), .A(n35), .B(n2), .ZN(n62) );
  NAND2_X1 U45 ( .A1(n64), .A2(n6), .ZN(n2) );
  AOI22_X1 U46 ( .A1(n7), .A2(n30), .B1(n65), .B2(n61), .ZN(n46) );
  AND2_X1 U47 ( .A1(n41), .A2(n66), .ZN(n61) );
  NAND3_X1 U48 ( .A1(n5), .A2(n3), .A3(n20), .ZN(Dout_1) );
  AOI211_X1 U49 ( .C1(n67), .C2(n68), .A(n69), .B(n70), .ZN(n5) );
  INV_X1 U50 ( .A(n25), .ZN(n70) );
  NAND2_X1 U51 ( .A1(n71), .A2(n6), .ZN(n25) );
  AND3_X1 U52 ( .A1(n56), .A2(n66), .A3(n55), .ZN(n69) );
  OAI211_X1 U53 ( .C1(n23), .C2(n63), .A(n20), .B(n72), .ZN(Dout_0) );
  AOI211_X1 U54 ( .C1(n68), .C2(n73), .A(n74), .B(n75), .ZN(n72) );
  INV_X1 U55 ( .A(n17), .ZN(n75) );
  NAND2_X1 U56 ( .A1(n76), .A2(n55), .ZN(n17) );
  INV_X1 U57 ( .A(n3), .ZN(n74) );
  NAND2_X1 U58 ( .A1(n29), .A2(n6), .ZN(n3) );
  INV_X1 U59 ( .A(n23), .ZN(n6) );
  AND4_X1 U60 ( .A1(n77), .A2(n78), .A3(n79), .A4(n80), .ZN(n68) );
  NOR2_X1 U61 ( .A1(n81), .A2(n82), .ZN(n80) );
  NAND4_X1 U62 ( .A1(Addr[14]), .A2(Addr[13]), .A3(Addr[12]), .A4(Addr[11]), 
        .ZN(n82) );
  NAND4_X1 U63 ( .A1(Addr[10]), .A2(Addr[3]), .A3(Addr[2]), .A4(Addr[4]), .ZN(
        n81) );
  NOR4_X1 U64 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(n79) );
  NAND4_X1 U65 ( .A1(Addr[18]), .A2(Addr[17]), .A3(Addr[16]), .A4(Addr[15]), 
        .ZN(n83) );
  AND4_X1 U66 ( .A1(n87), .A2(Addr[28]), .A3(Addr[26]), .A4(Addr[27]), .ZN(n78) );
  AND4_X1 U67 ( .A1(Addr[25]), .A2(Addr[24]), .A3(Addr[23]), .A4(Addr[22]), 
        .ZN(n87) );
  AND4_X1 U68 ( .A1(n88), .A2(Addr[9]), .A3(Addr[7]), .A4(Addr[8]), .ZN(n77)
         );
  AND4_X1 U69 ( .A1(Addr[6]), .A2(Addr[5]), .A3(Addr[30]), .A4(Addr[29]), .ZN(
        n88) );
  AND3_X1 U70 ( .A1(n11), .A2(n16), .A3(n89), .ZN(n20) );
  AOI21_X1 U71 ( .B1(n27), .B2(n55), .A(n14), .ZN(n89) );
  NAND3_X1 U72 ( .A1(n35), .A2(n90), .A3(n48), .ZN(n14) );
  AOI21_X1 U73 ( .B1(n43), .B2(n44), .A(n91), .ZN(n48) );
  INV_X1 U74 ( .A(n39), .ZN(n91) );
  NAND3_X1 U75 ( .A1(n53), .A2(n66), .A3(n56), .ZN(n39) );
  NAND2_X1 U76 ( .A1(n27), .A2(n53), .ZN(n11) );
  AND2_X1 U77 ( .A1(n64), .A2(n66), .ZN(n27) );
  OAI21_X1 U78 ( .B1(n55), .B2(n53), .A(n66), .ZN(n23) );
  NOR3_X1 U79 ( .A1(Addr[4]), .A2(Addr[5]), .A3(Addr[3]), .ZN(n55) );
  NAND3_X1 U80 ( .A1(Addr[3]), .A2(Addr[4]), .A3(n67), .ZN(n94) );
  AOI211_X1 U81 ( .C1(Addr[0]), .C2(n96), .A(Addr[2]), .B(n73), .ZN(n92) );
  NAND2_X1 U82 ( .A1(n1), .A2(n97), .ZN(Dout[29]) );
  NAND3_X1 U83 ( .A1(Addr[3]), .A2(n98), .A3(n56), .ZN(n97) );
  NOR2_X1 U84 ( .A1(n99), .A2(n100), .ZN(n56) );
  OAI21_X1 U85 ( .B1(n101), .B2(n102), .A(n103), .ZN(n1) );
  AOI21_X1 U86 ( .B1(n104), .B2(n96), .A(n67), .ZN(n102) );
  OAI221_X1 U87 ( .B1(n105), .B2(n93), .C1(Addr[4]), .C2(n106), .A(n107), .ZN(
        Dout[27]) );
  NAND3_X1 U88 ( .A1(n108), .A2(n95), .A3(n109), .ZN(Dout[26]) );
  MUX2_X1 U89 ( .A(n110), .B(n99), .S(Addr[4]), .Z(n109) );
  NAND2_X1 U90 ( .A1(Addr[2]), .A2(n111), .ZN(n110) );
  NAND2_X1 U91 ( .A1(Addr[5]), .A2(n71), .ZN(n95) );
  OAI21_X1 U92 ( .B1(n100), .B2(n96), .A(n103), .ZN(n108) );
  OAI221_X1 U93 ( .B1(n96), .B2(n112), .C1(n93), .C2(n113), .A(n107), .ZN(
        Dout[25]) );
  NAND3_X1 U94 ( .A1(Addr[0]), .A2(n100), .A3(n103), .ZN(n107) );
  INV_X1 U95 ( .A(n93), .ZN(n103) );
  NAND2_X1 U96 ( .A1(n114), .A2(n111), .ZN(n112) );
  OAI21_X1 U97 ( .B1(n105), .B2(n93), .A(n115), .ZN(Dout[24]) );
  NAND3_X1 U98 ( .A1(n114), .A2(n111), .A3(Addr[0]), .ZN(n115) );
  OAI21_X1 U99 ( .B1(Addr[3]), .B2(Addr[2]), .A(Addr[4]), .ZN(n114) );
  AOI21_X1 U100 ( .B1(n100), .B2(Addr[1]), .A(n101), .ZN(n105) );
  INV_X1 U101 ( .A(n113), .ZN(n101) );
  INV_X1 U102 ( .A(n116), .ZN(Dout[23]) );
  NAND2_X1 U103 ( .A1(n36), .A2(n116), .ZN(Dout[22]) );
  AOI22_X1 U104 ( .A1(n65), .A2(n76), .B1(n44), .B2(n30), .ZN(n36) );
  AOI21_X1 U105 ( .B1(n32), .B2(n117), .A(n52), .ZN(n30) );
  NAND3_X1 U106 ( .A1(Addr[5]), .A2(n98), .A3(n106), .ZN(n117) );
  INV_X1 U107 ( .A(Addr[4]), .ZN(n98) );
  INV_X1 U108 ( .A(n63), .ZN(n44) );
  NAND2_X1 U109 ( .A1(n73), .A2(n100), .ZN(n63) );
  OAI21_X1 U110 ( .B1(Addr[5]), .B2(n93), .A(n32), .ZN(n65) );
  NAND3_X1 U111 ( .A1(Addr[4]), .A2(n111), .A3(Addr[3]), .ZN(n32) );
  INV_X1 U112 ( .A(Addr[5]), .ZN(n111) );
  NAND2_X1 U113 ( .A1(n35), .A2(n116), .ZN(Dout[21]) );
  AOI211_X1 U114 ( .C1(n43), .C2(n41), .A(n31), .B(n45), .ZN(n116) );
  NAND3_X1 U115 ( .A1(n16), .A2(n13), .A3(n90), .ZN(n45) );
  NAND2_X1 U116 ( .A1(n7), .A2(n43), .ZN(n90) );
  NOR3_X1 U117 ( .A1(Addr[1]), .A2(Addr[2]), .A3(n104), .ZN(n7) );
  NAND2_X1 U118 ( .A1(n71), .A2(n43), .ZN(n13) );
  INV_X1 U119 ( .A(n58), .ZN(n71) );
  NAND2_X1 U120 ( .A1(n67), .A2(n100), .ZN(n58) );
  INV_X1 U121 ( .A(n99), .ZN(n67) );
  NAND2_X1 U122 ( .A1(Addr[1]), .A2(Addr[0]), .ZN(n99) );
  NAND2_X1 U123 ( .A1(n43), .A2(n29), .ZN(n16) );
  INV_X1 U124 ( .A(n57), .ZN(n29) );
  NAND3_X1 U125 ( .A1(n96), .A2(n100), .A3(n104), .ZN(n57) );
  INV_X1 U126 ( .A(Addr[2]), .ZN(n100) );
  INV_X1 U127 ( .A(n49), .ZN(n31) );
  NAND2_X1 U128 ( .A1(n43), .A2(n64), .ZN(n49) );
  NOR2_X1 U129 ( .A1(n113), .A2(Addr[0]), .ZN(n64) );
  NOR2_X1 U130 ( .A1(n113), .A2(n104), .ZN(n41) );
  INV_X1 U131 ( .A(Addr[0]), .ZN(n104) );
  NAND2_X1 U132 ( .A1(Addr[2]), .A2(n96), .ZN(n113) );
  NOR3_X1 U133 ( .A1(n93), .A2(Addr[5]), .A3(n52), .ZN(n43) );
  NAND2_X1 U134 ( .A1(Addr[4]), .A2(n106), .ZN(n93) );
  NAND2_X1 U135 ( .A1(n76), .A2(n53), .ZN(n35) );
  NOR3_X1 U136 ( .A1(Addr[4]), .A2(Addr[5]), .A3(n106), .ZN(n53) );
  INV_X1 U137 ( .A(Addr[3]), .ZN(n106) );
  AND3_X1 U138 ( .A1(n66), .A2(Addr[2]), .A3(n73), .ZN(n76) );
  NOR2_X1 U139 ( .A1(n96), .A2(Addr[0]), .ZN(n73) );
  INV_X1 U140 ( .A(Addr[1]), .ZN(n96) );
  INV_X1 U141 ( .A(n52), .ZN(n66) );
  NAND4_X1 U142 ( .A1(n118), .A2(n119), .A3(n120), .A4(n121), .ZN(n52) );
  NOR4_X1 U143 ( .A1(n122), .A2(Addr[28]), .A3(Addr[30]), .A4(Addr[29]), .ZN(
        n121) );
  OR4_X1 U144 ( .A1(Addr[6]), .A2(Addr[7]), .A3(Addr[8]), .A4(Addr[9]), .ZN(
        n122) );
  NOR4_X1 U145 ( .A1(n123), .A2(Addr[22]), .A3(Addr[24]), .A4(Addr[23]), .ZN(
        n120) );
  OR3_X1 U146 ( .A1(Addr[26]), .A2(Addr[27]), .A3(Addr[25]), .ZN(n123) );
  NOR4_X1 U147 ( .A1(n124), .A2(Addr[16]), .A3(Addr[18]), .A4(Addr[17]), .ZN(
        n119) );
  NAND3_X1 U148 ( .A1(n86), .A2(n84), .A3(n85), .ZN(n124) );
  INV_X1 U149 ( .A(Addr[19]), .ZN(n85) );
  INV_X1 U150 ( .A(Addr[21]), .ZN(n84) );
  INV_X1 U151 ( .A(Addr[20]), .ZN(n86) );
  NOR4_X1 U152 ( .A1(n125), .A2(Addr[10]), .A3(Addr[12]), .A4(Addr[11]), .ZN(
        n118) );
  OR3_X1 U153 ( .A1(Addr[14]), .A2(Addr[15]), .A3(Addr[13]), .ZN(n125) );
endmodule


module IRreg_N32 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  DFF_X1 \regOut_reg[31]  ( .D(n71), .CK(Clk), .Q(regOut[31]), .QN(n66) );
  DFF_X1 \regOut_reg[30]  ( .D(n70), .CK(Clk), .Q(regOut[30]) );
  DFF_X1 \regOut_reg[29]  ( .D(n72), .CK(Clk), .Q(regOut[29]), .QN(n65) );
  DFF_X1 \regOut_reg[28]  ( .D(n69), .CK(Clk), .Q(regOut[28]) );
  DFF_X1 \regOut_reg[27]  ( .D(n73), .CK(Clk), .Q(regOut[27]), .QN(n64) );
  DFF_X1 \regOut_reg[26]  ( .D(n68), .CK(Clk), .Q(regOut[26]) );
  DFF_X1 \regOut_reg[25]  ( .D(n74), .CK(Clk), .Q(regOut[25]), .QN(n63) );
  DFF_X1 \regOut_reg[24]  ( .D(n75), .CK(Clk), .Q(regOut[24]), .QN(n62) );
  DFF_X1 \regOut_reg[23]  ( .D(n67), .CK(Clk), .Q(regOut[23]), .QN(n61) );
  DFF_X1 \regOut_reg[21]  ( .D(n77), .CK(Clk), .QN(n59) );
  DFF_X1 \regOut_reg[20]  ( .D(n78), .CK(Clk), .Q(regOut[20]), .QN(n58) );
  DFF_X1 \regOut_reg[19]  ( .D(n79), .CK(Clk), .Q(regOut[19]), .QN(n57) );
  DFF_X1 \regOut_reg[18]  ( .D(n80), .CK(Clk), .Q(regOut[18]), .QN(n56) );
  DFF_X1 \regOut_reg[16]  ( .D(n82), .CK(Clk), .QN(n54) );
  DFF_X1 \regOut_reg[15]  ( .D(n83), .CK(Clk), .Q(regOut[15]), .QN(n53) );
  DFF_X1 \regOut_reg[14]  ( .D(n84), .CK(Clk), .Q(regOut[14]), .QN(n52) );
  DFF_X1 \regOut_reg[13]  ( .D(n85), .CK(Clk), .Q(regOut[13]), .QN(n51) );
  DFF_X1 \regOut_reg[12]  ( .D(n86), .CK(Clk), .Q(regOut[12]), .QN(n50) );
  DFF_X1 \regOut_reg[11]  ( .D(n87), .CK(Clk), .Q(regOut[11]), .QN(n49) );
  DFF_X1 \regOut_reg[10]  ( .D(n88), .CK(Clk), .Q(regOut[10]), .QN(n48) );
  DFF_X1 \regOut_reg[9]  ( .D(n89), .CK(Clk), .Q(regOut[9]), .QN(n47) );
  DFF_X1 \regOut_reg[8]  ( .D(n90), .CK(Clk), .Q(regOut[8]), .QN(n46) );
  DFF_X1 \regOut_reg[7]  ( .D(n91), .CK(Clk), .Q(regOut[7]), .QN(n45) );
  DFF_X1 \regOut_reg[6]  ( .D(n92), .CK(Clk), .Q(regOut[6]), .QN(n44) );
  DFF_X1 \regOut_reg[5]  ( .D(n93), .CK(Clk), .Q(regOut[5]), .QN(n43) );
  DFF_X1 \regOut_reg[4]  ( .D(n94), .CK(Clk), .Q(regOut[4]), .QN(n42) );
  DFF_X1 \regOut_reg[3]  ( .D(n95), .CK(Clk), .Q(regOut[3]), .QN(n41) );
  DFF_X1 \regOut_reg[2]  ( .D(n96), .CK(Clk), .Q(regOut[2]), .QN(n40) );
  DFF_X1 \regOut_reg[1]  ( .D(n97), .CK(Clk), .Q(regOut[1]), .QN(n39) );
  DFF_X1 \regOut_reg[0]  ( .D(n98), .CK(Clk), .Q(regOut[0]), .QN(n38) );
  DFF_X2 \regOut_reg[17]  ( .D(n81), .CK(Clk), .Q(regOut[17]), .QN(n55) );
  DFF_X2 \regOut_reg[22]  ( .D(n76), .CK(Clk), .Q(regOut[22]), .QN(n60) );
  INV_X2 U3 ( .A(n37), .ZN(n3) );
  OR2_X2 U4 ( .A1(n37), .A2(Reset), .ZN(n4) );
  INV_X4 U5 ( .A(n59), .ZN(regOut[21]) );
  INV_X4 U6 ( .A(n54), .ZN(regOut[16]) );
  OAI22_X1 U7 ( .A1(n3), .A2(n61), .B1(n4), .B2(n5), .ZN(n67) );
  INV_X1 U8 ( .A(regIn[23]), .ZN(n5) );
  OR2_X1 U9 ( .A1(Reset), .A2(n6), .ZN(n68) );
  MUX2_X1 U10 ( .A(regOut[26]), .B(regIn[26]), .S(n3), .Z(n6) );
  OR2_X1 U11 ( .A1(Reset), .A2(n7), .ZN(n69) );
  MUX2_X1 U12 ( .A(regOut[28]), .B(regIn[28]), .S(n3), .Z(n7) );
  OR2_X1 U13 ( .A1(Reset), .A2(n8), .ZN(n70) );
  MUX2_X1 U14 ( .A(regOut[30]), .B(regIn[30]), .S(n3), .Z(n8) );
  OAI22_X1 U15 ( .A1(n3), .A2(n66), .B1(n4), .B2(n9), .ZN(n71) );
  INV_X1 U16 ( .A(regIn[31]), .ZN(n9) );
  OAI22_X1 U17 ( .A1(n3), .A2(n65), .B1(n4), .B2(n10), .ZN(n72) );
  INV_X1 U18 ( .A(regIn[29]), .ZN(n10) );
  OAI22_X1 U19 ( .A1(n3), .A2(n64), .B1(n4), .B2(n11), .ZN(n73) );
  INV_X1 U20 ( .A(regIn[27]), .ZN(n11) );
  OAI22_X1 U21 ( .A1(n3), .A2(n63), .B1(n4), .B2(n12), .ZN(n74) );
  INV_X1 U22 ( .A(regIn[25]), .ZN(n12) );
  OAI22_X1 U23 ( .A1(n3), .A2(n62), .B1(n4), .B2(n13), .ZN(n75) );
  INV_X1 U24 ( .A(regIn[24]), .ZN(n13) );
  OAI22_X1 U25 ( .A1(n3), .A2(n60), .B1(n4), .B2(n14), .ZN(n76) );
  INV_X1 U26 ( .A(regIn[22]), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n3), .A2(n59), .B1(n4), .B2(n15), .ZN(n77) );
  INV_X1 U28 ( .A(regIn[21]), .ZN(n15) );
  OAI22_X1 U29 ( .A1(n3), .A2(n58), .B1(n4), .B2(n16), .ZN(n78) );
  INV_X1 U30 ( .A(regIn[20]), .ZN(n16) );
  OAI22_X1 U31 ( .A1(n3), .A2(n57), .B1(n4), .B2(n17), .ZN(n79) );
  INV_X1 U32 ( .A(regIn[19]), .ZN(n17) );
  OAI22_X1 U33 ( .A1(n3), .A2(n56), .B1(n4), .B2(n18), .ZN(n80) );
  INV_X1 U34 ( .A(regIn[18]), .ZN(n18) );
  OAI22_X1 U35 ( .A1(n3), .A2(n55), .B1(n4), .B2(n19), .ZN(n81) );
  INV_X1 U36 ( .A(regIn[17]), .ZN(n19) );
  OAI22_X1 U37 ( .A1(n3), .A2(n54), .B1(n4), .B2(n20), .ZN(n82) );
  INV_X1 U38 ( .A(regIn[16]), .ZN(n20) );
  OAI22_X1 U39 ( .A1(n3), .A2(n53), .B1(n4), .B2(n21), .ZN(n83) );
  INV_X1 U40 ( .A(regIn[15]), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n3), .A2(n52), .B1(n4), .B2(n22), .ZN(n84) );
  INV_X1 U42 ( .A(regIn[14]), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n3), .A2(n51), .B1(n4), .B2(n23), .ZN(n85) );
  INV_X1 U44 ( .A(regIn[13]), .ZN(n23) );
  OAI22_X1 U45 ( .A1(n3), .A2(n50), .B1(n4), .B2(n24), .ZN(n86) );
  INV_X1 U46 ( .A(regIn[12]), .ZN(n24) );
  OAI22_X1 U47 ( .A1(n3), .A2(n49), .B1(n4), .B2(n25), .ZN(n87) );
  INV_X1 U48 ( .A(regIn[11]), .ZN(n25) );
  OAI22_X1 U49 ( .A1(n3), .A2(n48), .B1(n4), .B2(n26), .ZN(n88) );
  INV_X1 U50 ( .A(regIn[10]), .ZN(n26) );
  OAI22_X1 U51 ( .A1(n3), .A2(n47), .B1(n4), .B2(n27), .ZN(n89) );
  INV_X1 U52 ( .A(regIn[9]), .ZN(n27) );
  OAI22_X1 U53 ( .A1(n3), .A2(n46), .B1(n4), .B2(n28), .ZN(n90) );
  INV_X1 U54 ( .A(regIn[8]), .ZN(n28) );
  OAI22_X1 U55 ( .A1(n3), .A2(n45), .B1(n4), .B2(n29), .ZN(n91) );
  INV_X1 U56 ( .A(regIn[7]), .ZN(n29) );
  OAI22_X1 U57 ( .A1(n3), .A2(n44), .B1(n4), .B2(n30), .ZN(n92) );
  INV_X1 U58 ( .A(regIn[6]), .ZN(n30) );
  OAI22_X1 U59 ( .A1(n3), .A2(n43), .B1(n4), .B2(n31), .ZN(n93) );
  INV_X1 U60 ( .A(regIn[5]), .ZN(n31) );
  OAI22_X1 U61 ( .A1(n3), .A2(n42), .B1(n4), .B2(n32), .ZN(n94) );
  INV_X1 U62 ( .A(regIn[4]), .ZN(n32) );
  OAI22_X1 U63 ( .A1(n3), .A2(n41), .B1(n4), .B2(n33), .ZN(n95) );
  INV_X1 U64 ( .A(regIn[3]), .ZN(n33) );
  OAI22_X1 U65 ( .A1(n3), .A2(n40), .B1(n4), .B2(n34), .ZN(n96) );
  INV_X1 U66 ( .A(regIn[2]), .ZN(n34) );
  OAI22_X1 U67 ( .A1(n3), .A2(n39), .B1(n4), .B2(n35), .ZN(n97) );
  INV_X1 U68 ( .A(regIn[1]), .ZN(n35) );
  OAI22_X1 U69 ( .A1(n3), .A2(n38), .B1(n4), .B2(n36), .ZN(n98) );
  INV_X1 U70 ( .A(regIn[0]), .ZN(n36) );
  NOR2_X1 U71 ( .A1(Reset), .A2(Enable), .ZN(n37) );
endmodule


module Adder_N32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U1 ( .A(A[4]), .B(n32), .Z(SUM[4]) );
  XOR2_X1 U2 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U3 ( .A(A[5]), .B(n30), .Z(SUM[5]) );
  XNOR2_X1 U4 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  XOR2_X1 U5 ( .A(A[30]), .B(n42), .Z(SUM[30]) );
  XOR2_X1 U6 ( .A(A[16]), .B(n40), .Z(SUM[16]) );
  XOR2_X1 U7 ( .A(A[12]), .B(n34), .Z(SUM[12]) );
  XOR2_X1 U8 ( .A(A[11]), .B(n36), .Z(SUM[11]) );
  XOR2_X1 U9 ( .A(A[10]), .B(n51), .Z(SUM[10]) );
  XOR2_X1 U10 ( .A(A[17]), .B(n33), .Z(SUM[17]) );
  XOR2_X1 U11 ( .A(A[18]), .B(n37), .Z(SUM[18]) );
  XOR2_X1 U12 ( .A(A[6]), .B(n31), .Z(SUM[6]) );
  XOR2_X1 U13 ( .A(A[7]), .B(n52), .Z(SUM[7]) );
  XOR2_X1 U14 ( .A(A[8]), .B(n49), .Z(SUM[8]) );
  XOR2_X1 U15 ( .A(A[9]), .B(n50), .Z(SUM[9]) );
  XOR2_X1 U16 ( .A(A[13]), .B(n35), .Z(SUM[13]) );
  XOR2_X1 U17 ( .A(A[14]), .B(n45), .Z(SUM[14]) );
  XOR2_X1 U18 ( .A(A[15]), .B(n46), .Z(SUM[15]) );
  XOR2_X1 U19 ( .A(A[22]), .B(n56), .Z(SUM[22]) );
  XOR2_X1 U20 ( .A(A[23]), .B(n39), .Z(SUM[23]) );
  XOR2_X1 U21 ( .A(A[24]), .B(n43), .Z(SUM[24]) );
  XOR2_X1 U22 ( .A(A[25]), .B(n44), .Z(SUM[25]) );
  XOR2_X1 U23 ( .A(A[26]), .B(n53), .Z(SUM[26]) );
  XOR2_X1 U24 ( .A(A[27]), .B(n47), .Z(SUM[27]) );
  XOR2_X1 U25 ( .A(A[28]), .B(n48), .Z(SUM[28]) );
  XOR2_X1 U26 ( .A(A[29]), .B(n41), .Z(SUM[29]) );
  XOR2_X1 U27 ( .A(A[19]), .B(n38), .Z(SUM[19]) );
  XOR2_X1 U28 ( .A(A[20]), .B(n54), .Z(SUM[20]) );
  XOR2_X1 U29 ( .A(A[21]), .B(n55), .Z(SUM[21]) );
  INV_X1 U30 ( .A(A[2]), .ZN(SUM[2]) );
  NAND2_X1 U31 ( .A1(A[30]), .A2(n42), .ZN(n57) );
  AND2_X1 U32 ( .A1(A[4]), .A2(n32), .ZN(n30) );
  AND2_X1 U33 ( .A1(A[5]), .A2(n30), .ZN(n31) );
  AND2_X1 U34 ( .A1(A[3]), .A2(A[2]), .ZN(n32) );
  AND2_X1 U35 ( .A1(A[16]), .A2(n40), .ZN(n33) );
  AND2_X1 U36 ( .A1(A[11]), .A2(n36), .ZN(n34) );
  AND2_X1 U37 ( .A1(A[12]), .A2(n34), .ZN(n35) );
  AND2_X1 U38 ( .A1(A[10]), .A2(n51), .ZN(n36) );
  AND2_X1 U39 ( .A1(A[17]), .A2(n33), .ZN(n37) );
  AND2_X1 U40 ( .A1(A[18]), .A2(n37), .ZN(n38) );
  AND2_X1 U41 ( .A1(A[22]), .A2(n56), .ZN(n39) );
  AND2_X1 U42 ( .A1(A[15]), .A2(n46), .ZN(n40) );
  AND2_X1 U43 ( .A1(A[28]), .A2(n48), .ZN(n41) );
  AND2_X1 U44 ( .A1(A[29]), .A2(n41), .ZN(n42) );
  AND2_X1 U45 ( .A1(A[23]), .A2(n39), .ZN(n43) );
  AND2_X1 U46 ( .A1(A[24]), .A2(n43), .ZN(n44) );
  AND2_X1 U47 ( .A1(A[13]), .A2(n35), .ZN(n45) );
  AND2_X1 U48 ( .A1(A[14]), .A2(n45), .ZN(n46) );
  AND2_X1 U49 ( .A1(A[26]), .A2(n53), .ZN(n47) );
  AND2_X1 U50 ( .A1(A[27]), .A2(n47), .ZN(n48) );
  AND2_X1 U51 ( .A1(A[7]), .A2(n52), .ZN(n49) );
  AND2_X1 U52 ( .A1(A[8]), .A2(n49), .ZN(n50) );
  AND2_X1 U53 ( .A1(A[9]), .A2(n50), .ZN(n51) );
  AND2_X1 U54 ( .A1(A[6]), .A2(n31), .ZN(n52) );
  AND2_X1 U55 ( .A1(A[25]), .A2(n44), .ZN(n53) );
  AND2_X1 U56 ( .A1(A[19]), .A2(n38), .ZN(n54) );
  AND2_X1 U57 ( .A1(A[20]), .A2(n54), .ZN(n55) );
  AND2_X1 U58 ( .A1(A[21]), .A2(n55), .ZN(n56) );
endmodule


module Adder_N32 ( PC, NPC );
  input [31:0] PC;
  output [31:0] NPC;


  Adder_N32_DW01_add_0 add_19 ( .A(PC), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM(NPC) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_0 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_191 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_190 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_189 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_188 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_187 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_186 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_185 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_184 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_183 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_182 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_181 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_180 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_179 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_178 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_177 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_176 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_175 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_174 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_173 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_172 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_171 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_170 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_169 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_168 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_167 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_166 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_165 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_164 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_163 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_162 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_161 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module ffd_266 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_265 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_264 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_263 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_262 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_261 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_260 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_259 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_258 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_257 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_256 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_255 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_254 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_253 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_252 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_251 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_250 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_249 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_248 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_247 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_246 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_245 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_244 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_243 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_242 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_241 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_240 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_239 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_238 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_237 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_236 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_235 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_8 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_266 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_265 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_264 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_263 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_262 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_261 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_260 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_259 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_258 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_257 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_256 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_255 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_254 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_253 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_252 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_251 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_250 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_249 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_248 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_247 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_246 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_245 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_244 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_243 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_242 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_241 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_240 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_239 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_238 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_237 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_236 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_235 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module FU_N32 ( IR_En, PC_En, NPC_En, Clk, RST, COND_REGOUT, FLUSH, ALU_OUT, 
        IR_IN, IR_OUT, NPC_OUT );
  input [31:0] ALU_OUT;
  output [31:0] IR_IN;
  output [31:0] IR_OUT;
  output [31:0] NPC_OUT;
  input IR_En, PC_En, NPC_En, Clk, RST, COND_REGOUT, FLUSH;
  wire   reset_IR;
  wire   [31:0] npc_regin;
  wire   [31:0] pc_regout;
  wire   [31:0] adder_out;

  regN_N32_0 unit_programCounter ( .regIn(npc_regin), .Clk(Clk), .Reset(RST), 
        .Enable(PC_En), .regOut(pc_regout) );
  IMemory_RAM_DEPTH40_I_SIZE8_NBIT32 unit_instructionMemory ( .Addr(pc_regout), 
        .Dout(IR_IN) );
  IRreg_N32 unit_instructionRegister ( .regIn(IR_IN), .Clk(Clk), .Reset(
        reset_IR), .Enable(IR_En), .regOut(IR_OUT) );
  Adder_N32 unit_adder ( .PC(pc_regout), .NPC(adder_out) );
  MUX21_GENERIC_NBIT32_0 unit_mpx ( .A(ALU_OUT), .B(adder_out), .SEL(
        COND_REGOUT), .Y(npc_regin) );
  regN_N32_8 unit_npcregister ( .regIn(npc_regin), .Clk(Clk), .Reset(RST), 
        .Enable(NPC_En), .regOut(NPC_OUT) );
  OR2_X1 U1 ( .A1(FLUSH), .A2(RST), .ZN(reset_IR) );
endmodule


module register_file_WORD_SIZE32_ADDR_SIZE5 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n2163), .CK(CLK), .Q(\REGISTERS[0][31] )
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n2162), .CK(CLK), .Q(\REGISTERS[0][30] )
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n2161), .CK(CLK), .Q(\REGISTERS[0][29] )
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n2160), .CK(CLK), .Q(\REGISTERS[0][28] )
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n2159), .CK(CLK), .Q(\REGISTERS[0][27] )
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n2158), .CK(CLK), .Q(\REGISTERS[0][26] )
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n2157), .CK(CLK), .Q(\REGISTERS[0][25] )
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n2156), .CK(CLK), .Q(\REGISTERS[0][24] )
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n2155), .CK(CLK), .Q(\REGISTERS[0][23] )
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n2154), .CK(CLK), .Q(\REGISTERS[0][22] )
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n2153), .CK(CLK), .Q(\REGISTERS[0][21] )
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n2152), .CK(CLK), .Q(\REGISTERS[0][20] )
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n2151), .CK(CLK), .Q(\REGISTERS[0][19] )
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n2150), .CK(CLK), .Q(\REGISTERS[0][18] )
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n2149), .CK(CLK), .Q(\REGISTERS[0][17] )
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n2148), .CK(CLK), .Q(\REGISTERS[0][16] )
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n2147), .CK(CLK), .Q(\REGISTERS[0][15] )
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n2146), .CK(CLK), .Q(\REGISTERS[0][14] )
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n2145), .CK(CLK), .Q(\REGISTERS[0][13] )
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n2144), .CK(CLK), .Q(\REGISTERS[0][12] )
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n2143), .CK(CLK), .Q(\REGISTERS[0][11] )
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n2142), .CK(CLK), .Q(\REGISTERS[0][10] )
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n2141), .CK(CLK), .Q(\REGISTERS[0][9] ) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n2140), .CK(CLK), .Q(\REGISTERS[0][8] ) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n2139), .CK(CLK), .Q(\REGISTERS[0][7] ) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n2138), .CK(CLK), .Q(\REGISTERS[0][6] ) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n2137), .CK(CLK), .Q(\REGISTERS[0][5] ) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n2136), .CK(CLK), .Q(\REGISTERS[0][4] ) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n2135), .CK(CLK), .Q(\REGISTERS[0][3] ) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n2134), .CK(CLK), .Q(\REGISTERS[0][2] ) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n2133), .CK(CLK), .Q(\REGISTERS[0][1] ) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n2132), .CK(CLK), .Q(\REGISTERS[0][0] ) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n2131), .CK(CLK), .Q(\REGISTERS[1][31] )
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n2130), .CK(CLK), .Q(\REGISTERS[1][30] )
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n2129), .CK(CLK), .Q(\REGISTERS[1][29] )
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n2128), .CK(CLK), .Q(\REGISTERS[1][28] )
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n2127), .CK(CLK), .Q(\REGISTERS[1][27] )
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n2126), .CK(CLK), .Q(\REGISTERS[1][26] )
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n2125), .CK(CLK), .Q(\REGISTERS[1][25] )
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n2124), .CK(CLK), .Q(\REGISTERS[1][24] )
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n2123), .CK(CLK), .Q(\REGISTERS[1][23] )
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n2122), .CK(CLK), .Q(\REGISTERS[1][22] )
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n2121), .CK(CLK), .Q(\REGISTERS[1][21] )
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n2120), .CK(CLK), .Q(\REGISTERS[1][20] )
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n2119), .CK(CLK), .Q(\REGISTERS[1][19] )
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n2118), .CK(CLK), .Q(\REGISTERS[1][18] )
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n2117), .CK(CLK), .Q(\REGISTERS[1][17] )
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n2116), .CK(CLK), .Q(\REGISTERS[1][16] )
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n2115), .CK(CLK), .Q(\REGISTERS[1][15] )
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n2114), .CK(CLK), .Q(\REGISTERS[1][14] )
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n2113), .CK(CLK), .Q(\REGISTERS[1][13] )
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n2112), .CK(CLK), .Q(\REGISTERS[1][12] )
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n2111), .CK(CLK), .Q(\REGISTERS[1][11] )
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n2110), .CK(CLK), .Q(\REGISTERS[1][10] )
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n2109), .CK(CLK), .Q(\REGISTERS[1][9] ) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n2108), .CK(CLK), .Q(\REGISTERS[1][8] ) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n2107), .CK(CLK), .Q(\REGISTERS[1][7] ) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n2106), .CK(CLK), .Q(\REGISTERS[1][6] ) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n2105), .CK(CLK), .Q(\REGISTERS[1][5] ) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n2104), .CK(CLK), .Q(\REGISTERS[1][4] ) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n2103), .CK(CLK), .Q(\REGISTERS[1][3] ) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n2102), .CK(CLK), .Q(\REGISTERS[1][2] ) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n2101), .CK(CLK), .Q(\REGISTERS[1][1] ) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n2100), .CK(CLK), .Q(\REGISTERS[1][0] ) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n2099), .CK(CLK), .Q(\REGISTERS[2][31] )
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n2098), .CK(CLK), .Q(\REGISTERS[2][30] )
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n2097), .CK(CLK), .Q(\REGISTERS[2][29] )
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n2096), .CK(CLK), .Q(\REGISTERS[2][28] )
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n2095), .CK(CLK), .Q(\REGISTERS[2][27] )
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n2094), .CK(CLK), .Q(\REGISTERS[2][26] )
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n2093), .CK(CLK), .Q(\REGISTERS[2][25] )
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n2092), .CK(CLK), .Q(\REGISTERS[2][24] )
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n2091), .CK(CLK), .Q(\REGISTERS[2][23] )
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n2090), .CK(CLK), .Q(\REGISTERS[2][22] )
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n2089), .CK(CLK), .Q(\REGISTERS[2][21] )
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n2088), .CK(CLK), .Q(\REGISTERS[2][20] )
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n2087), .CK(CLK), .Q(\REGISTERS[2][19] )
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n2086), .CK(CLK), .Q(\REGISTERS[2][18] )
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n2085), .CK(CLK), .Q(\REGISTERS[2][17] )
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n2084), .CK(CLK), .Q(\REGISTERS[2][16] )
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n2083), .CK(CLK), .Q(\REGISTERS[2][15] )
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n2082), .CK(CLK), .Q(\REGISTERS[2][14] )
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n2081), .CK(CLK), .Q(\REGISTERS[2][13] )
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n2080), .CK(CLK), .Q(\REGISTERS[2][12] )
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n2079), .CK(CLK), .Q(\REGISTERS[2][11] )
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n2078), .CK(CLK), .Q(\REGISTERS[2][10] )
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n2077), .CK(CLK), .Q(\REGISTERS[2][9] ) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n2076), .CK(CLK), .Q(\REGISTERS[2][8] ) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n2075), .CK(CLK), .Q(\REGISTERS[2][7] ) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n2074), .CK(CLK), .Q(\REGISTERS[2][6] ) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n2073), .CK(CLK), .Q(\REGISTERS[2][5] ) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n2072), .CK(CLK), .Q(\REGISTERS[2][4] ) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n2071), .CK(CLK), .Q(\REGISTERS[2][3] ) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n2070), .CK(CLK), .Q(\REGISTERS[2][2] ) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n2069), .CK(CLK), .Q(\REGISTERS[2][1] ) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n2068), .CK(CLK), .Q(\REGISTERS[2][0] ) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n2067), .CK(CLK), .Q(\REGISTERS[3][31] )
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n2066), .CK(CLK), .Q(\REGISTERS[3][30] )
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n2065), .CK(CLK), .Q(\REGISTERS[3][29] )
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n2064), .CK(CLK), .Q(\REGISTERS[3][28] )
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n2063), .CK(CLK), .Q(\REGISTERS[3][27] )
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n2062), .CK(CLK), .Q(\REGISTERS[3][26] )
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n2061), .CK(CLK), .Q(\REGISTERS[3][25] )
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n2060), .CK(CLK), .Q(\REGISTERS[3][24] )
         );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n2059), .CK(CLK), .Q(\REGISTERS[3][23] )
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n2058), .CK(CLK), .Q(\REGISTERS[3][22] )
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n2057), .CK(CLK), .Q(\REGISTERS[3][21] )
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n2056), .CK(CLK), .Q(\REGISTERS[3][20] )
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n2055), .CK(CLK), .Q(\REGISTERS[3][19] )
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n2054), .CK(CLK), .Q(\REGISTERS[3][18] )
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n2053), .CK(CLK), .Q(\REGISTERS[3][17] )
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n2052), .CK(CLK), .Q(\REGISTERS[3][16] )
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n2051), .CK(CLK), .Q(\REGISTERS[3][15] )
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n2050), .CK(CLK), .Q(\REGISTERS[3][14] )
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n2049), .CK(CLK), .Q(\REGISTERS[3][13] )
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n2048), .CK(CLK), .Q(\REGISTERS[3][12] )
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n2047), .CK(CLK), .Q(\REGISTERS[3][11] )
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n2046), .CK(CLK), .Q(\REGISTERS[3][10] )
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n2045), .CK(CLK), .Q(\REGISTERS[3][9] ) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n2044), .CK(CLK), .Q(\REGISTERS[3][8] ) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n2043), .CK(CLK), .Q(\REGISTERS[3][7] ) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n2042), .CK(CLK), .Q(\REGISTERS[3][6] ) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n2041), .CK(CLK), .Q(\REGISTERS[3][5] ) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n2040), .CK(CLK), .Q(\REGISTERS[3][4] ) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n2039), .CK(CLK), .Q(\REGISTERS[3][3] ) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n2038), .CK(CLK), .Q(\REGISTERS[3][2] ) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n2037), .CK(CLK), .Q(\REGISTERS[3][1] ) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n2036), .CK(CLK), .Q(\REGISTERS[3][0] ) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n2035), .CK(CLK), .Q(\REGISTERS[4][31] )
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n2034), .CK(CLK), .Q(\REGISTERS[4][30] )
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n2033), .CK(CLK), .Q(\REGISTERS[4][29] )
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n2032), .CK(CLK), .Q(\REGISTERS[4][28] )
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n2031), .CK(CLK), .Q(\REGISTERS[4][27] )
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n2030), .CK(CLK), .Q(\REGISTERS[4][26] )
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n2029), .CK(CLK), .Q(\REGISTERS[4][25] )
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n2028), .CK(CLK), .Q(\REGISTERS[4][24] )
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n2027), .CK(CLK), .Q(\REGISTERS[4][23] )
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n2026), .CK(CLK), .Q(\REGISTERS[4][22] )
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n2025), .CK(CLK), .Q(\REGISTERS[4][21] )
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n2024), .CK(CLK), .Q(\REGISTERS[4][20] )
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n2023), .CK(CLK), .Q(\REGISTERS[4][19] )
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n2022), .CK(CLK), .Q(\REGISTERS[4][18] )
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n2021), .CK(CLK), .Q(\REGISTERS[4][17] )
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n2020), .CK(CLK), .Q(\REGISTERS[4][16] )
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n2019), .CK(CLK), .Q(\REGISTERS[4][15] )
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n2018), .CK(CLK), .Q(\REGISTERS[4][14] )
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n2017), .CK(CLK), .Q(\REGISTERS[4][13] )
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n2016), .CK(CLK), .Q(\REGISTERS[4][12] )
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n2015), .CK(CLK), .Q(\REGISTERS[4][11] )
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n2014), .CK(CLK), .Q(\REGISTERS[4][10] )
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n2013), .CK(CLK), .Q(\REGISTERS[4][9] ) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n2012), .CK(CLK), .Q(\REGISTERS[4][8] ) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n2011), .CK(CLK), .Q(\REGISTERS[4][7] ) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n2010), .CK(CLK), .Q(\REGISTERS[4][6] ) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n2009), .CK(CLK), .Q(\REGISTERS[4][5] ) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n2008), .CK(CLK), .Q(\REGISTERS[4][4] ) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n2007), .CK(CLK), .Q(\REGISTERS[4][3] ) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n2006), .CK(CLK), .Q(\REGISTERS[4][2] ) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n2005), .CK(CLK), .Q(\REGISTERS[4][1] ) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n2004), .CK(CLK), .Q(\REGISTERS[4][0] ) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n2003), .CK(CLK), .Q(\REGISTERS[5][31] )
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n2002), .CK(CLK), .Q(\REGISTERS[5][30] )
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n2001), .CK(CLK), .Q(\REGISTERS[5][29] )
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n2000), .CK(CLK), .Q(\REGISTERS[5][28] )
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n1999), .CK(CLK), .Q(\REGISTERS[5][27] )
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n1998), .CK(CLK), .Q(\REGISTERS[5][26] )
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n1997), .CK(CLK), .Q(\REGISTERS[5][25] )
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n1996), .CK(CLK), .Q(\REGISTERS[5][24] )
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n1995), .CK(CLK), .Q(\REGISTERS[5][23] )
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n1994), .CK(CLK), .Q(\REGISTERS[5][22] )
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n1993), .CK(CLK), .Q(\REGISTERS[5][21] )
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n1992), .CK(CLK), .Q(\REGISTERS[5][20] )
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n1991), .CK(CLK), .Q(\REGISTERS[5][19] )
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n1990), .CK(CLK), .Q(\REGISTERS[5][18] )
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n1989), .CK(CLK), .Q(\REGISTERS[5][17] )
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n1988), .CK(CLK), .Q(\REGISTERS[5][16] )
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n1987), .CK(CLK), .Q(\REGISTERS[5][15] )
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n1986), .CK(CLK), .Q(\REGISTERS[5][14] )
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n1985), .CK(CLK), .Q(\REGISTERS[5][13] )
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n1984), .CK(CLK), .Q(\REGISTERS[5][12] )
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n1983), .CK(CLK), .Q(\REGISTERS[5][11] )
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n1982), .CK(CLK), .Q(\REGISTERS[5][10] )
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n1981), .CK(CLK), .Q(\REGISTERS[5][9] ) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n1980), .CK(CLK), .Q(\REGISTERS[5][8] ) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n1979), .CK(CLK), .Q(\REGISTERS[5][7] ) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n1978), .CK(CLK), .Q(\REGISTERS[5][6] ) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n1977), .CK(CLK), .Q(\REGISTERS[5][5] ) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n1976), .CK(CLK), .Q(\REGISTERS[5][4] ) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n1975), .CK(CLK), .Q(\REGISTERS[5][3] ) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n1974), .CK(CLK), .Q(\REGISTERS[5][2] ) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n1973), .CK(CLK), .Q(\REGISTERS[5][1] ) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n1972), .CK(CLK), .Q(\REGISTERS[5][0] ) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n1971), .CK(CLK), .Q(\REGISTERS[6][31] )
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n1970), .CK(CLK), .Q(\REGISTERS[6][30] )
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n1969), .CK(CLK), .Q(\REGISTERS[6][29] )
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n1968), .CK(CLK), .Q(\REGISTERS[6][28] )
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n1967), .CK(CLK), .Q(\REGISTERS[6][27] )
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n1966), .CK(CLK), .Q(\REGISTERS[6][26] )
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n1965), .CK(CLK), .Q(\REGISTERS[6][25] )
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n1964), .CK(CLK), .Q(\REGISTERS[6][24] )
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n1963), .CK(CLK), .Q(\REGISTERS[6][23] )
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n1962), .CK(CLK), .Q(\REGISTERS[6][22] )
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n1961), .CK(CLK), .Q(\REGISTERS[6][21] )
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n1960), .CK(CLK), .Q(\REGISTERS[6][20] )
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n1959), .CK(CLK), .Q(\REGISTERS[6][19] )
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n1958), .CK(CLK), .Q(\REGISTERS[6][18] )
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n1957), .CK(CLK), .Q(\REGISTERS[6][17] )
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n1956), .CK(CLK), .Q(\REGISTERS[6][16] )
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n1955), .CK(CLK), .Q(\REGISTERS[6][15] )
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n1954), .CK(CLK), .Q(\REGISTERS[6][14] )
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n1953), .CK(CLK), .Q(\REGISTERS[6][13] )
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n1952), .CK(CLK), .Q(\REGISTERS[6][12] )
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n1951), .CK(CLK), .Q(\REGISTERS[6][11] )
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n1950), .CK(CLK), .Q(\REGISTERS[6][10] )
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n1949), .CK(CLK), .Q(\REGISTERS[6][9] ) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n1948), .CK(CLK), .Q(\REGISTERS[6][8] ) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n1947), .CK(CLK), .Q(\REGISTERS[6][7] ) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n1946), .CK(CLK), .Q(\REGISTERS[6][6] ) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n1945), .CK(CLK), .Q(\REGISTERS[6][5] ) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n1944), .CK(CLK), .Q(\REGISTERS[6][4] ) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n1943), .CK(CLK), .Q(\REGISTERS[6][3] ) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n1942), .CK(CLK), .Q(\REGISTERS[6][2] ) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n1941), .CK(CLK), .Q(\REGISTERS[6][1] ) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n1940), .CK(CLK), .Q(\REGISTERS[6][0] ) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n1939), .CK(CLK), .Q(\REGISTERS[7][31] )
         );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n1938), .CK(CLK), .Q(\REGISTERS[7][30] )
         );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n1937), .CK(CLK), .Q(\REGISTERS[7][29] )
         );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n1936), .CK(CLK), .Q(\REGISTERS[7][28] )
         );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n1935), .CK(CLK), .Q(\REGISTERS[7][27] )
         );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n1934), .CK(CLK), .Q(\REGISTERS[7][26] )
         );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n1933), .CK(CLK), .Q(\REGISTERS[7][25] )
         );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n1932), .CK(CLK), .Q(\REGISTERS[7][24] )
         );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n1931), .CK(CLK), .Q(\REGISTERS[7][23] )
         );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n1930), .CK(CLK), .Q(\REGISTERS[7][22] )
         );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n1929), .CK(CLK), .Q(\REGISTERS[7][21] )
         );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n1928), .CK(CLK), .Q(\REGISTERS[7][20] )
         );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n1927), .CK(CLK), .Q(\REGISTERS[7][19] )
         );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n1926), .CK(CLK), .Q(\REGISTERS[7][18] )
         );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n1925), .CK(CLK), .Q(\REGISTERS[7][17] )
         );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n1924), .CK(CLK), .Q(\REGISTERS[7][16] )
         );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n1923), .CK(CLK), .Q(\REGISTERS[7][15] )
         );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n1922), .CK(CLK), .Q(\REGISTERS[7][14] )
         );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n1921), .CK(CLK), .Q(\REGISTERS[7][13] )
         );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n1920), .CK(CLK), .Q(\REGISTERS[7][12] )
         );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n1919), .CK(CLK), .Q(\REGISTERS[7][11] )
         );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n1918), .CK(CLK), .Q(\REGISTERS[7][10] )
         );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n1917), .CK(CLK), .Q(\REGISTERS[7][9] ) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n1916), .CK(CLK), .Q(\REGISTERS[7][8] ) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n1915), .CK(CLK), .Q(\REGISTERS[7][7] ) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n1914), .CK(CLK), .Q(\REGISTERS[7][6] ) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n1913), .CK(CLK), .Q(\REGISTERS[7][5] ) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n1912), .CK(CLK), .Q(\REGISTERS[7][4] ) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n1911), .CK(CLK), .Q(\REGISTERS[7][3] ) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n1910), .CK(CLK), .Q(\REGISTERS[7][2] ) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n1909), .CK(CLK), .Q(\REGISTERS[7][1] ) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n1908), .CK(CLK), .Q(\REGISTERS[7][0] ) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n1907), .CK(CLK), .Q(\REGISTERS[8][31] )
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n1906), .CK(CLK), .Q(\REGISTERS[8][30] )
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n1905), .CK(CLK), .Q(\REGISTERS[8][29] )
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n1904), .CK(CLK), .Q(\REGISTERS[8][28] )
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n1903), .CK(CLK), .Q(\REGISTERS[8][27] )
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n1902), .CK(CLK), .Q(\REGISTERS[8][26] )
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n1901), .CK(CLK), .Q(\REGISTERS[8][25] )
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n1900), .CK(CLK), .Q(\REGISTERS[8][24] )
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n1899), .CK(CLK), .Q(\REGISTERS[8][23] )
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n1898), .CK(CLK), .Q(\REGISTERS[8][22] )
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n1897), .CK(CLK), .Q(\REGISTERS[8][21] )
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n1896), .CK(CLK), .Q(\REGISTERS[8][20] )
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n1895), .CK(CLK), .Q(\REGISTERS[8][19] )
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n1894), .CK(CLK), .Q(\REGISTERS[8][18] )
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n1893), .CK(CLK), .Q(\REGISTERS[8][17] )
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n1892), .CK(CLK), .Q(\REGISTERS[8][16] )
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n1891), .CK(CLK), .Q(\REGISTERS[8][15] )
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n1890), .CK(CLK), .Q(\REGISTERS[8][14] )
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n1889), .CK(CLK), .Q(\REGISTERS[8][13] )
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n1888), .CK(CLK), .Q(\REGISTERS[8][12] )
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n1887), .CK(CLK), .Q(\REGISTERS[8][11] )
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n1886), .CK(CLK), .Q(\REGISTERS[8][10] )
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n1885), .CK(CLK), .Q(\REGISTERS[8][9] ) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n1884), .CK(CLK), .Q(\REGISTERS[8][8] ) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n1883), .CK(CLK), .Q(\REGISTERS[8][7] ) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n1882), .CK(CLK), .Q(\REGISTERS[8][6] ) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n1881), .CK(CLK), .Q(\REGISTERS[8][5] ) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n1880), .CK(CLK), .Q(\REGISTERS[8][4] ) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n1879), .CK(CLK), .Q(\REGISTERS[8][3] ) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n1878), .CK(CLK), .Q(\REGISTERS[8][2] ) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n1877), .CK(CLK), .Q(\REGISTERS[8][1] ) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n1876), .CK(CLK), .Q(\REGISTERS[8][0] ) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n1875), .CK(CLK), .Q(\REGISTERS[9][31] )
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n1874), .CK(CLK), .Q(\REGISTERS[9][30] )
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n1873), .CK(CLK), .Q(\REGISTERS[9][29] )
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n1872), .CK(CLK), .Q(\REGISTERS[9][28] )
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n1871), .CK(CLK), .Q(\REGISTERS[9][27] )
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n1870), .CK(CLK), .Q(\REGISTERS[9][26] )
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n1869), .CK(CLK), .Q(\REGISTERS[9][25] )
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n1868), .CK(CLK), .Q(\REGISTERS[9][24] )
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n1867), .CK(CLK), .Q(\REGISTERS[9][23] )
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n1866), .CK(CLK), .Q(\REGISTERS[9][22] )
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n1865), .CK(CLK), .Q(\REGISTERS[9][21] )
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n1864), .CK(CLK), .Q(\REGISTERS[9][20] )
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n1863), .CK(CLK), .Q(\REGISTERS[9][19] )
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n1862), .CK(CLK), .Q(\REGISTERS[9][18] )
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n1861), .CK(CLK), .Q(\REGISTERS[9][17] )
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n1860), .CK(CLK), .Q(\REGISTERS[9][16] )
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n1859), .CK(CLK), .Q(\REGISTERS[9][15] )
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n1858), .CK(CLK), .Q(\REGISTERS[9][14] )
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n1857), .CK(CLK), .Q(\REGISTERS[9][13] )
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n1856), .CK(CLK), .Q(\REGISTERS[9][12] )
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n1855), .CK(CLK), .Q(\REGISTERS[9][11] )
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n1854), .CK(CLK), .Q(\REGISTERS[9][10] )
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n1853), .CK(CLK), .Q(\REGISTERS[9][9] ) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n1852), .CK(CLK), .Q(\REGISTERS[9][8] ) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n1851), .CK(CLK), .Q(\REGISTERS[9][7] ) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n1850), .CK(CLK), .Q(\REGISTERS[9][6] ) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n1849), .CK(CLK), .Q(\REGISTERS[9][5] ) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n1848), .CK(CLK), .Q(\REGISTERS[9][4] ) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n1847), .CK(CLK), .Q(\REGISTERS[9][3] ) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n1846), .CK(CLK), .Q(\REGISTERS[9][2] ) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n1845), .CK(CLK), .Q(\REGISTERS[9][1] ) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n1844), .CK(CLK), .Q(\REGISTERS[9][0] ) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n1843), .CK(CLK), .Q(\REGISTERS[10][31] ) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n1842), .CK(CLK), .Q(\REGISTERS[10][30] ) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n1841), .CK(CLK), .Q(\REGISTERS[10][29] ) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n1840), .CK(CLK), .Q(\REGISTERS[10][28] ) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n1839), .CK(CLK), .Q(\REGISTERS[10][27] ) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n1838), .CK(CLK), .Q(\REGISTERS[10][26] ) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n1837), .CK(CLK), .Q(\REGISTERS[10][25] ) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n1836), .CK(CLK), .Q(\REGISTERS[10][24] ) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n1835), .CK(CLK), .Q(\REGISTERS[10][23] ) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n1834), .CK(CLK), .Q(\REGISTERS[10][22] ) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n1833), .CK(CLK), .Q(\REGISTERS[10][21] ) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n1832), .CK(CLK), .Q(\REGISTERS[10][20] ) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n1831), .CK(CLK), .Q(\REGISTERS[10][19] ) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n1830), .CK(CLK), .Q(\REGISTERS[10][18] ) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n1829), .CK(CLK), .Q(\REGISTERS[10][17] ) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n1828), .CK(CLK), .Q(\REGISTERS[10][16] ) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n1827), .CK(CLK), .Q(\REGISTERS[10][15] ) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n1826), .CK(CLK), .Q(\REGISTERS[10][14] ) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n1825), .CK(CLK), .Q(\REGISTERS[10][13] ) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n1824), .CK(CLK), .Q(\REGISTERS[10][12] ) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n1823), .CK(CLK), .Q(\REGISTERS[10][11] ) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n1822), .CK(CLK), .Q(\REGISTERS[10][10] ) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n1821), .CK(CLK), .Q(\REGISTERS[10][9] )
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n1820), .CK(CLK), .Q(\REGISTERS[10][8] )
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n1819), .CK(CLK), .Q(\REGISTERS[10][7] )
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n1818), .CK(CLK), .Q(\REGISTERS[10][6] )
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n1817), .CK(CLK), .Q(\REGISTERS[10][5] )
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n1816), .CK(CLK), .Q(\REGISTERS[10][4] )
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n1815), .CK(CLK), .Q(\REGISTERS[10][3] )
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n1814), .CK(CLK), .Q(\REGISTERS[10][2] )
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n1813), .CK(CLK), .Q(\REGISTERS[10][1] )
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n1812), .CK(CLK), .Q(\REGISTERS[10][0] )
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n1811), .CK(CLK), .Q(\REGISTERS[11][31] ) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n1810), .CK(CLK), .Q(\REGISTERS[11][30] ) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n1809), .CK(CLK), .Q(\REGISTERS[11][29] ) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n1808), .CK(CLK), .Q(\REGISTERS[11][28] ) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n1807), .CK(CLK), .Q(\REGISTERS[11][27] ) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n1806), .CK(CLK), .Q(\REGISTERS[11][26] ) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n1805), .CK(CLK), .Q(\REGISTERS[11][25] ) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n1804), .CK(CLK), .Q(\REGISTERS[11][24] ) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n1803), .CK(CLK), .Q(\REGISTERS[11][23] ) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n1802), .CK(CLK), .Q(\REGISTERS[11][22] ) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n1801), .CK(CLK), .Q(\REGISTERS[11][21] ) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n1800), .CK(CLK), .Q(\REGISTERS[11][20] ) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n1799), .CK(CLK), .Q(\REGISTERS[11][19] ) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n1798), .CK(CLK), .Q(\REGISTERS[11][18] ) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n1797), .CK(CLK), .Q(\REGISTERS[11][17] ) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n1796), .CK(CLK), .Q(\REGISTERS[11][16] ) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n1795), .CK(CLK), .Q(\REGISTERS[11][15] ) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n1794), .CK(CLK), .Q(\REGISTERS[11][14] ) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n1793), .CK(CLK), .Q(\REGISTERS[11][13] ) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n1792), .CK(CLK), .Q(\REGISTERS[11][12] ) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n1791), .CK(CLK), .Q(\REGISTERS[11][11] ) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n1790), .CK(CLK), .Q(\REGISTERS[11][10] ) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n1789), .CK(CLK), .Q(\REGISTERS[11][9] )
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n1788), .CK(CLK), .Q(\REGISTERS[11][8] )
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n1787), .CK(CLK), .Q(\REGISTERS[11][7] )
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n1786), .CK(CLK), .Q(\REGISTERS[11][6] )
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n1785), .CK(CLK), .Q(\REGISTERS[11][5] )
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n1784), .CK(CLK), .Q(\REGISTERS[11][4] )
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n1783), .CK(CLK), .Q(\REGISTERS[11][3] )
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n1782), .CK(CLK), .Q(\REGISTERS[11][2] )
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n1781), .CK(CLK), .Q(\REGISTERS[11][1] )
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n1780), .CK(CLK), .Q(\REGISTERS[11][0] )
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n1779), .CK(CLK), .Q(\REGISTERS[12][31] ) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n1778), .CK(CLK), .Q(\REGISTERS[12][30] ) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n1777), .CK(CLK), .Q(\REGISTERS[12][29] ) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n1776), .CK(CLK), .Q(\REGISTERS[12][28] ) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n1775), .CK(CLK), .Q(\REGISTERS[12][27] ) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n1774), .CK(CLK), .Q(\REGISTERS[12][26] ) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n1773), .CK(CLK), .Q(\REGISTERS[12][25] ) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n1772), .CK(CLK), .Q(\REGISTERS[12][24] ) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n1771), .CK(CLK), .Q(\REGISTERS[12][23] ) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n1770), .CK(CLK), .Q(\REGISTERS[12][22] ) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n1769), .CK(CLK), .Q(\REGISTERS[12][21] ) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n1768), .CK(CLK), .Q(\REGISTERS[12][20] ) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n1767), .CK(CLK), .Q(\REGISTERS[12][19] ) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n1766), .CK(CLK), .Q(\REGISTERS[12][18] ) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n1765), .CK(CLK), .Q(\REGISTERS[12][17] ) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n1764), .CK(CLK), .Q(\REGISTERS[12][16] ) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n1763), .CK(CLK), .Q(\REGISTERS[12][15] ) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n1762), .CK(CLK), .Q(\REGISTERS[12][14] ) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n1761), .CK(CLK), .Q(\REGISTERS[12][13] ) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n1760), .CK(CLK), .Q(\REGISTERS[12][12] ) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n1759), .CK(CLK), .Q(\REGISTERS[12][11] ) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n1758), .CK(CLK), .Q(\REGISTERS[12][10] ) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n1757), .CK(CLK), .Q(\REGISTERS[12][9] )
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n1756), .CK(CLK), .Q(\REGISTERS[12][8] )
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n1755), .CK(CLK), .Q(\REGISTERS[12][7] )
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n1754), .CK(CLK), .Q(\REGISTERS[12][6] )
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n1753), .CK(CLK), .Q(\REGISTERS[12][5] )
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n1752), .CK(CLK), .Q(\REGISTERS[12][4] )
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n1751), .CK(CLK), .Q(\REGISTERS[12][3] )
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n1750), .CK(CLK), .Q(\REGISTERS[12][2] )
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n1749), .CK(CLK), .Q(\REGISTERS[12][1] )
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n1748), .CK(CLK), .Q(\REGISTERS[12][0] )
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n1747), .CK(CLK), .Q(\REGISTERS[13][31] ) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n1746), .CK(CLK), .Q(\REGISTERS[13][30] ) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n1745), .CK(CLK), .Q(\REGISTERS[13][29] ) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n1744), .CK(CLK), .Q(\REGISTERS[13][28] ) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n1743), .CK(CLK), .Q(\REGISTERS[13][27] ) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n1742), .CK(CLK), .Q(\REGISTERS[13][26] ) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n1741), .CK(CLK), .Q(\REGISTERS[13][25] ) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n1740), .CK(CLK), .Q(\REGISTERS[13][24] ) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n1739), .CK(CLK), .Q(\REGISTERS[13][23] ) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n1738), .CK(CLK), .Q(\REGISTERS[13][22] ) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n1737), .CK(CLK), .Q(\REGISTERS[13][21] ) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n1736), .CK(CLK), .Q(\REGISTERS[13][20] ) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n1735), .CK(CLK), .Q(\REGISTERS[13][19] ) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n1734), .CK(CLK), .Q(\REGISTERS[13][18] ) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n1733), .CK(CLK), .Q(\REGISTERS[13][17] ) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n1732), .CK(CLK), .Q(\REGISTERS[13][16] ) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n1731), .CK(CLK), .Q(\REGISTERS[13][15] ) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n1730), .CK(CLK), .Q(\REGISTERS[13][14] ) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n1729), .CK(CLK), .Q(\REGISTERS[13][13] ) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n1728), .CK(CLK), .Q(\REGISTERS[13][12] ) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n1727), .CK(CLK), .Q(\REGISTERS[13][11] ) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n1726), .CK(CLK), .Q(\REGISTERS[13][10] ) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n1725), .CK(CLK), .Q(\REGISTERS[13][9] )
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n1724), .CK(CLK), .Q(\REGISTERS[13][8] )
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n1723), .CK(CLK), .Q(\REGISTERS[13][7] )
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n1722), .CK(CLK), .Q(\REGISTERS[13][6] )
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n1721), .CK(CLK), .Q(\REGISTERS[13][5] )
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n1720), .CK(CLK), .Q(\REGISTERS[13][4] )
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n1719), .CK(CLK), .Q(\REGISTERS[13][3] )
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n1718), .CK(CLK), .Q(\REGISTERS[13][2] )
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n1717), .CK(CLK), .Q(\REGISTERS[13][1] )
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n1716), .CK(CLK), .Q(\REGISTERS[13][0] )
         );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n1715), .CK(CLK), .Q(\REGISTERS[14][31] ) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n1714), .CK(CLK), .Q(\REGISTERS[14][30] ) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n1713), .CK(CLK), .Q(\REGISTERS[14][29] ) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n1712), .CK(CLK), .Q(\REGISTERS[14][28] ) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n1711), .CK(CLK), .Q(\REGISTERS[14][27] ) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n1710), .CK(CLK), .Q(\REGISTERS[14][26] ) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n1709), .CK(CLK), .Q(\REGISTERS[14][25] ) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n1708), .CK(CLK), .Q(\REGISTERS[14][24] ) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n1707), .CK(CLK), .Q(\REGISTERS[14][23] ) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n1706), .CK(CLK), .Q(\REGISTERS[14][22] ) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n1705), .CK(CLK), .Q(\REGISTERS[14][21] ) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n1704), .CK(CLK), .Q(\REGISTERS[14][20] ) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n1703), .CK(CLK), .Q(\REGISTERS[14][19] ) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n1702), .CK(CLK), .Q(\REGISTERS[14][18] ) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n1701), .CK(CLK), .Q(\REGISTERS[14][17] ) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n1700), .CK(CLK), .Q(\REGISTERS[14][16] ) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n1699), .CK(CLK), .Q(\REGISTERS[14][15] ) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n1698), .CK(CLK), .Q(\REGISTERS[14][14] ) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n1697), .CK(CLK), .Q(\REGISTERS[14][13] ) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n1696), .CK(CLK), .Q(\REGISTERS[14][12] ) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n1695), .CK(CLK), .Q(\REGISTERS[14][11] ) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n1694), .CK(CLK), .Q(\REGISTERS[14][10] ) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n1693), .CK(CLK), .Q(\REGISTERS[14][9] )
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n1692), .CK(CLK), .Q(\REGISTERS[14][8] )
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n1691), .CK(CLK), .Q(\REGISTERS[14][7] )
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n1690), .CK(CLK), .Q(\REGISTERS[14][6] )
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n1689), .CK(CLK), .Q(\REGISTERS[14][5] )
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n1688), .CK(CLK), .Q(\REGISTERS[14][4] )
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n1687), .CK(CLK), .Q(\REGISTERS[14][3] )
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n1686), .CK(CLK), .Q(\REGISTERS[14][2] )
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n1685), .CK(CLK), .Q(\REGISTERS[14][1] )
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n1684), .CK(CLK), .Q(\REGISTERS[14][0] )
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n1683), .CK(CLK), .Q(\REGISTERS[15][31] ) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n1682), .CK(CLK), .Q(\REGISTERS[15][30] ) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n1681), .CK(CLK), .Q(\REGISTERS[15][29] ) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n1680), .CK(CLK), .Q(\REGISTERS[15][28] ) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n1679), .CK(CLK), .Q(\REGISTERS[15][27] ) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n1678), .CK(CLK), .Q(\REGISTERS[15][26] ) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n1677), .CK(CLK), .Q(\REGISTERS[15][25] ) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n1676), .CK(CLK), .Q(\REGISTERS[15][24] ) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n1675), .CK(CLK), .Q(\REGISTERS[15][23] ) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n1674), .CK(CLK), .Q(\REGISTERS[15][22] ) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n1673), .CK(CLK), .Q(\REGISTERS[15][21] ) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n1672), .CK(CLK), .Q(\REGISTERS[15][20] ) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n1671), .CK(CLK), .Q(\REGISTERS[15][19] ) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n1670), .CK(CLK), .Q(\REGISTERS[15][18] ) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n1669), .CK(CLK), .Q(\REGISTERS[15][17] ) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n1668), .CK(CLK), .Q(\REGISTERS[15][16] ) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n1667), .CK(CLK), .Q(\REGISTERS[15][15] ) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n1666), .CK(CLK), .Q(\REGISTERS[15][14] ) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n1665), .CK(CLK), .Q(\REGISTERS[15][13] ) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n1664), .CK(CLK), .Q(\REGISTERS[15][12] ) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n1663), .CK(CLK), .Q(\REGISTERS[15][11] ) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n1662), .CK(CLK), .Q(\REGISTERS[15][10] ) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n1661), .CK(CLK), .Q(\REGISTERS[15][9] )
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n1660), .CK(CLK), .Q(\REGISTERS[15][8] )
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n1659), .CK(CLK), .Q(\REGISTERS[15][7] )
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n1658), .CK(CLK), .Q(\REGISTERS[15][6] )
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n1657), .CK(CLK), .Q(\REGISTERS[15][5] )
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n1656), .CK(CLK), .Q(\REGISTERS[15][4] )
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n1655), .CK(CLK), .Q(\REGISTERS[15][3] )
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n1654), .CK(CLK), .Q(\REGISTERS[15][2] )
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n1653), .CK(CLK), .Q(\REGISTERS[15][1] )
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n1652), .CK(CLK), .Q(\REGISTERS[15][0] )
         );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n1651), .CK(CLK), .Q(\REGISTERS[16][31] ) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n1650), .CK(CLK), .Q(\REGISTERS[16][30] ) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n1649), .CK(CLK), .Q(\REGISTERS[16][29] ) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n1648), .CK(CLK), .Q(\REGISTERS[16][28] ) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n1647), .CK(CLK), .Q(\REGISTERS[16][27] ) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n1646), .CK(CLK), .Q(\REGISTERS[16][26] ) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n1645), .CK(CLK), .Q(\REGISTERS[16][25] ) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n1644), .CK(CLK), .Q(\REGISTERS[16][24] ) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n1643), .CK(CLK), .Q(\REGISTERS[16][23] ) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n1642), .CK(CLK), .Q(\REGISTERS[16][22] ) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n1641), .CK(CLK), .Q(\REGISTERS[16][21] ) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n1640), .CK(CLK), .Q(\REGISTERS[16][20] ) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n1639), .CK(CLK), .Q(\REGISTERS[16][19] ) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n1638), .CK(CLK), .Q(\REGISTERS[16][18] ) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n1637), .CK(CLK), .Q(\REGISTERS[16][17] ) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n1636), .CK(CLK), .Q(\REGISTERS[16][16] ) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n1635), .CK(CLK), .Q(\REGISTERS[16][15] ) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n1634), .CK(CLK), .Q(\REGISTERS[16][14] ) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n1633), .CK(CLK), .Q(\REGISTERS[16][13] ) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n1632), .CK(CLK), .Q(\REGISTERS[16][12] ) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n1631), .CK(CLK), .Q(\REGISTERS[16][11] ) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n1630), .CK(CLK), .Q(\REGISTERS[16][10] ) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n1629), .CK(CLK), .Q(\REGISTERS[16][9] )
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n1628), .CK(CLK), .Q(\REGISTERS[16][8] )
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n1627), .CK(CLK), .Q(\REGISTERS[16][7] )
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n1626), .CK(CLK), .Q(\REGISTERS[16][6] )
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n1625), .CK(CLK), .Q(\REGISTERS[16][5] )
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n1624), .CK(CLK), .Q(\REGISTERS[16][4] )
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n1623), .CK(CLK), .Q(\REGISTERS[16][3] )
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n1622), .CK(CLK), .Q(\REGISTERS[16][2] )
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n1621), .CK(CLK), .Q(\REGISTERS[16][1] )
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n1620), .CK(CLK), .Q(\REGISTERS[16][0] )
         );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n1619), .CK(CLK), .Q(\REGISTERS[17][31] ) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n1618), .CK(CLK), .Q(\REGISTERS[17][30] ) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n1617), .CK(CLK), .Q(\REGISTERS[17][29] ) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n1616), .CK(CLK), .Q(\REGISTERS[17][28] ) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n1615), .CK(CLK), .Q(\REGISTERS[17][27] ) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n1614), .CK(CLK), .Q(\REGISTERS[17][26] ) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n1613), .CK(CLK), .Q(\REGISTERS[17][25] ) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n1612), .CK(CLK), .Q(\REGISTERS[17][24] ) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n1611), .CK(CLK), .Q(\REGISTERS[17][23] ) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n1610), .CK(CLK), .Q(\REGISTERS[17][22] ) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n1609), .CK(CLK), .Q(\REGISTERS[17][21] ) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n1608), .CK(CLK), .Q(\REGISTERS[17][20] ) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n1607), .CK(CLK), .Q(\REGISTERS[17][19] ) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n1606), .CK(CLK), .Q(\REGISTERS[17][18] ) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n1605), .CK(CLK), .Q(\REGISTERS[17][17] ) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n1604), .CK(CLK), .Q(\REGISTERS[17][16] ) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n1603), .CK(CLK), .Q(\REGISTERS[17][15] ) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n1602), .CK(CLK), .Q(\REGISTERS[17][14] ) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n1601), .CK(CLK), .Q(\REGISTERS[17][13] ) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n1600), .CK(CLK), .Q(\REGISTERS[17][12] ) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n1599), .CK(CLK), .Q(\REGISTERS[17][11] ) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n1598), .CK(CLK), .Q(\REGISTERS[17][10] ) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n1597), .CK(CLK), .Q(\REGISTERS[17][9] )
         );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n1596), .CK(CLK), .Q(\REGISTERS[17][8] )
         );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n1595), .CK(CLK), .Q(\REGISTERS[17][7] )
         );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n1594), .CK(CLK), .Q(\REGISTERS[17][6] )
         );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n1593), .CK(CLK), .Q(\REGISTERS[17][5] )
         );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n1592), .CK(CLK), .Q(\REGISTERS[17][4] )
         );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n1591), .CK(CLK), .Q(\REGISTERS[17][3] )
         );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n1590), .CK(CLK), .Q(\REGISTERS[17][2] )
         );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n1589), .CK(CLK), .Q(\REGISTERS[17][1] )
         );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n1588), .CK(CLK), .Q(\REGISTERS[17][0] )
         );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n1587), .CK(CLK), .Q(\REGISTERS[18][31] ) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n1586), .CK(CLK), .Q(\REGISTERS[18][30] ) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n1585), .CK(CLK), .Q(\REGISTERS[18][29] ) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n1584), .CK(CLK), .Q(\REGISTERS[18][28] ) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n1583), .CK(CLK), .Q(\REGISTERS[18][27] ) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n1582), .CK(CLK), .Q(\REGISTERS[18][26] ) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n1581), .CK(CLK), .Q(\REGISTERS[18][25] ) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n1580), .CK(CLK), .Q(\REGISTERS[18][24] ) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n1579), .CK(CLK), .Q(\REGISTERS[18][23] ) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n1578), .CK(CLK), .Q(\REGISTERS[18][22] ) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n1577), .CK(CLK), .Q(\REGISTERS[18][21] ) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n1576), .CK(CLK), .Q(\REGISTERS[18][20] ) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n1575), .CK(CLK), .Q(\REGISTERS[18][19] ) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n1574), .CK(CLK), .Q(\REGISTERS[18][18] ) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n1573), .CK(CLK), .Q(\REGISTERS[18][17] ) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n1572), .CK(CLK), .Q(\REGISTERS[18][16] ) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n1571), .CK(CLK), .Q(\REGISTERS[18][15] ) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n1570), .CK(CLK), .Q(\REGISTERS[18][14] ) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n1569), .CK(CLK), .Q(\REGISTERS[18][13] ) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n1568), .CK(CLK), .Q(\REGISTERS[18][12] ) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n1567), .CK(CLK), .Q(\REGISTERS[18][11] ) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n1566), .CK(CLK), .Q(\REGISTERS[18][10] ) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n1565), .CK(CLK), .Q(\REGISTERS[18][9] )
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n1564), .CK(CLK), .Q(\REGISTERS[18][8] )
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n1563), .CK(CLK), .Q(\REGISTERS[18][7] )
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n1562), .CK(CLK), .Q(\REGISTERS[18][6] )
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n1561), .CK(CLK), .Q(\REGISTERS[18][5] )
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n1560), .CK(CLK), .Q(\REGISTERS[18][4] )
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n1559), .CK(CLK), .Q(\REGISTERS[18][3] )
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n1558), .CK(CLK), .Q(\REGISTERS[18][2] )
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n1557), .CK(CLK), .Q(\REGISTERS[18][1] )
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n1556), .CK(CLK), .Q(\REGISTERS[18][0] )
         );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n1555), .CK(CLK), .Q(\REGISTERS[19][31] ) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n1554), .CK(CLK), .Q(\REGISTERS[19][30] ) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n1553), .CK(CLK), .Q(\REGISTERS[19][29] ) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n1552), .CK(CLK), .Q(\REGISTERS[19][28] ) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n1551), .CK(CLK), .Q(\REGISTERS[19][27] ) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n1550), .CK(CLK), .Q(\REGISTERS[19][26] ) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n1549), .CK(CLK), .Q(\REGISTERS[19][25] ) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n1548), .CK(CLK), .Q(\REGISTERS[19][24] ) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n1547), .CK(CLK), .Q(\REGISTERS[19][23] ) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n1546), .CK(CLK), .Q(\REGISTERS[19][22] ) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n1545), .CK(CLK), .Q(\REGISTERS[19][21] ) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n1544), .CK(CLK), .Q(\REGISTERS[19][20] ) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n1543), .CK(CLK), .Q(\REGISTERS[19][19] ) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n1542), .CK(CLK), .Q(\REGISTERS[19][18] ) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n1541), .CK(CLK), .Q(\REGISTERS[19][17] ) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n1540), .CK(CLK), .Q(\REGISTERS[19][16] ) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n1539), .CK(CLK), .Q(\REGISTERS[19][15] ) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n1538), .CK(CLK), .Q(\REGISTERS[19][14] ) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n1537), .CK(CLK), .Q(\REGISTERS[19][13] ) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n1536), .CK(CLK), .Q(\REGISTERS[19][12] ) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n1535), .CK(CLK), .Q(\REGISTERS[19][11] ) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n1534), .CK(CLK), .Q(\REGISTERS[19][10] ) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n1533), .CK(CLK), .Q(\REGISTERS[19][9] )
         );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n1532), .CK(CLK), .Q(\REGISTERS[19][8] )
         );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n1531), .CK(CLK), .Q(\REGISTERS[19][7] )
         );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n1530), .CK(CLK), .Q(\REGISTERS[19][6] )
         );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n1529), .CK(CLK), .Q(\REGISTERS[19][5] )
         );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n1528), .CK(CLK), .Q(\REGISTERS[19][4] )
         );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n1527), .CK(CLK), .Q(\REGISTERS[19][3] )
         );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n1526), .CK(CLK), .Q(\REGISTERS[19][2] )
         );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n1525), .CK(CLK), .Q(\REGISTERS[19][1] )
         );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n1524), .CK(CLK), .Q(\REGISTERS[19][0] )
         );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n1523), .CK(CLK), .Q(\REGISTERS[20][31] ) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n1522), .CK(CLK), .Q(\REGISTERS[20][30] ) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n1521), .CK(CLK), .Q(\REGISTERS[20][29] ) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n1520), .CK(CLK), .Q(\REGISTERS[20][28] ) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n1519), .CK(CLK), .Q(\REGISTERS[20][27] ) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n1518), .CK(CLK), .Q(\REGISTERS[20][26] ) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n1517), .CK(CLK), .Q(\REGISTERS[20][25] ) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n1516), .CK(CLK), .Q(\REGISTERS[20][24] ) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n1515), .CK(CLK), .Q(\REGISTERS[20][23] ) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n1514), .CK(CLK), .Q(\REGISTERS[20][22] ) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n1513), .CK(CLK), .Q(\REGISTERS[20][21] ) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n1512), .CK(CLK), .Q(\REGISTERS[20][20] ) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n1511), .CK(CLK), .Q(\REGISTERS[20][19] ) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n1510), .CK(CLK), .Q(\REGISTERS[20][18] ) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n1509), .CK(CLK), .Q(\REGISTERS[20][17] ) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n1508), .CK(CLK), .Q(\REGISTERS[20][16] ) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n1507), .CK(CLK), .Q(\REGISTERS[20][15] ) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n1506), .CK(CLK), .Q(\REGISTERS[20][14] ) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n1505), .CK(CLK), .Q(\REGISTERS[20][13] ) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n1504), .CK(CLK), .Q(\REGISTERS[20][12] ) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n1503), .CK(CLK), .Q(\REGISTERS[20][11] ) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n1502), .CK(CLK), .Q(\REGISTERS[20][10] ) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n1501), .CK(CLK), .Q(\REGISTERS[20][9] )
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n1500), .CK(CLK), .Q(\REGISTERS[20][8] )
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n1499), .CK(CLK), .Q(\REGISTERS[20][7] )
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n1498), .CK(CLK), .Q(\REGISTERS[20][6] )
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n1497), .CK(CLK), .Q(\REGISTERS[20][5] )
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n1496), .CK(CLK), .Q(\REGISTERS[20][4] )
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n1495), .CK(CLK), .Q(\REGISTERS[20][3] )
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n1494), .CK(CLK), .Q(\REGISTERS[20][2] )
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n1493), .CK(CLK), .Q(\REGISTERS[20][1] )
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n1492), .CK(CLK), .Q(\REGISTERS[20][0] )
         );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n1491), .CK(CLK), .Q(\REGISTERS[21][31] ) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n1490), .CK(CLK), .Q(\REGISTERS[21][30] ) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n1489), .CK(CLK), .Q(\REGISTERS[21][29] ) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n1488), .CK(CLK), .Q(\REGISTERS[21][28] ) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n1487), .CK(CLK), .Q(\REGISTERS[21][27] ) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n1486), .CK(CLK), .Q(\REGISTERS[21][26] ) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n1485), .CK(CLK), .Q(\REGISTERS[21][25] ) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n1484), .CK(CLK), .Q(\REGISTERS[21][24] ) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n1483), .CK(CLK), .Q(\REGISTERS[21][23] ) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n1482), .CK(CLK), .Q(\REGISTERS[21][22] ) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n1481), .CK(CLK), .Q(\REGISTERS[21][21] ) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n1480), .CK(CLK), .Q(\REGISTERS[21][20] ) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n1479), .CK(CLK), .Q(\REGISTERS[21][19] ) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n1478), .CK(CLK), .Q(\REGISTERS[21][18] ) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n1477), .CK(CLK), .Q(\REGISTERS[21][17] ) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n1476), .CK(CLK), .Q(\REGISTERS[21][16] ) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n1475), .CK(CLK), .Q(\REGISTERS[21][15] ) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n1474), .CK(CLK), .Q(\REGISTERS[21][14] ) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n1473), .CK(CLK), .Q(\REGISTERS[21][13] ) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n1472), .CK(CLK), .Q(\REGISTERS[21][12] ) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n1471), .CK(CLK), .Q(\REGISTERS[21][11] ) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n1470), .CK(CLK), .Q(\REGISTERS[21][10] ) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n1469), .CK(CLK), .Q(\REGISTERS[21][9] )
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n1468), .CK(CLK), .Q(\REGISTERS[21][8] )
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n1467), .CK(CLK), .Q(\REGISTERS[21][7] )
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n1466), .CK(CLK), .Q(\REGISTERS[21][6] )
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n1465), .CK(CLK), .Q(\REGISTERS[21][5] )
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n1464), .CK(CLK), .Q(\REGISTERS[21][4] )
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n1463), .CK(CLK), .Q(\REGISTERS[21][3] )
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n1462), .CK(CLK), .Q(\REGISTERS[21][2] )
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n1461), .CK(CLK), .Q(\REGISTERS[21][1] )
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n1460), .CK(CLK), .Q(\REGISTERS[21][0] )
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n1459), .CK(CLK), .Q(\REGISTERS[22][31] ) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n1458), .CK(CLK), .Q(\REGISTERS[22][30] ) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n1457), .CK(CLK), .Q(\REGISTERS[22][29] ) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n1456), .CK(CLK), .Q(\REGISTERS[22][28] ) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n1455), .CK(CLK), .Q(\REGISTERS[22][27] ) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n1454), .CK(CLK), .Q(\REGISTERS[22][26] ) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n1453), .CK(CLK), .Q(\REGISTERS[22][25] ) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n1452), .CK(CLK), .Q(\REGISTERS[22][24] ) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n1451), .CK(CLK), .Q(\REGISTERS[22][23] ) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n1450), .CK(CLK), .Q(\REGISTERS[22][22] ) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n1449), .CK(CLK), .Q(\REGISTERS[22][21] ) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n1448), .CK(CLK), .Q(\REGISTERS[22][20] ) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n1447), .CK(CLK), .Q(\REGISTERS[22][19] ) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n1446), .CK(CLK), .Q(\REGISTERS[22][18] ) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n1445), .CK(CLK), .Q(\REGISTERS[22][17] ) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n1444), .CK(CLK), .Q(\REGISTERS[22][16] ) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n1443), .CK(CLK), .Q(\REGISTERS[22][15] ) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n1442), .CK(CLK), .Q(\REGISTERS[22][14] ) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n1441), .CK(CLK), .Q(\REGISTERS[22][13] ) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n1440), .CK(CLK), .Q(\REGISTERS[22][12] ) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n1439), .CK(CLK), .Q(\REGISTERS[22][11] ) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n1438), .CK(CLK), .Q(\REGISTERS[22][10] ) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n1437), .CK(CLK), .Q(\REGISTERS[22][9] )
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n1436), .CK(CLK), .Q(\REGISTERS[22][8] )
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n1435), .CK(CLK), .Q(\REGISTERS[22][7] )
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n1434), .CK(CLK), .Q(\REGISTERS[22][6] )
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n1433), .CK(CLK), .Q(\REGISTERS[22][5] )
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n1432), .CK(CLK), .Q(\REGISTERS[22][4] )
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n1431), .CK(CLK), .Q(\REGISTERS[22][3] )
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n1430), .CK(CLK), .Q(\REGISTERS[22][2] )
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n1429), .CK(CLK), .Q(\REGISTERS[22][1] )
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n1428), .CK(CLK), .Q(\REGISTERS[22][0] )
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n1427), .CK(CLK), .Q(\REGISTERS[23][31] ) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n1426), .CK(CLK), .Q(\REGISTERS[23][30] ) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n1425), .CK(CLK), .Q(\REGISTERS[23][29] ) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n1424), .CK(CLK), .Q(\REGISTERS[23][28] ) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n1423), .CK(CLK), .Q(\REGISTERS[23][27] ) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n1422), .CK(CLK), .Q(\REGISTERS[23][26] ) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n1421), .CK(CLK), .Q(\REGISTERS[23][25] ) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n1420), .CK(CLK), .Q(\REGISTERS[23][24] ) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n1419), .CK(CLK), .Q(\REGISTERS[23][23] ) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n1418), .CK(CLK), .Q(\REGISTERS[23][22] ) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n1417), .CK(CLK), .Q(\REGISTERS[23][21] ) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n1416), .CK(CLK), .Q(\REGISTERS[23][20] ) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n1415), .CK(CLK), .Q(\REGISTERS[23][19] ) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n1414), .CK(CLK), .Q(\REGISTERS[23][18] ) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n1413), .CK(CLK), .Q(\REGISTERS[23][17] ) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n1412), .CK(CLK), .Q(\REGISTERS[23][16] ) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n1411), .CK(CLK), .Q(\REGISTERS[23][15] ) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n1410), .CK(CLK), .Q(\REGISTERS[23][14] ) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n1409), .CK(CLK), .Q(\REGISTERS[23][13] ) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n1408), .CK(CLK), .Q(\REGISTERS[23][12] ) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n1407), .CK(CLK), .Q(\REGISTERS[23][11] ) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n1406), .CK(CLK), .Q(\REGISTERS[23][10] ) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n1405), .CK(CLK), .Q(\REGISTERS[23][9] )
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n1404), .CK(CLK), .Q(\REGISTERS[23][8] )
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n1403), .CK(CLK), .Q(\REGISTERS[23][7] )
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n1402), .CK(CLK), .Q(\REGISTERS[23][6] )
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n1401), .CK(CLK), .Q(\REGISTERS[23][5] )
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n1400), .CK(CLK), .Q(\REGISTERS[23][4] )
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n1399), .CK(CLK), .Q(\REGISTERS[23][3] )
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n1398), .CK(CLK), .Q(\REGISTERS[23][2] )
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n1397), .CK(CLK), .Q(\REGISTERS[23][1] )
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n1396), .CK(CLK), .Q(\REGISTERS[23][0] )
         );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n1395), .CK(CLK), .Q(\REGISTERS[24][31] ) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n1394), .CK(CLK), .Q(\REGISTERS[24][30] ) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n1393), .CK(CLK), .Q(\REGISTERS[24][29] ) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n1392), .CK(CLK), .Q(\REGISTERS[24][28] ) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n1391), .CK(CLK), .Q(\REGISTERS[24][27] ) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n1390), .CK(CLK), .Q(\REGISTERS[24][26] ) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n1389), .CK(CLK), .Q(\REGISTERS[24][25] ) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n1388), .CK(CLK), .Q(\REGISTERS[24][24] ) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n1387), .CK(CLK), .Q(\REGISTERS[24][23] ) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n1386), .CK(CLK), .Q(\REGISTERS[24][22] ) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n1385), .CK(CLK), .Q(\REGISTERS[24][21] ) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n1384), .CK(CLK), .Q(\REGISTERS[24][20] ) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n1383), .CK(CLK), .Q(\REGISTERS[24][19] ) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n1382), .CK(CLK), .Q(\REGISTERS[24][18] ) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n1381), .CK(CLK), .Q(\REGISTERS[24][17] ) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n1380), .CK(CLK), .Q(\REGISTERS[24][16] ) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n1379), .CK(CLK), .Q(\REGISTERS[24][15] ) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n1378), .CK(CLK), .Q(\REGISTERS[24][14] ) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n1377), .CK(CLK), .Q(\REGISTERS[24][13] ) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n1376), .CK(CLK), .Q(\REGISTERS[24][12] ) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n1375), .CK(CLK), .Q(\REGISTERS[24][11] ) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n1374), .CK(CLK), .Q(\REGISTERS[24][10] ) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n1373), .CK(CLK), .Q(\REGISTERS[24][9] )
         );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n1372), .CK(CLK), .Q(\REGISTERS[24][8] )
         );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n1371), .CK(CLK), .Q(\REGISTERS[24][7] )
         );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n1370), .CK(CLK), .Q(\REGISTERS[24][6] )
         );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n1369), .CK(CLK), .Q(\REGISTERS[24][5] )
         );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n1368), .CK(CLK), .Q(\REGISTERS[24][4] )
         );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n1367), .CK(CLK), .Q(\REGISTERS[24][3] )
         );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n1366), .CK(CLK), .Q(\REGISTERS[24][2] )
         );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n1365), .CK(CLK), .Q(\REGISTERS[24][1] )
         );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n1364), .CK(CLK), .Q(\REGISTERS[24][0] )
         );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n1363), .CK(CLK), .Q(\REGISTERS[25][31] ) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n1362), .CK(CLK), .Q(\REGISTERS[25][30] ) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n1361), .CK(CLK), .Q(\REGISTERS[25][29] ) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n1360), .CK(CLK), .Q(\REGISTERS[25][28] ) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n1359), .CK(CLK), .Q(\REGISTERS[25][27] ) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n1358), .CK(CLK), .Q(\REGISTERS[25][26] ) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n1357), .CK(CLK), .Q(\REGISTERS[25][25] ) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n1356), .CK(CLK), .Q(\REGISTERS[25][24] ) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n1355), .CK(CLK), .Q(\REGISTERS[25][23] ) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n1354), .CK(CLK), .Q(\REGISTERS[25][22] ) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n1353), .CK(CLK), .Q(\REGISTERS[25][21] ) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n1352), .CK(CLK), .Q(\REGISTERS[25][20] ) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n1351), .CK(CLK), .Q(\REGISTERS[25][19] ) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n1350), .CK(CLK), .Q(\REGISTERS[25][18] ) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n1349), .CK(CLK), .Q(\REGISTERS[25][17] ) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n1348), .CK(CLK), .Q(\REGISTERS[25][16] ) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n1347), .CK(CLK), .Q(\REGISTERS[25][15] ) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n1346), .CK(CLK), .Q(\REGISTERS[25][14] ) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n1345), .CK(CLK), .Q(\REGISTERS[25][13] ) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n1344), .CK(CLK), .Q(\REGISTERS[25][12] ) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n1343), .CK(CLK), .Q(\REGISTERS[25][11] ) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n1342), .CK(CLK), .Q(\REGISTERS[25][10] ) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n1341), .CK(CLK), .Q(\REGISTERS[25][9] )
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n1340), .CK(CLK), .Q(\REGISTERS[25][8] )
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n1339), .CK(CLK), .Q(\REGISTERS[25][7] )
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n1338), .CK(CLK), .Q(\REGISTERS[25][6] )
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n1337), .CK(CLK), .Q(\REGISTERS[25][5] )
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n1336), .CK(CLK), .Q(\REGISTERS[25][4] )
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n1335), .CK(CLK), .Q(\REGISTERS[25][3] )
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n1334), .CK(CLK), .Q(\REGISTERS[25][2] )
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n1333), .CK(CLK), .Q(\REGISTERS[25][1] )
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n1332), .CK(CLK), .Q(\REGISTERS[25][0] )
         );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n1331), .CK(CLK), .Q(\REGISTERS[26][31] ) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n1330), .CK(CLK), .Q(\REGISTERS[26][30] ) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n1329), .CK(CLK), .Q(\REGISTERS[26][29] ) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n1328), .CK(CLK), .Q(\REGISTERS[26][28] ) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n1327), .CK(CLK), .Q(\REGISTERS[26][27] ) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n1326), .CK(CLK), .Q(\REGISTERS[26][26] ) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n1325), .CK(CLK), .Q(\REGISTERS[26][25] ) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n1324), .CK(CLK), .Q(\REGISTERS[26][24] ) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n1323), .CK(CLK), .Q(\REGISTERS[26][23] ) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n1322), .CK(CLK), .Q(\REGISTERS[26][22] ) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n1321), .CK(CLK), .Q(\REGISTERS[26][21] ) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n1320), .CK(CLK), .Q(\REGISTERS[26][20] ) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n1319), .CK(CLK), .Q(\REGISTERS[26][19] ) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n1318), .CK(CLK), .Q(\REGISTERS[26][18] ) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n1317), .CK(CLK), .Q(\REGISTERS[26][17] ) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n1316), .CK(CLK), .Q(\REGISTERS[26][16] ) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n1315), .CK(CLK), .Q(\REGISTERS[26][15] ) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n1314), .CK(CLK), .Q(\REGISTERS[26][14] ) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n1313), .CK(CLK), .Q(\REGISTERS[26][13] ) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n1312), .CK(CLK), .Q(\REGISTERS[26][12] ) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n1311), .CK(CLK), .Q(\REGISTERS[26][11] ) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n1310), .CK(CLK), .Q(\REGISTERS[26][10] ) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n1309), .CK(CLK), .Q(\REGISTERS[26][9] )
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n1308), .CK(CLK), .Q(\REGISTERS[26][8] )
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n1307), .CK(CLK), .Q(\REGISTERS[26][7] )
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n1306), .CK(CLK), .Q(\REGISTERS[26][6] )
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n1305), .CK(CLK), .Q(\REGISTERS[26][5] )
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n1304), .CK(CLK), .Q(\REGISTERS[26][4] )
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n1303), .CK(CLK), .Q(\REGISTERS[26][3] )
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n1302), .CK(CLK), .Q(\REGISTERS[26][2] )
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n1301), .CK(CLK), .Q(\REGISTERS[26][1] )
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n1300), .CK(CLK), .Q(\REGISTERS[26][0] )
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n1299), .CK(CLK), .Q(\REGISTERS[27][31] ) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n1298), .CK(CLK), .Q(\REGISTERS[27][30] ) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n1297), .CK(CLK), .Q(\REGISTERS[27][29] ) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n1296), .CK(CLK), .Q(\REGISTERS[27][28] ) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n1295), .CK(CLK), .Q(\REGISTERS[27][27] ) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n1294), .CK(CLK), .Q(\REGISTERS[27][26] ) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n1293), .CK(CLK), .Q(\REGISTERS[27][25] ) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n1292), .CK(CLK), .Q(\REGISTERS[27][24] ) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n1291), .CK(CLK), .Q(\REGISTERS[27][23] ) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n1290), .CK(CLK), .Q(\REGISTERS[27][22] ) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n1289), .CK(CLK), .Q(\REGISTERS[27][21] ) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n1288), .CK(CLK), .Q(\REGISTERS[27][20] ) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n1287), .CK(CLK), .Q(\REGISTERS[27][19] ) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n1286), .CK(CLK), .Q(\REGISTERS[27][18] ) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n1285), .CK(CLK), .Q(\REGISTERS[27][17] ) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n1284), .CK(CLK), .Q(\REGISTERS[27][16] ) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n1283), .CK(CLK), .Q(\REGISTERS[27][15] ) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n1282), .CK(CLK), .Q(\REGISTERS[27][14] ) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n1281), .CK(CLK), .Q(\REGISTERS[27][13] ) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n1280), .CK(CLK), .Q(\REGISTERS[27][12] ) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n1279), .CK(CLK), .Q(\REGISTERS[27][11] ) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n1278), .CK(CLK), .Q(\REGISTERS[27][10] ) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n1277), .CK(CLK), .Q(\REGISTERS[27][9] )
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n1276), .CK(CLK), .Q(\REGISTERS[27][8] )
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n1275), .CK(CLK), .Q(\REGISTERS[27][7] )
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n1274), .CK(CLK), .Q(\REGISTERS[27][6] )
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n1273), .CK(CLK), .Q(\REGISTERS[27][5] )
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n1272), .CK(CLK), .Q(\REGISTERS[27][4] )
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n1271), .CK(CLK), .Q(\REGISTERS[27][3] )
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n1270), .CK(CLK), .Q(\REGISTERS[27][2] )
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n1269), .CK(CLK), .Q(\REGISTERS[27][1] )
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n1268), .CK(CLK), .Q(\REGISTERS[27][0] )
         );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n1267), .CK(CLK), .Q(\REGISTERS[28][31] ) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n1266), .CK(CLK), .Q(\REGISTERS[28][30] ) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n1265), .CK(CLK), .Q(\REGISTERS[28][29] ) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n1264), .CK(CLK), .Q(\REGISTERS[28][28] ) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n1263), .CK(CLK), .Q(\REGISTERS[28][27] ) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n1262), .CK(CLK), .Q(\REGISTERS[28][26] ) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n1261), .CK(CLK), .Q(\REGISTERS[28][25] ) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n1260), .CK(CLK), .Q(\REGISTERS[28][24] ) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n1259), .CK(CLK), .Q(\REGISTERS[28][23] ) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n1258), .CK(CLK), .Q(\REGISTERS[28][22] ) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n1257), .CK(CLK), .Q(\REGISTERS[28][21] ) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n1256), .CK(CLK), .Q(\REGISTERS[28][20] ) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n1255), .CK(CLK), .Q(\REGISTERS[28][19] ) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n1254), .CK(CLK), .Q(\REGISTERS[28][18] ) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n1253), .CK(CLK), .Q(\REGISTERS[28][17] ) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n1252), .CK(CLK), .Q(\REGISTERS[28][16] ) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n1251), .CK(CLK), .Q(\REGISTERS[28][15] ) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n1250), .CK(CLK), .Q(\REGISTERS[28][14] ) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n1249), .CK(CLK), .Q(\REGISTERS[28][13] ) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n1248), .CK(CLK), .Q(\REGISTERS[28][12] ) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n1247), .CK(CLK), .Q(\REGISTERS[28][11] ) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n1246), .CK(CLK), .Q(\REGISTERS[28][10] ) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n1245), .CK(CLK), .Q(\REGISTERS[28][9] )
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n1244), .CK(CLK), .Q(\REGISTERS[28][8] )
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n1243), .CK(CLK), .Q(\REGISTERS[28][7] )
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n1242), .CK(CLK), .Q(\REGISTERS[28][6] )
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n1241), .CK(CLK), .Q(\REGISTERS[28][5] )
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n1240), .CK(CLK), .Q(\REGISTERS[28][4] )
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n1239), .CK(CLK), .Q(\REGISTERS[28][3] )
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n1238), .CK(CLK), .Q(\REGISTERS[28][2] )
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n1237), .CK(CLK), .Q(\REGISTERS[28][1] )
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n1236), .CK(CLK), .Q(\REGISTERS[28][0] )
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n1235), .CK(CLK), .Q(\REGISTERS[29][31] ) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n1234), .CK(CLK), .Q(\REGISTERS[29][30] ) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n1233), .CK(CLK), .Q(\REGISTERS[29][29] ) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n1232), .CK(CLK), .Q(\REGISTERS[29][28] ) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n1231), .CK(CLK), .Q(\REGISTERS[29][27] ) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n1230), .CK(CLK), .Q(\REGISTERS[29][26] ) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n1229), .CK(CLK), .Q(\REGISTERS[29][25] ) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n1228), .CK(CLK), .Q(\REGISTERS[29][24] ) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n1227), .CK(CLK), .Q(\REGISTERS[29][23] ) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n1226), .CK(CLK), .Q(\REGISTERS[29][22] ) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n1225), .CK(CLK), .Q(\REGISTERS[29][21] ) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n1224), .CK(CLK), .Q(\REGISTERS[29][20] ) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n1223), .CK(CLK), .Q(\REGISTERS[29][19] ) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n1222), .CK(CLK), .Q(\REGISTERS[29][18] ) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n1221), .CK(CLK), .Q(\REGISTERS[29][17] ) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n1220), .CK(CLK), .Q(\REGISTERS[29][16] ) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n1219), .CK(CLK), .Q(\REGISTERS[29][15] ) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n1218), .CK(CLK), .Q(\REGISTERS[29][14] ) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n1217), .CK(CLK), .Q(\REGISTERS[29][13] ) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n1216), .CK(CLK), .Q(\REGISTERS[29][12] ) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n1215), .CK(CLK), .Q(\REGISTERS[29][11] ) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n1214), .CK(CLK), .Q(\REGISTERS[29][10] ) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n1213), .CK(CLK), .Q(\REGISTERS[29][9] )
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n1212), .CK(CLK), .Q(\REGISTERS[29][8] )
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n1211), .CK(CLK), .Q(\REGISTERS[29][7] )
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n1210), .CK(CLK), .Q(\REGISTERS[29][6] )
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n1209), .CK(CLK), .Q(\REGISTERS[29][5] )
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n1208), .CK(CLK), .Q(\REGISTERS[29][4] )
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n1207), .CK(CLK), .Q(\REGISTERS[29][3] )
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n1206), .CK(CLK), .Q(\REGISTERS[29][2] )
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n1205), .CK(CLK), .Q(\REGISTERS[29][1] )
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n1204), .CK(CLK), .Q(\REGISTERS[29][0] )
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n1203), .CK(CLK), .Q(\REGISTERS[30][31] ) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n1202), .CK(CLK), .Q(\REGISTERS[30][30] ) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n1201), .CK(CLK), .Q(\REGISTERS[30][29] ) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n1200), .CK(CLK), .Q(\REGISTERS[30][28] ) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n1199), .CK(CLK), .Q(\REGISTERS[30][27] ) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n1198), .CK(CLK), .Q(\REGISTERS[30][26] ) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n1197), .CK(CLK), .Q(\REGISTERS[30][25] ) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n1196), .CK(CLK), .Q(\REGISTERS[30][24] ) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n1195), .CK(CLK), .Q(\REGISTERS[30][23] ) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n1194), .CK(CLK), .Q(\REGISTERS[30][22] ) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n1193), .CK(CLK), .Q(\REGISTERS[30][21] ) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n1192), .CK(CLK), .Q(\REGISTERS[30][20] ) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n1191), .CK(CLK), .Q(\REGISTERS[30][19] ) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n1190), .CK(CLK), .Q(\REGISTERS[30][18] ) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n1189), .CK(CLK), .Q(\REGISTERS[30][17] ) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n1188), .CK(CLK), .Q(\REGISTERS[30][16] ) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n1187), .CK(CLK), .Q(\REGISTERS[30][15] ) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n1186), .CK(CLK), .Q(\REGISTERS[30][14] ) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n1185), .CK(CLK), .Q(\REGISTERS[30][13] ) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n1184), .CK(CLK), .Q(\REGISTERS[30][12] ) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n1183), .CK(CLK), .Q(\REGISTERS[30][11] ) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n1182), .CK(CLK), .Q(\REGISTERS[30][10] ) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n1181), .CK(CLK), .Q(\REGISTERS[30][9] )
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n1180), .CK(CLK), .Q(\REGISTERS[30][8] )
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n1179), .CK(CLK), .Q(\REGISTERS[30][7] )
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n1178), .CK(CLK), .Q(\REGISTERS[30][6] )
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n1177), .CK(CLK), .Q(\REGISTERS[30][5] )
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n1176), .CK(CLK), .Q(\REGISTERS[30][4] )
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n1175), .CK(CLK), .Q(\REGISTERS[30][3] )
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n1174), .CK(CLK), .Q(\REGISTERS[30][2] )
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n1173), .CK(CLK), .Q(\REGISTERS[30][1] )
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n1172), .CK(CLK), .Q(\REGISTERS[30][0] )
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n1171), .CK(CLK), .Q(\REGISTERS[31][31] ) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n1170), .CK(CLK), .Q(\REGISTERS[31][30] ) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n1169), .CK(CLK), .Q(\REGISTERS[31][29] ) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n1168), .CK(CLK), .Q(\REGISTERS[31][28] ) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n1167), .CK(CLK), .Q(\REGISTERS[31][27] ) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n1166), .CK(CLK), .Q(\REGISTERS[31][26] ) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n1165), .CK(CLK), .Q(\REGISTERS[31][25] ) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n1164), .CK(CLK), .Q(\REGISTERS[31][24] ) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n1163), .CK(CLK), .Q(\REGISTERS[31][23] ) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n1162), .CK(CLK), .Q(\REGISTERS[31][22] ) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n1161), .CK(CLK), .Q(\REGISTERS[31][21] ) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n1160), .CK(CLK), .Q(\REGISTERS[31][20] ) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n1159), .CK(CLK), .Q(\REGISTERS[31][19] ) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n1158), .CK(CLK), .Q(\REGISTERS[31][18] ) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n1157), .CK(CLK), .Q(\REGISTERS[31][17] ) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n1156), .CK(CLK), .Q(\REGISTERS[31][16] ) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n1155), .CK(CLK), .Q(\REGISTERS[31][15] ) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n1154), .CK(CLK), .Q(\REGISTERS[31][14] ) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n1153), .CK(CLK), .Q(\REGISTERS[31][13] ) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n1152), .CK(CLK), .Q(\REGISTERS[31][12] ) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n1151), .CK(CLK), .Q(\REGISTERS[31][11] ) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n1150), .CK(CLK), .Q(\REGISTERS[31][10] ) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n1149), .CK(CLK), .Q(\REGISTERS[31][9] )
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n1148), .CK(CLK), .Q(\REGISTERS[31][8] )
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n1147), .CK(CLK), .Q(\REGISTERS[31][7] )
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n1146), .CK(CLK), .Q(\REGISTERS[31][6] )
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n1145), .CK(CLK), .Q(\REGISTERS[31][5] )
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n1144), .CK(CLK), .Q(\REGISTERS[31][4] )
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n1143), .CK(CLK), .Q(\REGISTERS[31][3] )
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n1142), .CK(CLK), .Q(\REGISTERS[31][2] )
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n1141), .CK(CLK), .Q(\REGISTERS[31][1] )
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n1140), .CK(CLK), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT1_reg[31]  ( .G(N444), .D(N410), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N444), .D(N409), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N444), .D(N408), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N444), .D(N407), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N444), .D(N406), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N444), .D(N405), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N444), .D(N404), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N444), .D(N403), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N444), .D(N402), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N444), .D(N401), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N444), .D(N400), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N444), .D(N399), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N444), .D(N398), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N444), .D(N397), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N444), .D(N396), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N444), .D(N395), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N444), .D(N394), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N444), .D(N393), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N444), .D(N392), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N444), .D(N391), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N444), .D(N390), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N444), .D(N389), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N444), .D(N388), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N444), .D(N387), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N444), .D(N386), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N444), .D(N385), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N444), .D(N384), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N444), .D(N383), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N444), .D(N382), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N444), .D(N381), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N444), .D(N380), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N444), .D(N379), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N445), .D(N443), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N445), .D(N442), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N445), .D(N441), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N445), .D(N440), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N445), .D(N439), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N445), .D(N438), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N445), .D(N437), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N445), .D(N436), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N445), .D(N435), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N445), .D(N434), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N445), .D(N433), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N445), .D(N432), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N445), .D(N431), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N445), .D(N430), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N445), .D(N429), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N445), .D(N428), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N445), .D(N427), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N445), .D(N426), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N445), .D(N425), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N445), .D(N424), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N445), .D(N423), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N445), .D(N422), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N445), .D(N421), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N445), .D(N420), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N445), .D(N419), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N445), .D(N418), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N445), .D(N417), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N445), .D(N416), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N445), .D(N415), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N445), .D(N414), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N445), .D(N413), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N445), .D(N412), .Q(OUT2[0]) );
  INV_X1 U3 ( .A(n3243), .ZN(n1) );
  INV_X2 U4 ( .A(n1), .ZN(n2) );
  INV_X1 U5 ( .A(n3244), .ZN(n3) );
  INV_X2 U6 ( .A(n3), .ZN(n4) );
  INV_X1 U7 ( .A(n3245), .ZN(n5) );
  INV_X2 U8 ( .A(n5), .ZN(n6) );
  INV_X1 U9 ( .A(n3246), .ZN(n7) );
  INV_X2 U10 ( .A(n7), .ZN(n8) );
  INV_X1 U11 ( .A(n3247), .ZN(n9) );
  INV_X2 U12 ( .A(n9), .ZN(n10) );
  INV_X1 U13 ( .A(n3248), .ZN(n11) );
  INV_X2 U14 ( .A(n11), .ZN(n12) );
  INV_X1 U15 ( .A(n3253), .ZN(n13) );
  INV_X2 U16 ( .A(n13), .ZN(n14) );
  INV_X1 U17 ( .A(n3254), .ZN(n15) );
  INV_X2 U18 ( .A(n15), .ZN(n16) );
  INV_X1 U19 ( .A(n3255), .ZN(n17) );
  INV_X2 U20 ( .A(n17), .ZN(n18) );
  INV_X1 U21 ( .A(n3256), .ZN(n19) );
  INV_X2 U22 ( .A(n19), .ZN(n20) );
  INV_X1 U23 ( .A(n3257), .ZN(n21) );
  INV_X2 U24 ( .A(n21), .ZN(n22) );
  INV_X1 U25 ( .A(n3258), .ZN(n23) );
  INV_X2 U26 ( .A(n23), .ZN(n24) );
  INV_X1 U27 ( .A(n3259), .ZN(n25) );
  INV_X2 U28 ( .A(n25), .ZN(n26) );
  INV_X1 U29 ( .A(n3241), .ZN(n27) );
  INV_X2 U30 ( .A(n27), .ZN(n28) );
  INV_X1 U31 ( .A(n3242), .ZN(n29) );
  INV_X2 U32 ( .A(n29), .ZN(n30) );
  INV_X1 U33 ( .A(n3238), .ZN(n31) );
  INV_X2 U34 ( .A(n31), .ZN(n32) );
  INV_X1 U35 ( .A(n3239), .ZN(n33) );
  INV_X2 U36 ( .A(n33), .ZN(n34) );
  INV_X1 U37 ( .A(n3236), .ZN(n35) );
  INV_X2 U38 ( .A(n35), .ZN(n36) );
  INV_X1 U39 ( .A(n3237), .ZN(n37) );
  INV_X2 U40 ( .A(n37), .ZN(n38) );
  INV_X1 U41 ( .A(n3234), .ZN(n39) );
  INV_X2 U42 ( .A(n39), .ZN(n40) );
  INV_X1 U43 ( .A(n3235), .ZN(n41) );
  INV_X2 U44 ( .A(n41), .ZN(n42) );
  INV_X1 U45 ( .A(n3232), .ZN(n43) );
  INV_X2 U46 ( .A(n43), .ZN(n44) );
  INV_X1 U47 ( .A(n3233), .ZN(n45) );
  INV_X2 U48 ( .A(n45), .ZN(n46) );
  INV_X1 U49 ( .A(n3225), .ZN(n47) );
  INV_X2 U50 ( .A(n47), .ZN(n48) );
  INV_X1 U51 ( .A(n3230), .ZN(n49) );
  INV_X2 U52 ( .A(n49), .ZN(n50) );
  INV_X1 U53 ( .A(n3221), .ZN(n51) );
  INV_X2 U54 ( .A(n51), .ZN(n52) );
  INV_X1 U55 ( .A(n3223), .ZN(n53) );
  INV_X2 U56 ( .A(n53), .ZN(n54) );
  INV_X1 U57 ( .A(n3217), .ZN(n55) );
  INV_X2 U58 ( .A(n55), .ZN(n56) );
  INV_X1 U59 ( .A(n3219), .ZN(n57) );
  INV_X2 U60 ( .A(n57), .ZN(n58) );
  INV_X1 U61 ( .A(n3213), .ZN(n59) );
  INV_X2 U62 ( .A(n59), .ZN(n60) );
  INV_X1 U63 ( .A(n3215), .ZN(n61) );
  INV_X2 U64 ( .A(n61), .ZN(n62) );
  OAI21_X4 U65 ( .B1(n3210), .B2(n3211), .A(n3212), .ZN(n3178) );
  INV_X4 U66 ( .A(RESET), .ZN(n3212) );
  BUF_X1 U67 ( .A(ADD_RD1[4]), .Z(n231) );
  BUF_X1 U68 ( .A(ADD_RD1[4]), .Z(n230) );
  BUF_X1 U69 ( .A(ADD_RD1[4]), .Z(n229) );
  BUF_X1 U70 ( .A(ADD_RD1[4]), .Z(n228) );
  BUF_X1 U71 ( .A(ADD_RD1[4]), .Z(n227) );
  BUF_X1 U72 ( .A(ADD_RD1[4]), .Z(n226) );
  BUF_X1 U73 ( .A(ADD_RD1[4]), .Z(n225) );
  BUF_X1 U74 ( .A(ADD_RD1[4]), .Z(n224) );
  BUF_X1 U75 ( .A(ADD_RD2[4]), .Z(n146) );
  BUF_X1 U76 ( .A(ADD_RD2[4]), .Z(n145) );
  BUF_X1 U77 ( .A(ADD_RD2[4]), .Z(n144) );
  BUF_X1 U78 ( .A(ADD_RD2[4]), .Z(n143) );
  BUF_X1 U79 ( .A(ADD_RD2[4]), .Z(n142) );
  BUF_X1 U80 ( .A(ADD_RD2[4]), .Z(n141) );
  BUF_X1 U81 ( .A(ADD_RD2[4]), .Z(n140) );
  BUF_X1 U82 ( .A(ADD_RD2[4]), .Z(n139) );
  BUF_X1 U83 ( .A(ADD_RD1[4]), .Z(n232) );
  BUF_X1 U84 ( .A(ADD_RD2[4]), .Z(n147) );
  CLKBUF_X1 U85 ( .A(ADD_RD2[2]), .Z(n63) );
  CLKBUF_X1 U86 ( .A(ADD_RD2[2]), .Z(n64) );
  CLKBUF_X1 U87 ( .A(ADD_RD2[2]), .Z(n65) );
  CLKBUF_X1 U88 ( .A(ADD_RD2[2]), .Z(n66) );
  CLKBUF_X1 U89 ( .A(ADD_RD2[2]), .Z(n67) );
  CLKBUF_X1 U90 ( .A(ADD_RD2[2]), .Z(n68) );
  CLKBUF_X1 U91 ( .A(ADD_RD2[2]), .Z(n69) );
  CLKBUF_X1 U92 ( .A(ADD_RD2[2]), .Z(n70) );
  CLKBUF_X1 U93 ( .A(ADD_RD2[2]), .Z(n71) );
  CLKBUF_X1 U94 ( .A(ADD_RD2[2]), .Z(n72) );
  CLKBUF_X1 U95 ( .A(ADD_RD2[2]), .Z(n73) );
  CLKBUF_X1 U96 ( .A(ADD_RD2[3]), .Z(n74) );
  CLKBUF_X1 U97 ( .A(ADD_RD2[3]), .Z(n75) );
  CLKBUF_X1 U98 ( .A(ADD_RD2[3]), .Z(n76) );
  CLKBUF_X1 U99 ( .A(ADD_RD2[3]), .Z(n77) );
  CLKBUF_X1 U100 ( .A(ADD_RD2[3]), .Z(n78) );
  CLKBUF_X1 U101 ( .A(ADD_RD2[3]), .Z(n79) );
  CLKBUF_X1 U102 ( .A(ADD_RD2[3]), .Z(n80) );
  CLKBUF_X1 U103 ( .A(ADD_RD2[3]), .Z(n81) );
  CLKBUF_X1 U104 ( .A(ADD_RD2[3]), .Z(n82) );
  CLKBUF_X1 U105 ( .A(ADD_RD2[3]), .Z(n83) );
  CLKBUF_X1 U106 ( .A(ADD_RD2[3]), .Z(n84) );
  CLKBUF_X1 U107 ( .A(ADD_RD2[3]), .Z(n85) );
  CLKBUF_X1 U108 ( .A(ADD_RD2[3]), .Z(n86) );
  CLKBUF_X1 U109 ( .A(ADD_RD2[3]), .Z(n87) );
  CLKBUF_X1 U110 ( .A(ADD_RD2[3]), .Z(n88) );
  CLKBUF_X1 U111 ( .A(ADD_RD2[3]), .Z(n89) );
  CLKBUF_X1 U112 ( .A(ADD_RD2[3]), .Z(n90) );
  CLKBUF_X1 U113 ( .A(ADD_RD2[3]), .Z(n91) );
  CLKBUF_X1 U114 ( .A(ADD_RD2[3]), .Z(n92) );
  CLKBUF_X1 U115 ( .A(ADD_RD2[3]), .Z(n93) );
  CLKBUF_X1 U116 ( .A(ADD_RD2[3]), .Z(n94) );
  CLKBUF_X1 U117 ( .A(ADD_RD2[3]), .Z(n95) );
  CLKBUF_X1 U118 ( .A(n147), .Z(n96) );
  CLKBUF_X1 U119 ( .A(n147), .Z(n97) );
  CLKBUF_X1 U120 ( .A(n147), .Z(n98) );
  CLKBUF_X1 U121 ( .A(n146), .Z(n99) );
  CLKBUF_X1 U122 ( .A(n146), .Z(n100) );
  CLKBUF_X1 U123 ( .A(n146), .Z(n101) );
  CLKBUF_X1 U124 ( .A(n146), .Z(n102) );
  CLKBUF_X1 U125 ( .A(n146), .Z(n103) );
  CLKBUF_X1 U126 ( .A(n145), .Z(n104) );
  CLKBUF_X1 U127 ( .A(n145), .Z(n105) );
  CLKBUF_X1 U128 ( .A(n145), .Z(n106) );
  CLKBUF_X1 U129 ( .A(n145), .Z(n107) );
  CLKBUF_X1 U130 ( .A(n145), .Z(n108) );
  CLKBUF_X1 U131 ( .A(n144), .Z(n109) );
  CLKBUF_X1 U132 ( .A(n144), .Z(n110) );
  CLKBUF_X1 U133 ( .A(n144), .Z(n111) );
  CLKBUF_X1 U134 ( .A(n144), .Z(n112) );
  CLKBUF_X1 U135 ( .A(n144), .Z(n113) );
  CLKBUF_X1 U136 ( .A(n143), .Z(n114) );
  CLKBUF_X1 U137 ( .A(n143), .Z(n115) );
  CLKBUF_X1 U138 ( .A(n143), .Z(n116) );
  CLKBUF_X1 U139 ( .A(n143), .Z(n117) );
  CLKBUF_X1 U140 ( .A(n143), .Z(n118) );
  CLKBUF_X1 U141 ( .A(n142), .Z(n119) );
  CLKBUF_X1 U142 ( .A(n142), .Z(n120) );
  CLKBUF_X1 U143 ( .A(n142), .Z(n121) );
  CLKBUF_X1 U144 ( .A(n142), .Z(n122) );
  CLKBUF_X1 U145 ( .A(n142), .Z(n123) );
  CLKBUF_X1 U146 ( .A(n141), .Z(n124) );
  CLKBUF_X1 U147 ( .A(n141), .Z(n125) );
  CLKBUF_X1 U148 ( .A(n141), .Z(n126) );
  CLKBUF_X1 U149 ( .A(n141), .Z(n127) );
  CLKBUF_X1 U150 ( .A(n141), .Z(n128) );
  CLKBUF_X1 U151 ( .A(n140), .Z(n129) );
  CLKBUF_X1 U152 ( .A(n140), .Z(n130) );
  CLKBUF_X1 U153 ( .A(n140), .Z(n131) );
  CLKBUF_X1 U154 ( .A(n140), .Z(n132) );
  CLKBUF_X1 U155 ( .A(n140), .Z(n133) );
  CLKBUF_X1 U156 ( .A(n139), .Z(n134) );
  CLKBUF_X1 U157 ( .A(n139), .Z(n135) );
  CLKBUF_X1 U158 ( .A(n139), .Z(n136) );
  CLKBUF_X1 U159 ( .A(n139), .Z(n137) );
  CLKBUF_X1 U160 ( .A(n139), .Z(n138) );
  CLKBUF_X1 U161 ( .A(ADD_RD1[2]), .Z(n148) );
  CLKBUF_X1 U162 ( .A(ADD_RD1[2]), .Z(n149) );
  CLKBUF_X1 U163 ( .A(ADD_RD1[2]), .Z(n150) );
  CLKBUF_X1 U164 ( .A(ADD_RD1[2]), .Z(n151) );
  CLKBUF_X1 U165 ( .A(ADD_RD1[2]), .Z(n152) );
  CLKBUF_X1 U166 ( .A(ADD_RD1[2]), .Z(n153) );
  CLKBUF_X1 U167 ( .A(ADD_RD1[2]), .Z(n154) );
  CLKBUF_X1 U168 ( .A(ADD_RD1[2]), .Z(n155) );
  CLKBUF_X1 U169 ( .A(ADD_RD1[2]), .Z(n156) );
  CLKBUF_X1 U170 ( .A(ADD_RD1[2]), .Z(n157) );
  CLKBUF_X1 U171 ( .A(ADD_RD1[2]), .Z(n158) );
  CLKBUF_X1 U172 ( .A(ADD_RD1[3]), .Z(n159) );
  CLKBUF_X1 U173 ( .A(ADD_RD1[3]), .Z(n160) );
  CLKBUF_X1 U174 ( .A(ADD_RD1[3]), .Z(n161) );
  CLKBUF_X1 U175 ( .A(ADD_RD1[3]), .Z(n162) );
  CLKBUF_X1 U176 ( .A(ADD_RD1[3]), .Z(n163) );
  CLKBUF_X1 U177 ( .A(ADD_RD1[3]), .Z(n164) );
  CLKBUF_X1 U178 ( .A(ADD_RD1[3]), .Z(n165) );
  CLKBUF_X1 U179 ( .A(ADD_RD1[3]), .Z(n166) );
  CLKBUF_X1 U180 ( .A(ADD_RD1[3]), .Z(n167) );
  CLKBUF_X1 U181 ( .A(ADD_RD1[3]), .Z(n168) );
  CLKBUF_X1 U182 ( .A(ADD_RD1[3]), .Z(n169) );
  CLKBUF_X1 U183 ( .A(ADD_RD1[3]), .Z(n170) );
  CLKBUF_X1 U184 ( .A(ADD_RD1[3]), .Z(n171) );
  CLKBUF_X1 U185 ( .A(ADD_RD1[3]), .Z(n172) );
  CLKBUF_X1 U186 ( .A(ADD_RD1[3]), .Z(n173) );
  CLKBUF_X1 U187 ( .A(ADD_RD1[3]), .Z(n174) );
  CLKBUF_X1 U188 ( .A(ADD_RD1[3]), .Z(n175) );
  CLKBUF_X1 U189 ( .A(ADD_RD1[3]), .Z(n176) );
  CLKBUF_X1 U190 ( .A(ADD_RD1[3]), .Z(n177) );
  CLKBUF_X1 U191 ( .A(ADD_RD1[3]), .Z(n178) );
  CLKBUF_X1 U192 ( .A(ADD_RD1[3]), .Z(n179) );
  CLKBUF_X1 U193 ( .A(ADD_RD1[3]), .Z(n180) );
  CLKBUF_X1 U194 ( .A(n232), .Z(n181) );
  CLKBUF_X1 U195 ( .A(n232), .Z(n182) );
  CLKBUF_X1 U196 ( .A(n232), .Z(n183) );
  CLKBUF_X1 U197 ( .A(n231), .Z(n184) );
  CLKBUF_X1 U198 ( .A(n231), .Z(n185) );
  CLKBUF_X1 U199 ( .A(n231), .Z(n186) );
  CLKBUF_X1 U200 ( .A(n231), .Z(n187) );
  CLKBUF_X1 U201 ( .A(n231), .Z(n188) );
  CLKBUF_X1 U202 ( .A(n230), .Z(n189) );
  CLKBUF_X1 U203 ( .A(n230), .Z(n190) );
  CLKBUF_X1 U204 ( .A(n230), .Z(n191) );
  CLKBUF_X1 U205 ( .A(n230), .Z(n192) );
  CLKBUF_X1 U206 ( .A(n230), .Z(n193) );
  CLKBUF_X1 U207 ( .A(n229), .Z(n194) );
  CLKBUF_X1 U208 ( .A(n229), .Z(n195) );
  CLKBUF_X1 U209 ( .A(n229), .Z(n196) );
  CLKBUF_X1 U210 ( .A(n229), .Z(n197) );
  CLKBUF_X1 U211 ( .A(n229), .Z(n198) );
  CLKBUF_X1 U212 ( .A(n228), .Z(n199) );
  CLKBUF_X1 U213 ( .A(n228), .Z(n200) );
  CLKBUF_X1 U214 ( .A(n228), .Z(n201) );
  CLKBUF_X1 U215 ( .A(n228), .Z(n202) );
  CLKBUF_X1 U216 ( .A(n228), .Z(n203) );
  CLKBUF_X1 U217 ( .A(n227), .Z(n204) );
  CLKBUF_X1 U218 ( .A(n227), .Z(n205) );
  CLKBUF_X1 U219 ( .A(n227), .Z(n206) );
  CLKBUF_X1 U220 ( .A(n227), .Z(n207) );
  CLKBUF_X1 U221 ( .A(n227), .Z(n208) );
  CLKBUF_X1 U222 ( .A(n226), .Z(n209) );
  CLKBUF_X1 U223 ( .A(n226), .Z(n210) );
  CLKBUF_X1 U224 ( .A(n226), .Z(n211) );
  CLKBUF_X1 U225 ( .A(n226), .Z(n212) );
  CLKBUF_X1 U226 ( .A(n226), .Z(n213) );
  CLKBUF_X1 U227 ( .A(n225), .Z(n214) );
  CLKBUF_X1 U228 ( .A(n225), .Z(n215) );
  CLKBUF_X1 U229 ( .A(n225), .Z(n216) );
  CLKBUF_X1 U230 ( .A(n225), .Z(n217) );
  CLKBUF_X1 U231 ( .A(n225), .Z(n218) );
  CLKBUF_X1 U232 ( .A(n224), .Z(n219) );
  CLKBUF_X1 U233 ( .A(n224), .Z(n220) );
  CLKBUF_X1 U234 ( .A(n224), .Z(n221) );
  CLKBUF_X1 U235 ( .A(n224), .Z(n222) );
  CLKBUF_X1 U236 ( .A(n224), .Z(n223) );
  MUX2_X1 U237 ( .A(\REGISTERS[15][0] ), .B(\REGISTERS[31][0] ), .S(n96), .Z(
        n233) );
  MUX2_X1 U238 ( .A(\REGISTERS[7][0] ), .B(\REGISTERS[23][0] ), .S(n96), .Z(
        n234) );
  MUX2_X1 U239 ( .A(n234), .B(n233), .S(n74), .Z(n235) );
  MUX2_X1 U240 ( .A(\REGISTERS[11][0] ), .B(\REGISTERS[27][0] ), .S(n96), .Z(
        n236) );
  MUX2_X1 U241 ( .A(\REGISTERS[3][0] ), .B(\REGISTERS[19][0] ), .S(n96), .Z(
        n237) );
  MUX2_X1 U242 ( .A(n237), .B(n236), .S(n74), .Z(n238) );
  MUX2_X1 U243 ( .A(n238), .B(n235), .S(n63), .Z(n239) );
  MUX2_X1 U244 ( .A(\REGISTERS[14][0] ), .B(\REGISTERS[30][0] ), .S(n96), .Z(
        n240) );
  MUX2_X1 U245 ( .A(\REGISTERS[6][0] ), .B(\REGISTERS[22][0] ), .S(n96), .Z(
        n241) );
  MUX2_X1 U246 ( .A(n241), .B(n240), .S(n74), .Z(n242) );
  MUX2_X1 U247 ( .A(\REGISTERS[10][0] ), .B(\REGISTERS[26][0] ), .S(n96), .Z(
        n243) );
  MUX2_X1 U248 ( .A(\REGISTERS[2][0] ), .B(\REGISTERS[18][0] ), .S(n96), .Z(
        n244) );
  MUX2_X1 U249 ( .A(n244), .B(n243), .S(n74), .Z(n245) );
  MUX2_X1 U250 ( .A(n245), .B(n242), .S(n63), .Z(n246) );
  MUX2_X1 U251 ( .A(n246), .B(n239), .S(ADD_RD2[0]), .Z(n247) );
  MUX2_X1 U252 ( .A(\REGISTERS[13][0] ), .B(\REGISTERS[29][0] ), .S(n96), .Z(
        n248) );
  MUX2_X1 U253 ( .A(\REGISTERS[5][0] ), .B(\REGISTERS[21][0] ), .S(n96), .Z(
        n249) );
  MUX2_X1 U254 ( .A(n249), .B(n248), .S(n74), .Z(n250) );
  MUX2_X1 U255 ( .A(\REGISTERS[9][0] ), .B(\REGISTERS[25][0] ), .S(n96), .Z(
        n251) );
  MUX2_X1 U256 ( .A(\REGISTERS[1][0] ), .B(\REGISTERS[17][0] ), .S(n96), .Z(
        n252) );
  MUX2_X1 U257 ( .A(n252), .B(n251), .S(n74), .Z(n253) );
  MUX2_X1 U258 ( .A(n253), .B(n250), .S(n63), .Z(n254) );
  MUX2_X1 U259 ( .A(\REGISTERS[12][0] ), .B(\REGISTERS[28][0] ), .S(n97), .Z(
        n255) );
  MUX2_X1 U260 ( .A(\REGISTERS[4][0] ), .B(\REGISTERS[20][0] ), .S(n97), .Z(
        n256) );
  MUX2_X1 U261 ( .A(n256), .B(n255), .S(n74), .Z(n257) );
  MUX2_X1 U262 ( .A(\REGISTERS[8][0] ), .B(\REGISTERS[24][0] ), .S(n97), .Z(
        n258) );
  MUX2_X1 U263 ( .A(\REGISTERS[0][0] ), .B(\REGISTERS[16][0] ), .S(n97), .Z(
        n259) );
  MUX2_X1 U264 ( .A(n259), .B(n258), .S(n74), .Z(n260) );
  MUX2_X1 U265 ( .A(n260), .B(n257), .S(n63), .Z(n261) );
  MUX2_X1 U266 ( .A(n261), .B(n254), .S(ADD_RD2[0]), .Z(n262) );
  MUX2_X1 U267 ( .A(n262), .B(n247), .S(ADD_RD2[1]), .Z(N412) );
  MUX2_X1 U268 ( .A(\REGISTERS[15][1] ), .B(\REGISTERS[31][1] ), .S(n97), .Z(
        n263) );
  MUX2_X1 U269 ( .A(\REGISTERS[7][1] ), .B(\REGISTERS[23][1] ), .S(n97), .Z(
        n264) );
  MUX2_X1 U270 ( .A(n264), .B(n263), .S(n74), .Z(n265) );
  MUX2_X1 U271 ( .A(\REGISTERS[11][1] ), .B(\REGISTERS[27][1] ), .S(n97), .Z(
        n266) );
  MUX2_X1 U272 ( .A(\REGISTERS[3][1] ), .B(\REGISTERS[19][1] ), .S(n97), .Z(
        n267) );
  MUX2_X1 U273 ( .A(n267), .B(n266), .S(n74), .Z(n268) );
  MUX2_X1 U274 ( .A(n268), .B(n265), .S(n63), .Z(n269) );
  MUX2_X1 U275 ( .A(\REGISTERS[14][1] ), .B(\REGISTERS[30][1] ), .S(n97), .Z(
        n270) );
  MUX2_X1 U276 ( .A(\REGISTERS[6][1] ), .B(\REGISTERS[22][1] ), .S(n97), .Z(
        n271) );
  MUX2_X1 U277 ( .A(n271), .B(n270), .S(n74), .Z(n272) );
  MUX2_X1 U278 ( .A(\REGISTERS[10][1] ), .B(\REGISTERS[26][1] ), .S(n97), .Z(
        n273) );
  MUX2_X1 U279 ( .A(\REGISTERS[2][1] ), .B(\REGISTERS[18][1] ), .S(n97), .Z(
        n274) );
  MUX2_X1 U280 ( .A(n274), .B(n273), .S(n74), .Z(n275) );
  MUX2_X1 U281 ( .A(n275), .B(n272), .S(n63), .Z(n276) );
  MUX2_X1 U282 ( .A(n276), .B(n269), .S(ADD_RD2[0]), .Z(n277) );
  MUX2_X1 U283 ( .A(\REGISTERS[13][1] ), .B(\REGISTERS[29][1] ), .S(n98), .Z(
        n278) );
  MUX2_X1 U284 ( .A(\REGISTERS[5][1] ), .B(\REGISTERS[21][1] ), .S(n98), .Z(
        n279) );
  MUX2_X1 U285 ( .A(n279), .B(n278), .S(n75), .Z(n280) );
  MUX2_X1 U286 ( .A(\REGISTERS[9][1] ), .B(\REGISTERS[25][1] ), .S(n98), .Z(
        n281) );
  MUX2_X1 U287 ( .A(\REGISTERS[1][1] ), .B(\REGISTERS[17][1] ), .S(n98), .Z(
        n282) );
  MUX2_X1 U288 ( .A(n282), .B(n281), .S(n75), .Z(n283) );
  MUX2_X1 U289 ( .A(n283), .B(n280), .S(n63), .Z(n284) );
  MUX2_X1 U290 ( .A(\REGISTERS[12][1] ), .B(\REGISTERS[28][1] ), .S(n98), .Z(
        n285) );
  MUX2_X1 U291 ( .A(\REGISTERS[4][1] ), .B(\REGISTERS[20][1] ), .S(n98), .Z(
        n286) );
  MUX2_X1 U292 ( .A(n286), .B(n285), .S(n75), .Z(n287) );
  MUX2_X1 U293 ( .A(\REGISTERS[8][1] ), .B(\REGISTERS[24][1] ), .S(n98), .Z(
        n288) );
  MUX2_X1 U294 ( .A(\REGISTERS[0][1] ), .B(\REGISTERS[16][1] ), .S(n98), .Z(
        n289) );
  MUX2_X1 U295 ( .A(n289), .B(n288), .S(n75), .Z(n290) );
  MUX2_X1 U296 ( .A(n290), .B(n287), .S(n63), .Z(n291) );
  MUX2_X1 U297 ( .A(n291), .B(n284), .S(ADD_RD2[0]), .Z(n292) );
  MUX2_X1 U298 ( .A(n292), .B(n277), .S(ADD_RD2[1]), .Z(N413) );
  MUX2_X1 U299 ( .A(\REGISTERS[15][2] ), .B(\REGISTERS[31][2] ), .S(n98), .Z(
        n293) );
  MUX2_X1 U300 ( .A(\REGISTERS[7][2] ), .B(\REGISTERS[23][2] ), .S(n98), .Z(
        n294) );
  MUX2_X1 U301 ( .A(n294), .B(n293), .S(n75), .Z(n295) );
  MUX2_X1 U302 ( .A(\REGISTERS[11][2] ), .B(\REGISTERS[27][2] ), .S(n98), .Z(
        n296) );
  MUX2_X1 U303 ( .A(\REGISTERS[3][2] ), .B(\REGISTERS[19][2] ), .S(n98), .Z(
        n297) );
  MUX2_X1 U304 ( .A(n297), .B(n296), .S(n75), .Z(n298) );
  MUX2_X1 U305 ( .A(n298), .B(n295), .S(n63), .Z(n299) );
  MUX2_X1 U306 ( .A(\REGISTERS[14][2] ), .B(\REGISTERS[30][2] ), .S(n99), .Z(
        n300) );
  MUX2_X1 U307 ( .A(\REGISTERS[6][2] ), .B(\REGISTERS[22][2] ), .S(n99), .Z(
        n301) );
  MUX2_X1 U308 ( .A(n301), .B(n300), .S(n75), .Z(n302) );
  MUX2_X1 U309 ( .A(\REGISTERS[10][2] ), .B(\REGISTERS[26][2] ), .S(n99), .Z(
        n303) );
  MUX2_X1 U310 ( .A(\REGISTERS[2][2] ), .B(\REGISTERS[18][2] ), .S(n99), .Z(
        n304) );
  MUX2_X1 U311 ( .A(n304), .B(n303), .S(n75), .Z(n305) );
  MUX2_X1 U312 ( .A(n305), .B(n302), .S(n63), .Z(n306) );
  MUX2_X1 U313 ( .A(n306), .B(n299), .S(ADD_RD2[0]), .Z(n307) );
  MUX2_X1 U314 ( .A(\REGISTERS[13][2] ), .B(\REGISTERS[29][2] ), .S(n99), .Z(
        n308) );
  MUX2_X1 U315 ( .A(\REGISTERS[5][2] ), .B(\REGISTERS[21][2] ), .S(n99), .Z(
        n309) );
  MUX2_X1 U316 ( .A(n309), .B(n308), .S(n75), .Z(n310) );
  MUX2_X1 U317 ( .A(\REGISTERS[9][2] ), .B(\REGISTERS[25][2] ), .S(n99), .Z(
        n311) );
  MUX2_X1 U318 ( .A(\REGISTERS[1][2] ), .B(\REGISTERS[17][2] ), .S(n99), .Z(
        n312) );
  MUX2_X1 U319 ( .A(n312), .B(n311), .S(n75), .Z(n313) );
  MUX2_X1 U320 ( .A(n313), .B(n310), .S(n63), .Z(n314) );
  MUX2_X1 U321 ( .A(\REGISTERS[12][2] ), .B(\REGISTERS[28][2] ), .S(n99), .Z(
        n315) );
  MUX2_X1 U322 ( .A(\REGISTERS[4][2] ), .B(\REGISTERS[20][2] ), .S(n99), .Z(
        n316) );
  MUX2_X1 U323 ( .A(n316), .B(n315), .S(n75), .Z(n317) );
  MUX2_X1 U324 ( .A(\REGISTERS[8][2] ), .B(\REGISTERS[24][2] ), .S(n99), .Z(
        n318) );
  MUX2_X1 U325 ( .A(\REGISTERS[0][2] ), .B(\REGISTERS[16][2] ), .S(n99), .Z(
        n319) );
  MUX2_X1 U326 ( .A(n319), .B(n318), .S(n75), .Z(n320) );
  MUX2_X1 U327 ( .A(n320), .B(n317), .S(n63), .Z(n321) );
  MUX2_X1 U328 ( .A(n321), .B(n314), .S(ADD_RD2[0]), .Z(n322) );
  MUX2_X1 U329 ( .A(n322), .B(n307), .S(ADD_RD2[1]), .Z(N414) );
  MUX2_X1 U330 ( .A(\REGISTERS[15][3] ), .B(\REGISTERS[31][3] ), .S(n100), .Z(
        n323) );
  MUX2_X1 U331 ( .A(\REGISTERS[7][3] ), .B(\REGISTERS[23][3] ), .S(n100), .Z(
        n324) );
  MUX2_X1 U332 ( .A(n324), .B(n323), .S(n76), .Z(n325) );
  MUX2_X1 U333 ( .A(\REGISTERS[11][3] ), .B(\REGISTERS[27][3] ), .S(n100), .Z(
        n326) );
  MUX2_X1 U334 ( .A(\REGISTERS[3][3] ), .B(\REGISTERS[19][3] ), .S(n100), .Z(
        n327) );
  MUX2_X1 U335 ( .A(n327), .B(n326), .S(n76), .Z(n328) );
  MUX2_X1 U336 ( .A(n328), .B(n325), .S(n64), .Z(n329) );
  MUX2_X1 U337 ( .A(\REGISTERS[14][3] ), .B(\REGISTERS[30][3] ), .S(n100), .Z(
        n330) );
  MUX2_X1 U338 ( .A(\REGISTERS[6][3] ), .B(\REGISTERS[22][3] ), .S(n100), .Z(
        n331) );
  MUX2_X1 U339 ( .A(n331), .B(n330), .S(n76), .Z(n332) );
  MUX2_X1 U340 ( .A(\REGISTERS[10][3] ), .B(\REGISTERS[26][3] ), .S(n100), .Z(
        n333) );
  MUX2_X1 U341 ( .A(\REGISTERS[2][3] ), .B(\REGISTERS[18][3] ), .S(n100), .Z(
        n334) );
  MUX2_X1 U342 ( .A(n334), .B(n333), .S(n76), .Z(n335) );
  MUX2_X1 U343 ( .A(n335), .B(n332), .S(n64), .Z(n336) );
  MUX2_X1 U344 ( .A(n336), .B(n329), .S(ADD_RD2[0]), .Z(n337) );
  MUX2_X1 U345 ( .A(\REGISTERS[13][3] ), .B(\REGISTERS[29][3] ), .S(n100), .Z(
        n338) );
  MUX2_X1 U346 ( .A(\REGISTERS[5][3] ), .B(\REGISTERS[21][3] ), .S(n100), .Z(
        n339) );
  MUX2_X1 U347 ( .A(n339), .B(n338), .S(n76), .Z(n340) );
  MUX2_X1 U348 ( .A(\REGISTERS[9][3] ), .B(\REGISTERS[25][3] ), .S(n100), .Z(
        n341) );
  MUX2_X1 U349 ( .A(\REGISTERS[1][3] ), .B(\REGISTERS[17][3] ), .S(n100), .Z(
        n342) );
  MUX2_X1 U350 ( .A(n342), .B(n341), .S(n76), .Z(n343) );
  MUX2_X1 U351 ( .A(n343), .B(n340), .S(n64), .Z(n344) );
  MUX2_X1 U352 ( .A(\REGISTERS[12][3] ), .B(\REGISTERS[28][3] ), .S(n101), .Z(
        n345) );
  MUX2_X1 U353 ( .A(\REGISTERS[4][3] ), .B(\REGISTERS[20][3] ), .S(n101), .Z(
        n346) );
  MUX2_X1 U354 ( .A(n346), .B(n345), .S(n76), .Z(n347) );
  MUX2_X1 U355 ( .A(\REGISTERS[8][3] ), .B(\REGISTERS[24][3] ), .S(n101), .Z(
        n348) );
  MUX2_X1 U356 ( .A(\REGISTERS[0][3] ), .B(\REGISTERS[16][3] ), .S(n101), .Z(
        n349) );
  MUX2_X1 U357 ( .A(n349), .B(n348), .S(n76), .Z(n350) );
  MUX2_X1 U358 ( .A(n350), .B(n347), .S(n64), .Z(n351) );
  MUX2_X1 U359 ( .A(n351), .B(n344), .S(ADD_RD2[0]), .Z(n352) );
  MUX2_X1 U360 ( .A(n352), .B(n337), .S(ADD_RD2[1]), .Z(N415) );
  MUX2_X1 U361 ( .A(\REGISTERS[15][4] ), .B(\REGISTERS[31][4] ), .S(n101), .Z(
        n353) );
  MUX2_X1 U362 ( .A(\REGISTERS[7][4] ), .B(\REGISTERS[23][4] ), .S(n101), .Z(
        n354) );
  MUX2_X1 U363 ( .A(n354), .B(n353), .S(n76), .Z(n355) );
  MUX2_X1 U364 ( .A(\REGISTERS[11][4] ), .B(\REGISTERS[27][4] ), .S(n101), .Z(
        n356) );
  MUX2_X1 U365 ( .A(\REGISTERS[3][4] ), .B(\REGISTERS[19][4] ), .S(n101), .Z(
        n357) );
  MUX2_X1 U366 ( .A(n357), .B(n356), .S(n76), .Z(n358) );
  MUX2_X1 U367 ( .A(n358), .B(n355), .S(n64), .Z(n359) );
  MUX2_X1 U368 ( .A(\REGISTERS[14][4] ), .B(\REGISTERS[30][4] ), .S(n101), .Z(
        n360) );
  MUX2_X1 U369 ( .A(\REGISTERS[6][4] ), .B(\REGISTERS[22][4] ), .S(n101), .Z(
        n361) );
  MUX2_X1 U370 ( .A(n361), .B(n360), .S(n76), .Z(n362) );
  MUX2_X1 U371 ( .A(\REGISTERS[10][4] ), .B(\REGISTERS[26][4] ), .S(n101), .Z(
        n363) );
  MUX2_X1 U372 ( .A(\REGISTERS[2][4] ), .B(\REGISTERS[18][4] ), .S(n101), .Z(
        n364) );
  MUX2_X1 U373 ( .A(n364), .B(n363), .S(n76), .Z(n365) );
  MUX2_X1 U374 ( .A(n365), .B(n362), .S(n64), .Z(n366) );
  MUX2_X1 U375 ( .A(n366), .B(n359), .S(ADD_RD2[0]), .Z(n367) );
  MUX2_X1 U376 ( .A(\REGISTERS[13][4] ), .B(\REGISTERS[29][4] ), .S(n102), .Z(
        n368) );
  MUX2_X1 U377 ( .A(\REGISTERS[5][4] ), .B(\REGISTERS[21][4] ), .S(n102), .Z(
        n369) );
  MUX2_X1 U378 ( .A(n369), .B(n368), .S(n77), .Z(n370) );
  MUX2_X1 U379 ( .A(\REGISTERS[9][4] ), .B(\REGISTERS[25][4] ), .S(n102), .Z(
        n371) );
  MUX2_X1 U380 ( .A(\REGISTERS[1][4] ), .B(\REGISTERS[17][4] ), .S(n102), .Z(
        n372) );
  MUX2_X1 U381 ( .A(n372), .B(n371), .S(n77), .Z(n373) );
  MUX2_X1 U382 ( .A(n373), .B(n370), .S(n64), .Z(n374) );
  MUX2_X1 U383 ( .A(\REGISTERS[12][4] ), .B(\REGISTERS[28][4] ), .S(n102), .Z(
        n375) );
  MUX2_X1 U384 ( .A(\REGISTERS[4][4] ), .B(\REGISTERS[20][4] ), .S(n102), .Z(
        n376) );
  MUX2_X1 U385 ( .A(n376), .B(n375), .S(n77), .Z(n377) );
  MUX2_X1 U386 ( .A(\REGISTERS[8][4] ), .B(\REGISTERS[24][4] ), .S(n102), .Z(
        n378) );
  MUX2_X1 U387 ( .A(\REGISTERS[0][4] ), .B(\REGISTERS[16][4] ), .S(n102), .Z(
        n379) );
  MUX2_X1 U388 ( .A(n379), .B(n378), .S(n77), .Z(n380) );
  MUX2_X1 U389 ( .A(n380), .B(n377), .S(n64), .Z(n381) );
  MUX2_X1 U390 ( .A(n381), .B(n374), .S(ADD_RD2[0]), .Z(n382) );
  MUX2_X1 U391 ( .A(n382), .B(n367), .S(ADD_RD2[1]), .Z(N416) );
  MUX2_X1 U392 ( .A(\REGISTERS[15][5] ), .B(\REGISTERS[31][5] ), .S(n102), .Z(
        n383) );
  MUX2_X1 U393 ( .A(\REGISTERS[7][5] ), .B(\REGISTERS[23][5] ), .S(n102), .Z(
        n384) );
  MUX2_X1 U394 ( .A(n384), .B(n383), .S(n77), .Z(n385) );
  MUX2_X1 U395 ( .A(\REGISTERS[11][5] ), .B(\REGISTERS[27][5] ), .S(n102), .Z(
        n386) );
  MUX2_X1 U396 ( .A(\REGISTERS[3][5] ), .B(\REGISTERS[19][5] ), .S(n102), .Z(
        n387) );
  MUX2_X1 U397 ( .A(n387), .B(n386), .S(n77), .Z(n388) );
  MUX2_X1 U398 ( .A(n388), .B(n385), .S(n64), .Z(n389) );
  MUX2_X1 U399 ( .A(\REGISTERS[14][5] ), .B(\REGISTERS[30][5] ), .S(n103), .Z(
        n390) );
  MUX2_X1 U400 ( .A(\REGISTERS[6][5] ), .B(\REGISTERS[22][5] ), .S(n103), .Z(
        n391) );
  MUX2_X1 U401 ( .A(n391), .B(n390), .S(n77), .Z(n392) );
  MUX2_X1 U402 ( .A(\REGISTERS[10][5] ), .B(\REGISTERS[26][5] ), .S(n103), .Z(
        n393) );
  MUX2_X1 U403 ( .A(\REGISTERS[2][5] ), .B(\REGISTERS[18][5] ), .S(n103), .Z(
        n394) );
  MUX2_X1 U404 ( .A(n394), .B(n393), .S(n77), .Z(n395) );
  MUX2_X1 U405 ( .A(n395), .B(n392), .S(n64), .Z(n396) );
  MUX2_X1 U406 ( .A(n396), .B(n389), .S(ADD_RD2[0]), .Z(n397) );
  MUX2_X1 U407 ( .A(\REGISTERS[13][5] ), .B(\REGISTERS[29][5] ), .S(n103), .Z(
        n398) );
  MUX2_X1 U408 ( .A(\REGISTERS[5][5] ), .B(\REGISTERS[21][5] ), .S(n103), .Z(
        n399) );
  MUX2_X1 U409 ( .A(n399), .B(n398), .S(n77), .Z(n400) );
  MUX2_X1 U410 ( .A(\REGISTERS[9][5] ), .B(\REGISTERS[25][5] ), .S(n103), .Z(
        n401) );
  MUX2_X1 U411 ( .A(\REGISTERS[1][5] ), .B(\REGISTERS[17][5] ), .S(n103), .Z(
        n402) );
  MUX2_X1 U412 ( .A(n402), .B(n401), .S(n77), .Z(n403) );
  MUX2_X1 U413 ( .A(n403), .B(n400), .S(n64), .Z(n404) );
  MUX2_X1 U414 ( .A(\REGISTERS[12][5] ), .B(\REGISTERS[28][5] ), .S(n103), .Z(
        n405) );
  MUX2_X1 U415 ( .A(\REGISTERS[4][5] ), .B(\REGISTERS[20][5] ), .S(n103), .Z(
        n406) );
  MUX2_X1 U416 ( .A(n406), .B(n405), .S(n77), .Z(n407) );
  MUX2_X1 U417 ( .A(\REGISTERS[8][5] ), .B(\REGISTERS[24][5] ), .S(n103), .Z(
        n408) );
  MUX2_X1 U418 ( .A(\REGISTERS[0][5] ), .B(\REGISTERS[16][5] ), .S(n103), .Z(
        n409) );
  MUX2_X1 U419 ( .A(n409), .B(n408), .S(n77), .Z(n410) );
  MUX2_X1 U420 ( .A(n410), .B(n407), .S(n64), .Z(n411) );
  MUX2_X1 U421 ( .A(n411), .B(n404), .S(ADD_RD2[0]), .Z(n412) );
  MUX2_X1 U422 ( .A(n412), .B(n397), .S(ADD_RD2[1]), .Z(N417) );
  MUX2_X1 U423 ( .A(\REGISTERS[15][6] ), .B(\REGISTERS[31][6] ), .S(n104), .Z(
        n413) );
  MUX2_X1 U424 ( .A(\REGISTERS[7][6] ), .B(\REGISTERS[23][6] ), .S(n104), .Z(
        n414) );
  MUX2_X1 U425 ( .A(n414), .B(n413), .S(n78), .Z(n415) );
  MUX2_X1 U426 ( .A(\REGISTERS[11][6] ), .B(\REGISTERS[27][6] ), .S(n104), .Z(
        n416) );
  MUX2_X1 U427 ( .A(\REGISTERS[3][6] ), .B(\REGISTERS[19][6] ), .S(n104), .Z(
        n417) );
  MUX2_X1 U428 ( .A(n417), .B(n416), .S(n78), .Z(n418) );
  MUX2_X1 U429 ( .A(n418), .B(n415), .S(n65), .Z(n419) );
  MUX2_X1 U430 ( .A(\REGISTERS[14][6] ), .B(\REGISTERS[30][6] ), .S(n104), .Z(
        n420) );
  MUX2_X1 U431 ( .A(\REGISTERS[6][6] ), .B(\REGISTERS[22][6] ), .S(n104), .Z(
        n421) );
  MUX2_X1 U432 ( .A(n421), .B(n420), .S(n78), .Z(n422) );
  MUX2_X1 U433 ( .A(\REGISTERS[10][6] ), .B(\REGISTERS[26][6] ), .S(n104), .Z(
        n423) );
  MUX2_X1 U434 ( .A(\REGISTERS[2][6] ), .B(\REGISTERS[18][6] ), .S(n104), .Z(
        n424) );
  MUX2_X1 U435 ( .A(n424), .B(n423), .S(n78), .Z(n425) );
  MUX2_X1 U436 ( .A(n425), .B(n422), .S(n65), .Z(n426) );
  MUX2_X1 U437 ( .A(n426), .B(n419), .S(ADD_RD2[0]), .Z(n427) );
  MUX2_X1 U438 ( .A(\REGISTERS[13][6] ), .B(\REGISTERS[29][6] ), .S(n104), .Z(
        n428) );
  MUX2_X1 U439 ( .A(\REGISTERS[5][6] ), .B(\REGISTERS[21][6] ), .S(n104), .Z(
        n429) );
  MUX2_X1 U440 ( .A(n429), .B(n428), .S(n78), .Z(n430) );
  MUX2_X1 U441 ( .A(\REGISTERS[9][6] ), .B(\REGISTERS[25][6] ), .S(n104), .Z(
        n431) );
  MUX2_X1 U442 ( .A(\REGISTERS[1][6] ), .B(\REGISTERS[17][6] ), .S(n104), .Z(
        n432) );
  MUX2_X1 U443 ( .A(n432), .B(n431), .S(n78), .Z(n433) );
  MUX2_X1 U444 ( .A(n433), .B(n430), .S(n65), .Z(n434) );
  MUX2_X1 U445 ( .A(\REGISTERS[12][6] ), .B(\REGISTERS[28][6] ), .S(n105), .Z(
        n435) );
  MUX2_X1 U446 ( .A(\REGISTERS[4][6] ), .B(\REGISTERS[20][6] ), .S(n105), .Z(
        n436) );
  MUX2_X1 U447 ( .A(n436), .B(n435), .S(n78), .Z(n437) );
  MUX2_X1 U448 ( .A(\REGISTERS[8][6] ), .B(\REGISTERS[24][6] ), .S(n105), .Z(
        n438) );
  MUX2_X1 U449 ( .A(\REGISTERS[0][6] ), .B(\REGISTERS[16][6] ), .S(n105), .Z(
        n439) );
  MUX2_X1 U450 ( .A(n439), .B(n438), .S(n78), .Z(n440) );
  MUX2_X1 U451 ( .A(n440), .B(n437), .S(n65), .Z(n441) );
  MUX2_X1 U452 ( .A(n441), .B(n434), .S(ADD_RD2[0]), .Z(n442) );
  MUX2_X1 U453 ( .A(n442), .B(n427), .S(ADD_RD2[1]), .Z(N418) );
  MUX2_X1 U454 ( .A(\REGISTERS[15][7] ), .B(\REGISTERS[31][7] ), .S(n105), .Z(
        n443) );
  MUX2_X1 U455 ( .A(\REGISTERS[7][7] ), .B(\REGISTERS[23][7] ), .S(n105), .Z(
        n444) );
  MUX2_X1 U456 ( .A(n444), .B(n443), .S(n78), .Z(n445) );
  MUX2_X1 U457 ( .A(\REGISTERS[11][7] ), .B(\REGISTERS[27][7] ), .S(n105), .Z(
        n446) );
  MUX2_X1 U458 ( .A(\REGISTERS[3][7] ), .B(\REGISTERS[19][7] ), .S(n105), .Z(
        n447) );
  MUX2_X1 U459 ( .A(n447), .B(n446), .S(n78), .Z(n448) );
  MUX2_X1 U460 ( .A(n448), .B(n445), .S(n65), .Z(n449) );
  MUX2_X1 U461 ( .A(\REGISTERS[14][7] ), .B(\REGISTERS[30][7] ), .S(n105), .Z(
        n450) );
  MUX2_X1 U462 ( .A(\REGISTERS[6][7] ), .B(\REGISTERS[22][7] ), .S(n105), .Z(
        n451) );
  MUX2_X1 U463 ( .A(n451), .B(n450), .S(n78), .Z(n452) );
  MUX2_X1 U464 ( .A(\REGISTERS[10][7] ), .B(\REGISTERS[26][7] ), .S(n105), .Z(
        n453) );
  MUX2_X1 U465 ( .A(\REGISTERS[2][7] ), .B(\REGISTERS[18][7] ), .S(n105), .Z(
        n454) );
  MUX2_X1 U466 ( .A(n454), .B(n453), .S(n78), .Z(n455) );
  MUX2_X1 U467 ( .A(n455), .B(n452), .S(n65), .Z(n456) );
  MUX2_X1 U468 ( .A(n456), .B(n449), .S(ADD_RD2[0]), .Z(n457) );
  MUX2_X1 U469 ( .A(\REGISTERS[13][7] ), .B(\REGISTERS[29][7] ), .S(n106), .Z(
        n458) );
  MUX2_X1 U470 ( .A(\REGISTERS[5][7] ), .B(\REGISTERS[21][7] ), .S(n106), .Z(
        n459) );
  MUX2_X1 U471 ( .A(n459), .B(n458), .S(n79), .Z(n460) );
  MUX2_X1 U472 ( .A(\REGISTERS[9][7] ), .B(\REGISTERS[25][7] ), .S(n106), .Z(
        n461) );
  MUX2_X1 U473 ( .A(\REGISTERS[1][7] ), .B(\REGISTERS[17][7] ), .S(n106), .Z(
        n462) );
  MUX2_X1 U474 ( .A(n462), .B(n461), .S(n79), .Z(n463) );
  MUX2_X1 U475 ( .A(n463), .B(n460), .S(n65), .Z(n464) );
  MUX2_X1 U476 ( .A(\REGISTERS[12][7] ), .B(\REGISTERS[28][7] ), .S(n106), .Z(
        n465) );
  MUX2_X1 U477 ( .A(\REGISTERS[4][7] ), .B(\REGISTERS[20][7] ), .S(n106), .Z(
        n466) );
  MUX2_X1 U478 ( .A(n466), .B(n465), .S(n79), .Z(n467) );
  MUX2_X1 U479 ( .A(\REGISTERS[8][7] ), .B(\REGISTERS[24][7] ), .S(n106), .Z(
        n468) );
  MUX2_X1 U480 ( .A(\REGISTERS[0][7] ), .B(\REGISTERS[16][7] ), .S(n106), .Z(
        n469) );
  MUX2_X1 U481 ( .A(n469), .B(n468), .S(n79), .Z(n470) );
  MUX2_X1 U482 ( .A(n470), .B(n467), .S(n65), .Z(n471) );
  MUX2_X1 U483 ( .A(n471), .B(n464), .S(ADD_RD2[0]), .Z(n472) );
  MUX2_X1 U484 ( .A(n472), .B(n457), .S(ADD_RD2[1]), .Z(N419) );
  MUX2_X1 U485 ( .A(\REGISTERS[15][8] ), .B(\REGISTERS[31][8] ), .S(n106), .Z(
        n473) );
  MUX2_X1 U486 ( .A(\REGISTERS[7][8] ), .B(\REGISTERS[23][8] ), .S(n106), .Z(
        n474) );
  MUX2_X1 U487 ( .A(n474), .B(n473), .S(n79), .Z(n475) );
  MUX2_X1 U488 ( .A(\REGISTERS[11][8] ), .B(\REGISTERS[27][8] ), .S(n106), .Z(
        n476) );
  MUX2_X1 U489 ( .A(\REGISTERS[3][8] ), .B(\REGISTERS[19][8] ), .S(n106), .Z(
        n477) );
  MUX2_X1 U490 ( .A(n477), .B(n476), .S(n79), .Z(n478) );
  MUX2_X1 U491 ( .A(n478), .B(n475), .S(n65), .Z(n479) );
  MUX2_X1 U492 ( .A(\REGISTERS[14][8] ), .B(\REGISTERS[30][8] ), .S(n107), .Z(
        n480) );
  MUX2_X1 U493 ( .A(\REGISTERS[6][8] ), .B(\REGISTERS[22][8] ), .S(n107), .Z(
        n481) );
  MUX2_X1 U494 ( .A(n481), .B(n480), .S(n79), .Z(n482) );
  MUX2_X1 U495 ( .A(\REGISTERS[10][8] ), .B(\REGISTERS[26][8] ), .S(n107), .Z(
        n483) );
  MUX2_X1 U496 ( .A(\REGISTERS[2][8] ), .B(\REGISTERS[18][8] ), .S(n107), .Z(
        n484) );
  MUX2_X1 U497 ( .A(n484), .B(n483), .S(n79), .Z(n485) );
  MUX2_X1 U498 ( .A(n485), .B(n482), .S(n65), .Z(n486) );
  MUX2_X1 U499 ( .A(n486), .B(n479), .S(ADD_RD2[0]), .Z(n487) );
  MUX2_X1 U500 ( .A(\REGISTERS[13][8] ), .B(\REGISTERS[29][8] ), .S(n107), .Z(
        n488) );
  MUX2_X1 U501 ( .A(\REGISTERS[5][8] ), .B(\REGISTERS[21][8] ), .S(n107), .Z(
        n489) );
  MUX2_X1 U502 ( .A(n489), .B(n488), .S(n79), .Z(n490) );
  MUX2_X1 U503 ( .A(\REGISTERS[9][8] ), .B(\REGISTERS[25][8] ), .S(n107), .Z(
        n491) );
  MUX2_X1 U504 ( .A(\REGISTERS[1][8] ), .B(\REGISTERS[17][8] ), .S(n107), .Z(
        n492) );
  MUX2_X1 U505 ( .A(n492), .B(n491), .S(n79), .Z(n493) );
  MUX2_X1 U506 ( .A(n493), .B(n490), .S(n65), .Z(n494) );
  MUX2_X1 U507 ( .A(\REGISTERS[12][8] ), .B(\REGISTERS[28][8] ), .S(n107), .Z(
        n495) );
  MUX2_X1 U508 ( .A(\REGISTERS[4][8] ), .B(\REGISTERS[20][8] ), .S(n107), .Z(
        n496) );
  MUX2_X1 U509 ( .A(n496), .B(n495), .S(n79), .Z(n497) );
  MUX2_X1 U510 ( .A(\REGISTERS[8][8] ), .B(\REGISTERS[24][8] ), .S(n107), .Z(
        n498) );
  MUX2_X1 U511 ( .A(\REGISTERS[0][8] ), .B(\REGISTERS[16][8] ), .S(n107), .Z(
        n499) );
  MUX2_X1 U512 ( .A(n499), .B(n498), .S(n79), .Z(n500) );
  MUX2_X1 U513 ( .A(n500), .B(n497), .S(n65), .Z(n501) );
  MUX2_X1 U514 ( .A(n501), .B(n494), .S(ADD_RD2[0]), .Z(n502) );
  MUX2_X1 U515 ( .A(n502), .B(n487), .S(ADD_RD2[1]), .Z(N420) );
  MUX2_X1 U516 ( .A(\REGISTERS[15][9] ), .B(\REGISTERS[31][9] ), .S(n108), .Z(
        n503) );
  MUX2_X1 U517 ( .A(\REGISTERS[7][9] ), .B(\REGISTERS[23][9] ), .S(n108), .Z(
        n504) );
  MUX2_X1 U518 ( .A(n504), .B(n503), .S(n80), .Z(n505) );
  MUX2_X1 U519 ( .A(\REGISTERS[11][9] ), .B(\REGISTERS[27][9] ), .S(n108), .Z(
        n506) );
  MUX2_X1 U520 ( .A(\REGISTERS[3][9] ), .B(\REGISTERS[19][9] ), .S(n108), .Z(
        n507) );
  MUX2_X1 U521 ( .A(n507), .B(n506), .S(n80), .Z(n508) );
  MUX2_X1 U522 ( .A(n508), .B(n505), .S(n66), .Z(n509) );
  MUX2_X1 U523 ( .A(\REGISTERS[14][9] ), .B(\REGISTERS[30][9] ), .S(n108), .Z(
        n510) );
  MUX2_X1 U524 ( .A(\REGISTERS[6][9] ), .B(\REGISTERS[22][9] ), .S(n108), .Z(
        n511) );
  MUX2_X1 U525 ( .A(n511), .B(n510), .S(n80), .Z(n512) );
  MUX2_X1 U526 ( .A(\REGISTERS[10][9] ), .B(\REGISTERS[26][9] ), .S(n108), .Z(
        n513) );
  MUX2_X1 U527 ( .A(\REGISTERS[2][9] ), .B(\REGISTERS[18][9] ), .S(n108), .Z(
        n514) );
  MUX2_X1 U528 ( .A(n514), .B(n513), .S(n80), .Z(n515) );
  MUX2_X1 U529 ( .A(n515), .B(n512), .S(n66), .Z(n516) );
  MUX2_X1 U530 ( .A(n516), .B(n509), .S(ADD_RD2[0]), .Z(n517) );
  MUX2_X1 U531 ( .A(\REGISTERS[13][9] ), .B(\REGISTERS[29][9] ), .S(n108), .Z(
        n518) );
  MUX2_X1 U532 ( .A(\REGISTERS[5][9] ), .B(\REGISTERS[21][9] ), .S(n108), .Z(
        n519) );
  MUX2_X1 U533 ( .A(n519), .B(n518), .S(n80), .Z(n520) );
  MUX2_X1 U534 ( .A(\REGISTERS[9][9] ), .B(\REGISTERS[25][9] ), .S(n108), .Z(
        n521) );
  MUX2_X1 U535 ( .A(\REGISTERS[1][9] ), .B(\REGISTERS[17][9] ), .S(n108), .Z(
        n522) );
  MUX2_X1 U536 ( .A(n522), .B(n521), .S(n80), .Z(n523) );
  MUX2_X1 U537 ( .A(n523), .B(n520), .S(n66), .Z(n524) );
  MUX2_X1 U538 ( .A(\REGISTERS[12][9] ), .B(\REGISTERS[28][9] ), .S(n109), .Z(
        n525) );
  MUX2_X1 U539 ( .A(\REGISTERS[4][9] ), .B(\REGISTERS[20][9] ), .S(n109), .Z(
        n526) );
  MUX2_X1 U540 ( .A(n526), .B(n525), .S(n80), .Z(n527) );
  MUX2_X1 U541 ( .A(\REGISTERS[8][9] ), .B(\REGISTERS[24][9] ), .S(n109), .Z(
        n528) );
  MUX2_X1 U542 ( .A(\REGISTERS[0][9] ), .B(\REGISTERS[16][9] ), .S(n109), .Z(
        n529) );
  MUX2_X1 U543 ( .A(n529), .B(n528), .S(n80), .Z(n530) );
  MUX2_X1 U544 ( .A(n530), .B(n527), .S(n66), .Z(n531) );
  MUX2_X1 U545 ( .A(n531), .B(n524), .S(ADD_RD2[0]), .Z(n532) );
  MUX2_X1 U546 ( .A(n532), .B(n517), .S(ADD_RD2[1]), .Z(N421) );
  MUX2_X1 U547 ( .A(\REGISTERS[15][10] ), .B(\REGISTERS[31][10] ), .S(n109), 
        .Z(n533) );
  MUX2_X1 U548 ( .A(\REGISTERS[7][10] ), .B(\REGISTERS[23][10] ), .S(n109), 
        .Z(n534) );
  MUX2_X1 U549 ( .A(n534), .B(n533), .S(n80), .Z(n535) );
  MUX2_X1 U550 ( .A(\REGISTERS[11][10] ), .B(\REGISTERS[27][10] ), .S(n109), 
        .Z(n536) );
  MUX2_X1 U551 ( .A(\REGISTERS[3][10] ), .B(\REGISTERS[19][10] ), .S(n109), 
        .Z(n537) );
  MUX2_X1 U552 ( .A(n537), .B(n536), .S(n80), .Z(n538) );
  MUX2_X1 U553 ( .A(n538), .B(n535), .S(n66), .Z(n539) );
  MUX2_X1 U554 ( .A(\REGISTERS[14][10] ), .B(\REGISTERS[30][10] ), .S(n109), 
        .Z(n540) );
  MUX2_X1 U555 ( .A(\REGISTERS[6][10] ), .B(\REGISTERS[22][10] ), .S(n109), 
        .Z(n541) );
  MUX2_X1 U556 ( .A(n541), .B(n540), .S(n80), .Z(n542) );
  MUX2_X1 U557 ( .A(\REGISTERS[10][10] ), .B(\REGISTERS[26][10] ), .S(n109), 
        .Z(n543) );
  MUX2_X1 U558 ( .A(\REGISTERS[2][10] ), .B(\REGISTERS[18][10] ), .S(n109), 
        .Z(n544) );
  MUX2_X1 U559 ( .A(n544), .B(n543), .S(n80), .Z(n545) );
  MUX2_X1 U560 ( .A(n545), .B(n542), .S(n66), .Z(n546) );
  MUX2_X1 U561 ( .A(n546), .B(n539), .S(ADD_RD2[0]), .Z(n547) );
  MUX2_X1 U562 ( .A(\REGISTERS[13][10] ), .B(\REGISTERS[29][10] ), .S(n110), 
        .Z(n548) );
  MUX2_X1 U563 ( .A(\REGISTERS[5][10] ), .B(\REGISTERS[21][10] ), .S(n110), 
        .Z(n549) );
  MUX2_X1 U564 ( .A(n549), .B(n548), .S(n81), .Z(n550) );
  MUX2_X1 U565 ( .A(\REGISTERS[9][10] ), .B(\REGISTERS[25][10] ), .S(n110), 
        .Z(n551) );
  MUX2_X1 U566 ( .A(\REGISTERS[1][10] ), .B(\REGISTERS[17][10] ), .S(n110), 
        .Z(n552) );
  MUX2_X1 U567 ( .A(n552), .B(n551), .S(n81), .Z(n553) );
  MUX2_X1 U568 ( .A(n553), .B(n550), .S(n66), .Z(n554) );
  MUX2_X1 U569 ( .A(\REGISTERS[12][10] ), .B(\REGISTERS[28][10] ), .S(n110), 
        .Z(n555) );
  MUX2_X1 U570 ( .A(\REGISTERS[4][10] ), .B(\REGISTERS[20][10] ), .S(n110), 
        .Z(n556) );
  MUX2_X1 U571 ( .A(n556), .B(n555), .S(n81), .Z(n557) );
  MUX2_X1 U572 ( .A(\REGISTERS[8][10] ), .B(\REGISTERS[24][10] ), .S(n110), 
        .Z(n558) );
  MUX2_X1 U573 ( .A(\REGISTERS[0][10] ), .B(\REGISTERS[16][10] ), .S(n110), 
        .Z(n559) );
  MUX2_X1 U574 ( .A(n559), .B(n558), .S(n81), .Z(n560) );
  MUX2_X1 U575 ( .A(n560), .B(n557), .S(n66), .Z(n561) );
  MUX2_X1 U576 ( .A(n561), .B(n554), .S(ADD_RD2[0]), .Z(n562) );
  MUX2_X1 U577 ( .A(n562), .B(n547), .S(ADD_RD2[1]), .Z(N422) );
  MUX2_X1 U578 ( .A(\REGISTERS[15][11] ), .B(\REGISTERS[31][11] ), .S(n110), 
        .Z(n563) );
  MUX2_X1 U579 ( .A(\REGISTERS[7][11] ), .B(\REGISTERS[23][11] ), .S(n110), 
        .Z(n564) );
  MUX2_X1 U580 ( .A(n564), .B(n563), .S(n81), .Z(n565) );
  MUX2_X1 U581 ( .A(\REGISTERS[11][11] ), .B(\REGISTERS[27][11] ), .S(n110), 
        .Z(n566) );
  MUX2_X1 U582 ( .A(\REGISTERS[3][11] ), .B(\REGISTERS[19][11] ), .S(n110), 
        .Z(n567) );
  MUX2_X1 U583 ( .A(n567), .B(n566), .S(n81), .Z(n568) );
  MUX2_X1 U584 ( .A(n568), .B(n565), .S(n66), .Z(n569) );
  MUX2_X1 U585 ( .A(\REGISTERS[14][11] ), .B(\REGISTERS[30][11] ), .S(n111), 
        .Z(n570) );
  MUX2_X1 U586 ( .A(\REGISTERS[6][11] ), .B(\REGISTERS[22][11] ), .S(n111), 
        .Z(n571) );
  MUX2_X1 U587 ( .A(n571), .B(n570), .S(n81), .Z(n572) );
  MUX2_X1 U588 ( .A(\REGISTERS[10][11] ), .B(\REGISTERS[26][11] ), .S(n111), 
        .Z(n573) );
  MUX2_X1 U589 ( .A(\REGISTERS[2][11] ), .B(\REGISTERS[18][11] ), .S(n111), 
        .Z(n574) );
  MUX2_X1 U590 ( .A(n574), .B(n573), .S(n81), .Z(n575) );
  MUX2_X1 U591 ( .A(n575), .B(n572), .S(n66), .Z(n576) );
  MUX2_X1 U592 ( .A(n576), .B(n569), .S(ADD_RD2[0]), .Z(n577) );
  MUX2_X1 U593 ( .A(\REGISTERS[13][11] ), .B(\REGISTERS[29][11] ), .S(n111), 
        .Z(n578) );
  MUX2_X1 U594 ( .A(\REGISTERS[5][11] ), .B(\REGISTERS[21][11] ), .S(n111), 
        .Z(n579) );
  MUX2_X1 U595 ( .A(n579), .B(n578), .S(n81), .Z(n580) );
  MUX2_X1 U596 ( .A(\REGISTERS[9][11] ), .B(\REGISTERS[25][11] ), .S(n111), 
        .Z(n581) );
  MUX2_X1 U597 ( .A(\REGISTERS[1][11] ), .B(\REGISTERS[17][11] ), .S(n111), 
        .Z(n582) );
  MUX2_X1 U598 ( .A(n582), .B(n581), .S(n81), .Z(n583) );
  MUX2_X1 U599 ( .A(n583), .B(n580), .S(n66), .Z(n584) );
  MUX2_X1 U600 ( .A(\REGISTERS[12][11] ), .B(\REGISTERS[28][11] ), .S(n111), 
        .Z(n585) );
  MUX2_X1 U601 ( .A(\REGISTERS[4][11] ), .B(\REGISTERS[20][11] ), .S(n111), 
        .Z(n586) );
  MUX2_X1 U602 ( .A(n586), .B(n585), .S(n81), .Z(n587) );
  MUX2_X1 U603 ( .A(\REGISTERS[8][11] ), .B(\REGISTERS[24][11] ), .S(n111), 
        .Z(n588) );
  MUX2_X1 U604 ( .A(\REGISTERS[0][11] ), .B(\REGISTERS[16][11] ), .S(n111), 
        .Z(n589) );
  MUX2_X1 U605 ( .A(n589), .B(n588), .S(n81), .Z(n590) );
  MUX2_X1 U606 ( .A(n590), .B(n587), .S(n66), .Z(n591) );
  MUX2_X1 U607 ( .A(n591), .B(n584), .S(ADD_RD2[0]), .Z(n592) );
  MUX2_X1 U608 ( .A(n592), .B(n577), .S(ADD_RD2[1]), .Z(N423) );
  MUX2_X1 U609 ( .A(\REGISTERS[15][12] ), .B(\REGISTERS[31][12] ), .S(n112), 
        .Z(n593) );
  MUX2_X1 U610 ( .A(\REGISTERS[7][12] ), .B(\REGISTERS[23][12] ), .S(n112), 
        .Z(n594) );
  MUX2_X1 U611 ( .A(n594), .B(n593), .S(n82), .Z(n595) );
  MUX2_X1 U612 ( .A(\REGISTERS[11][12] ), .B(\REGISTERS[27][12] ), .S(n112), 
        .Z(n596) );
  MUX2_X1 U613 ( .A(\REGISTERS[3][12] ), .B(\REGISTERS[19][12] ), .S(n112), 
        .Z(n597) );
  MUX2_X1 U614 ( .A(n597), .B(n596), .S(n82), .Z(n598) );
  MUX2_X1 U615 ( .A(n598), .B(n595), .S(n67), .Z(n599) );
  MUX2_X1 U616 ( .A(\REGISTERS[14][12] ), .B(\REGISTERS[30][12] ), .S(n112), 
        .Z(n600) );
  MUX2_X1 U617 ( .A(\REGISTERS[6][12] ), .B(\REGISTERS[22][12] ), .S(n112), 
        .Z(n601) );
  MUX2_X1 U618 ( .A(n601), .B(n600), .S(n82), .Z(n602) );
  MUX2_X1 U619 ( .A(\REGISTERS[10][12] ), .B(\REGISTERS[26][12] ), .S(n112), 
        .Z(n603) );
  MUX2_X1 U620 ( .A(\REGISTERS[2][12] ), .B(\REGISTERS[18][12] ), .S(n112), 
        .Z(n604) );
  MUX2_X1 U621 ( .A(n604), .B(n603), .S(n82), .Z(n605) );
  MUX2_X1 U622 ( .A(n605), .B(n602), .S(n67), .Z(n606) );
  MUX2_X1 U623 ( .A(n606), .B(n599), .S(ADD_RD2[0]), .Z(n607) );
  MUX2_X1 U624 ( .A(\REGISTERS[13][12] ), .B(\REGISTERS[29][12] ), .S(n112), 
        .Z(n608) );
  MUX2_X1 U625 ( .A(\REGISTERS[5][12] ), .B(\REGISTERS[21][12] ), .S(n112), 
        .Z(n609) );
  MUX2_X1 U626 ( .A(n609), .B(n608), .S(n82), .Z(n610) );
  MUX2_X1 U627 ( .A(\REGISTERS[9][12] ), .B(\REGISTERS[25][12] ), .S(n112), 
        .Z(n611) );
  MUX2_X1 U628 ( .A(\REGISTERS[1][12] ), .B(\REGISTERS[17][12] ), .S(n112), 
        .Z(n612) );
  MUX2_X1 U629 ( .A(n612), .B(n611), .S(n82), .Z(n613) );
  MUX2_X1 U630 ( .A(n613), .B(n610), .S(n67), .Z(n614) );
  MUX2_X1 U631 ( .A(\REGISTERS[12][12] ), .B(\REGISTERS[28][12] ), .S(n113), 
        .Z(n615) );
  MUX2_X1 U632 ( .A(\REGISTERS[4][12] ), .B(\REGISTERS[20][12] ), .S(n113), 
        .Z(n616) );
  MUX2_X1 U633 ( .A(n616), .B(n615), .S(n82), .Z(n617) );
  MUX2_X1 U634 ( .A(\REGISTERS[8][12] ), .B(\REGISTERS[24][12] ), .S(n113), 
        .Z(n618) );
  MUX2_X1 U635 ( .A(\REGISTERS[0][12] ), .B(\REGISTERS[16][12] ), .S(n113), 
        .Z(n619) );
  MUX2_X1 U636 ( .A(n619), .B(n618), .S(n82), .Z(n620) );
  MUX2_X1 U637 ( .A(n620), .B(n617), .S(n67), .Z(n621) );
  MUX2_X1 U638 ( .A(n621), .B(n614), .S(ADD_RD2[0]), .Z(n622) );
  MUX2_X1 U639 ( .A(n622), .B(n607), .S(ADD_RD2[1]), .Z(N424) );
  MUX2_X1 U640 ( .A(\REGISTERS[15][13] ), .B(\REGISTERS[31][13] ), .S(n113), 
        .Z(n623) );
  MUX2_X1 U641 ( .A(\REGISTERS[7][13] ), .B(\REGISTERS[23][13] ), .S(n113), 
        .Z(n624) );
  MUX2_X1 U642 ( .A(n624), .B(n623), .S(n82), .Z(n625) );
  MUX2_X1 U643 ( .A(\REGISTERS[11][13] ), .B(\REGISTERS[27][13] ), .S(n113), 
        .Z(n626) );
  MUX2_X1 U644 ( .A(\REGISTERS[3][13] ), .B(\REGISTERS[19][13] ), .S(n113), 
        .Z(n627) );
  MUX2_X1 U645 ( .A(n627), .B(n626), .S(n82), .Z(n628) );
  MUX2_X1 U646 ( .A(n628), .B(n625), .S(n67), .Z(n629) );
  MUX2_X1 U647 ( .A(\REGISTERS[14][13] ), .B(\REGISTERS[30][13] ), .S(n113), 
        .Z(n630) );
  MUX2_X1 U648 ( .A(\REGISTERS[6][13] ), .B(\REGISTERS[22][13] ), .S(n113), 
        .Z(n631) );
  MUX2_X1 U649 ( .A(n631), .B(n630), .S(n82), .Z(n632) );
  MUX2_X1 U650 ( .A(\REGISTERS[10][13] ), .B(\REGISTERS[26][13] ), .S(n113), 
        .Z(n633) );
  MUX2_X1 U651 ( .A(\REGISTERS[2][13] ), .B(\REGISTERS[18][13] ), .S(n113), 
        .Z(n634) );
  MUX2_X1 U652 ( .A(n634), .B(n633), .S(n82), .Z(n635) );
  MUX2_X1 U653 ( .A(n635), .B(n632), .S(n67), .Z(n636) );
  MUX2_X1 U654 ( .A(n636), .B(n629), .S(ADD_RD2[0]), .Z(n637) );
  MUX2_X1 U655 ( .A(\REGISTERS[13][13] ), .B(\REGISTERS[29][13] ), .S(n114), 
        .Z(n638) );
  MUX2_X1 U656 ( .A(\REGISTERS[5][13] ), .B(\REGISTERS[21][13] ), .S(n114), 
        .Z(n639) );
  MUX2_X1 U657 ( .A(n639), .B(n638), .S(n83), .Z(n640) );
  MUX2_X1 U658 ( .A(\REGISTERS[9][13] ), .B(\REGISTERS[25][13] ), .S(n114), 
        .Z(n641) );
  MUX2_X1 U659 ( .A(\REGISTERS[1][13] ), .B(\REGISTERS[17][13] ), .S(n114), 
        .Z(n642) );
  MUX2_X1 U660 ( .A(n642), .B(n641), .S(n83), .Z(n643) );
  MUX2_X1 U661 ( .A(n643), .B(n640), .S(n67), .Z(n644) );
  MUX2_X1 U662 ( .A(\REGISTERS[12][13] ), .B(\REGISTERS[28][13] ), .S(n114), 
        .Z(n645) );
  MUX2_X1 U663 ( .A(\REGISTERS[4][13] ), .B(\REGISTERS[20][13] ), .S(n114), 
        .Z(n646) );
  MUX2_X1 U664 ( .A(n646), .B(n645), .S(n83), .Z(n647) );
  MUX2_X1 U665 ( .A(\REGISTERS[8][13] ), .B(\REGISTERS[24][13] ), .S(n114), 
        .Z(n648) );
  MUX2_X1 U666 ( .A(\REGISTERS[0][13] ), .B(\REGISTERS[16][13] ), .S(n114), 
        .Z(n649) );
  MUX2_X1 U667 ( .A(n649), .B(n648), .S(n83), .Z(n650) );
  MUX2_X1 U668 ( .A(n650), .B(n647), .S(n67), .Z(n651) );
  MUX2_X1 U669 ( .A(n651), .B(n644), .S(ADD_RD2[0]), .Z(n652) );
  MUX2_X1 U670 ( .A(n652), .B(n637), .S(ADD_RD2[1]), .Z(N425) );
  MUX2_X1 U671 ( .A(\REGISTERS[15][14] ), .B(\REGISTERS[31][14] ), .S(n114), 
        .Z(n653) );
  MUX2_X1 U672 ( .A(\REGISTERS[7][14] ), .B(\REGISTERS[23][14] ), .S(n114), 
        .Z(n654) );
  MUX2_X1 U673 ( .A(n654), .B(n653), .S(n83), .Z(n655) );
  MUX2_X1 U674 ( .A(\REGISTERS[11][14] ), .B(\REGISTERS[27][14] ), .S(n114), 
        .Z(n656) );
  MUX2_X1 U675 ( .A(\REGISTERS[3][14] ), .B(\REGISTERS[19][14] ), .S(n114), 
        .Z(n657) );
  MUX2_X1 U676 ( .A(n657), .B(n656), .S(n83), .Z(n658) );
  MUX2_X1 U677 ( .A(n658), .B(n655), .S(n67), .Z(n659) );
  MUX2_X1 U678 ( .A(\REGISTERS[14][14] ), .B(\REGISTERS[30][14] ), .S(n115), 
        .Z(n660) );
  MUX2_X1 U679 ( .A(\REGISTERS[6][14] ), .B(\REGISTERS[22][14] ), .S(n115), 
        .Z(n661) );
  MUX2_X1 U680 ( .A(n661), .B(n660), .S(n83), .Z(n662) );
  MUX2_X1 U681 ( .A(\REGISTERS[10][14] ), .B(\REGISTERS[26][14] ), .S(n115), 
        .Z(n663) );
  MUX2_X1 U682 ( .A(\REGISTERS[2][14] ), .B(\REGISTERS[18][14] ), .S(n115), 
        .Z(n664) );
  MUX2_X1 U683 ( .A(n664), .B(n663), .S(n83), .Z(n665) );
  MUX2_X1 U684 ( .A(n665), .B(n662), .S(n67), .Z(n666) );
  MUX2_X1 U685 ( .A(n666), .B(n659), .S(ADD_RD2[0]), .Z(n667) );
  MUX2_X1 U686 ( .A(\REGISTERS[13][14] ), .B(\REGISTERS[29][14] ), .S(n115), 
        .Z(n668) );
  MUX2_X1 U687 ( .A(\REGISTERS[5][14] ), .B(\REGISTERS[21][14] ), .S(n115), 
        .Z(n669) );
  MUX2_X1 U688 ( .A(n669), .B(n668), .S(n83), .Z(n670) );
  MUX2_X1 U689 ( .A(\REGISTERS[9][14] ), .B(\REGISTERS[25][14] ), .S(n115), 
        .Z(n671) );
  MUX2_X1 U690 ( .A(\REGISTERS[1][14] ), .B(\REGISTERS[17][14] ), .S(n115), 
        .Z(n672) );
  MUX2_X1 U691 ( .A(n672), .B(n671), .S(n83), .Z(n673) );
  MUX2_X1 U692 ( .A(n673), .B(n670), .S(n67), .Z(n674) );
  MUX2_X1 U693 ( .A(\REGISTERS[12][14] ), .B(\REGISTERS[28][14] ), .S(n115), 
        .Z(n675) );
  MUX2_X1 U694 ( .A(\REGISTERS[4][14] ), .B(\REGISTERS[20][14] ), .S(n115), 
        .Z(n676) );
  MUX2_X1 U695 ( .A(n676), .B(n675), .S(n83), .Z(n677) );
  MUX2_X1 U696 ( .A(\REGISTERS[8][14] ), .B(\REGISTERS[24][14] ), .S(n115), 
        .Z(n678) );
  MUX2_X1 U697 ( .A(\REGISTERS[0][14] ), .B(\REGISTERS[16][14] ), .S(n115), 
        .Z(n679) );
  MUX2_X1 U698 ( .A(n679), .B(n678), .S(n83), .Z(n680) );
  MUX2_X1 U699 ( .A(n680), .B(n677), .S(n67), .Z(n681) );
  MUX2_X1 U700 ( .A(n681), .B(n674), .S(ADD_RD2[0]), .Z(n682) );
  MUX2_X1 U701 ( .A(n682), .B(n667), .S(ADD_RD2[1]), .Z(N426) );
  MUX2_X1 U702 ( .A(\REGISTERS[15][15] ), .B(\REGISTERS[31][15] ), .S(n116), 
        .Z(n683) );
  MUX2_X1 U703 ( .A(\REGISTERS[7][15] ), .B(\REGISTERS[23][15] ), .S(n116), 
        .Z(n684) );
  MUX2_X1 U704 ( .A(n684), .B(n683), .S(n84), .Z(n685) );
  MUX2_X1 U705 ( .A(\REGISTERS[11][15] ), .B(\REGISTERS[27][15] ), .S(n116), 
        .Z(n686) );
  MUX2_X1 U706 ( .A(\REGISTERS[3][15] ), .B(\REGISTERS[19][15] ), .S(n116), 
        .Z(n687) );
  MUX2_X1 U707 ( .A(n687), .B(n686), .S(n84), .Z(n688) );
  MUX2_X1 U708 ( .A(n688), .B(n685), .S(n68), .Z(n689) );
  MUX2_X1 U709 ( .A(\REGISTERS[14][15] ), .B(\REGISTERS[30][15] ), .S(n116), 
        .Z(n690) );
  MUX2_X1 U710 ( .A(\REGISTERS[6][15] ), .B(\REGISTERS[22][15] ), .S(n116), 
        .Z(n691) );
  MUX2_X1 U711 ( .A(n691), .B(n690), .S(n84), .Z(n692) );
  MUX2_X1 U712 ( .A(\REGISTERS[10][15] ), .B(\REGISTERS[26][15] ), .S(n116), 
        .Z(n693) );
  MUX2_X1 U713 ( .A(\REGISTERS[2][15] ), .B(\REGISTERS[18][15] ), .S(n116), 
        .Z(n694) );
  MUX2_X1 U714 ( .A(n694), .B(n693), .S(n84), .Z(n695) );
  MUX2_X1 U715 ( .A(n695), .B(n692), .S(n68), .Z(n696) );
  MUX2_X1 U716 ( .A(n696), .B(n689), .S(ADD_RD2[0]), .Z(n697) );
  MUX2_X1 U717 ( .A(\REGISTERS[13][15] ), .B(\REGISTERS[29][15] ), .S(n116), 
        .Z(n698) );
  MUX2_X1 U718 ( .A(\REGISTERS[5][15] ), .B(\REGISTERS[21][15] ), .S(n116), 
        .Z(n699) );
  MUX2_X1 U719 ( .A(n699), .B(n698), .S(n84), .Z(n700) );
  MUX2_X1 U720 ( .A(\REGISTERS[9][15] ), .B(\REGISTERS[25][15] ), .S(n116), 
        .Z(n701) );
  MUX2_X1 U721 ( .A(\REGISTERS[1][15] ), .B(\REGISTERS[17][15] ), .S(n116), 
        .Z(n702) );
  MUX2_X1 U722 ( .A(n702), .B(n701), .S(n84), .Z(n703) );
  MUX2_X1 U723 ( .A(n703), .B(n700), .S(n68), .Z(n704) );
  MUX2_X1 U724 ( .A(\REGISTERS[12][15] ), .B(\REGISTERS[28][15] ), .S(n117), 
        .Z(n705) );
  MUX2_X1 U725 ( .A(\REGISTERS[4][15] ), .B(\REGISTERS[20][15] ), .S(n117), 
        .Z(n706) );
  MUX2_X1 U726 ( .A(n706), .B(n705), .S(n84), .Z(n707) );
  MUX2_X1 U727 ( .A(\REGISTERS[8][15] ), .B(\REGISTERS[24][15] ), .S(n117), 
        .Z(n708) );
  MUX2_X1 U728 ( .A(\REGISTERS[0][15] ), .B(\REGISTERS[16][15] ), .S(n117), 
        .Z(n709) );
  MUX2_X1 U729 ( .A(n709), .B(n708), .S(n84), .Z(n710) );
  MUX2_X1 U730 ( .A(n710), .B(n707), .S(n68), .Z(n711) );
  MUX2_X1 U731 ( .A(n711), .B(n704), .S(ADD_RD2[0]), .Z(n712) );
  MUX2_X1 U732 ( .A(n712), .B(n697), .S(ADD_RD2[1]), .Z(N427) );
  MUX2_X1 U733 ( .A(\REGISTERS[15][16] ), .B(\REGISTERS[31][16] ), .S(n117), 
        .Z(n713) );
  MUX2_X1 U734 ( .A(\REGISTERS[7][16] ), .B(\REGISTERS[23][16] ), .S(n117), 
        .Z(n714) );
  MUX2_X1 U735 ( .A(n714), .B(n713), .S(n84), .Z(n715) );
  MUX2_X1 U736 ( .A(\REGISTERS[11][16] ), .B(\REGISTERS[27][16] ), .S(n117), 
        .Z(n716) );
  MUX2_X1 U737 ( .A(\REGISTERS[3][16] ), .B(\REGISTERS[19][16] ), .S(n117), 
        .Z(n717) );
  MUX2_X1 U738 ( .A(n717), .B(n716), .S(n84), .Z(n718) );
  MUX2_X1 U739 ( .A(n718), .B(n715), .S(n68), .Z(n719) );
  MUX2_X1 U740 ( .A(\REGISTERS[14][16] ), .B(\REGISTERS[30][16] ), .S(n117), 
        .Z(n720) );
  MUX2_X1 U741 ( .A(\REGISTERS[6][16] ), .B(\REGISTERS[22][16] ), .S(n117), 
        .Z(n721) );
  MUX2_X1 U742 ( .A(n721), .B(n720), .S(n84), .Z(n722) );
  MUX2_X1 U743 ( .A(\REGISTERS[10][16] ), .B(\REGISTERS[26][16] ), .S(n117), 
        .Z(n723) );
  MUX2_X1 U744 ( .A(\REGISTERS[2][16] ), .B(\REGISTERS[18][16] ), .S(n117), 
        .Z(n724) );
  MUX2_X1 U745 ( .A(n724), .B(n723), .S(n84), .Z(n725) );
  MUX2_X1 U746 ( .A(n725), .B(n722), .S(n68), .Z(n726) );
  MUX2_X1 U747 ( .A(n726), .B(n719), .S(ADD_RD2[0]), .Z(n727) );
  MUX2_X1 U748 ( .A(\REGISTERS[13][16] ), .B(\REGISTERS[29][16] ), .S(n118), 
        .Z(n728) );
  MUX2_X1 U749 ( .A(\REGISTERS[5][16] ), .B(\REGISTERS[21][16] ), .S(n118), 
        .Z(n729) );
  MUX2_X1 U750 ( .A(n729), .B(n728), .S(n85), .Z(n730) );
  MUX2_X1 U751 ( .A(\REGISTERS[9][16] ), .B(\REGISTERS[25][16] ), .S(n118), 
        .Z(n731) );
  MUX2_X1 U752 ( .A(\REGISTERS[1][16] ), .B(\REGISTERS[17][16] ), .S(n118), 
        .Z(n732) );
  MUX2_X1 U753 ( .A(n732), .B(n731), .S(n85), .Z(n733) );
  MUX2_X1 U754 ( .A(n733), .B(n730), .S(n68), .Z(n734) );
  MUX2_X1 U755 ( .A(\REGISTERS[12][16] ), .B(\REGISTERS[28][16] ), .S(n118), 
        .Z(n735) );
  MUX2_X1 U756 ( .A(\REGISTERS[4][16] ), .B(\REGISTERS[20][16] ), .S(n118), 
        .Z(n736) );
  MUX2_X1 U757 ( .A(n736), .B(n735), .S(n85), .Z(n737) );
  MUX2_X1 U758 ( .A(\REGISTERS[8][16] ), .B(\REGISTERS[24][16] ), .S(n118), 
        .Z(n738) );
  MUX2_X1 U759 ( .A(\REGISTERS[0][16] ), .B(\REGISTERS[16][16] ), .S(n118), 
        .Z(n739) );
  MUX2_X1 U760 ( .A(n739), .B(n738), .S(n85), .Z(n740) );
  MUX2_X1 U761 ( .A(n740), .B(n737), .S(n68), .Z(n741) );
  MUX2_X1 U762 ( .A(n741), .B(n734), .S(ADD_RD2[0]), .Z(n742) );
  MUX2_X1 U763 ( .A(n742), .B(n727), .S(ADD_RD2[1]), .Z(N428) );
  MUX2_X1 U764 ( .A(\REGISTERS[15][17] ), .B(\REGISTERS[31][17] ), .S(n118), 
        .Z(n743) );
  MUX2_X1 U765 ( .A(\REGISTERS[7][17] ), .B(\REGISTERS[23][17] ), .S(n118), 
        .Z(n744) );
  MUX2_X1 U766 ( .A(n744), .B(n743), .S(n85), .Z(n745) );
  MUX2_X1 U767 ( .A(\REGISTERS[11][17] ), .B(\REGISTERS[27][17] ), .S(n118), 
        .Z(n746) );
  MUX2_X1 U768 ( .A(\REGISTERS[3][17] ), .B(\REGISTERS[19][17] ), .S(n118), 
        .Z(n747) );
  MUX2_X1 U769 ( .A(n747), .B(n746), .S(n85), .Z(n748) );
  MUX2_X1 U770 ( .A(n748), .B(n745), .S(n68), .Z(n749) );
  MUX2_X1 U771 ( .A(\REGISTERS[14][17] ), .B(\REGISTERS[30][17] ), .S(n119), 
        .Z(n750) );
  MUX2_X1 U772 ( .A(\REGISTERS[6][17] ), .B(\REGISTERS[22][17] ), .S(n119), 
        .Z(n751) );
  MUX2_X1 U773 ( .A(n751), .B(n750), .S(n85), .Z(n752) );
  MUX2_X1 U774 ( .A(\REGISTERS[10][17] ), .B(\REGISTERS[26][17] ), .S(n119), 
        .Z(n753) );
  MUX2_X1 U775 ( .A(\REGISTERS[2][17] ), .B(\REGISTERS[18][17] ), .S(n119), 
        .Z(n754) );
  MUX2_X1 U776 ( .A(n754), .B(n753), .S(n85), .Z(n755) );
  MUX2_X1 U777 ( .A(n755), .B(n752), .S(n68), .Z(n756) );
  MUX2_X1 U778 ( .A(n756), .B(n749), .S(ADD_RD2[0]), .Z(n757) );
  MUX2_X1 U779 ( .A(\REGISTERS[13][17] ), .B(\REGISTERS[29][17] ), .S(n119), 
        .Z(n758) );
  MUX2_X1 U780 ( .A(\REGISTERS[5][17] ), .B(\REGISTERS[21][17] ), .S(n119), 
        .Z(n759) );
  MUX2_X1 U781 ( .A(n759), .B(n758), .S(n85), .Z(n760) );
  MUX2_X1 U782 ( .A(\REGISTERS[9][17] ), .B(\REGISTERS[25][17] ), .S(n119), 
        .Z(n761) );
  MUX2_X1 U783 ( .A(\REGISTERS[1][17] ), .B(\REGISTERS[17][17] ), .S(n119), 
        .Z(n762) );
  MUX2_X1 U784 ( .A(n762), .B(n761), .S(n85), .Z(n763) );
  MUX2_X1 U785 ( .A(n763), .B(n760), .S(n68), .Z(n764) );
  MUX2_X1 U786 ( .A(\REGISTERS[12][17] ), .B(\REGISTERS[28][17] ), .S(n119), 
        .Z(n765) );
  MUX2_X1 U787 ( .A(\REGISTERS[4][17] ), .B(\REGISTERS[20][17] ), .S(n119), 
        .Z(n766) );
  MUX2_X1 U788 ( .A(n766), .B(n765), .S(n85), .Z(n767) );
  MUX2_X1 U789 ( .A(\REGISTERS[8][17] ), .B(\REGISTERS[24][17] ), .S(n119), 
        .Z(n768) );
  MUX2_X1 U790 ( .A(\REGISTERS[0][17] ), .B(\REGISTERS[16][17] ), .S(n119), 
        .Z(n769) );
  MUX2_X1 U791 ( .A(n769), .B(n768), .S(n85), .Z(n770) );
  MUX2_X1 U792 ( .A(n770), .B(n767), .S(n68), .Z(n771) );
  MUX2_X1 U793 ( .A(n771), .B(n764), .S(ADD_RD2[0]), .Z(n772) );
  MUX2_X1 U794 ( .A(n772), .B(n757), .S(ADD_RD2[1]), .Z(N429) );
  MUX2_X1 U795 ( .A(\REGISTERS[15][18] ), .B(\REGISTERS[31][18] ), .S(n120), 
        .Z(n773) );
  MUX2_X1 U796 ( .A(\REGISTERS[7][18] ), .B(\REGISTERS[23][18] ), .S(n120), 
        .Z(n774) );
  MUX2_X1 U797 ( .A(n774), .B(n773), .S(n86), .Z(n775) );
  MUX2_X1 U798 ( .A(\REGISTERS[11][18] ), .B(\REGISTERS[27][18] ), .S(n120), 
        .Z(n776) );
  MUX2_X1 U799 ( .A(\REGISTERS[3][18] ), .B(\REGISTERS[19][18] ), .S(n120), 
        .Z(n777) );
  MUX2_X1 U800 ( .A(n777), .B(n776), .S(n86), .Z(n778) );
  MUX2_X1 U801 ( .A(n778), .B(n775), .S(n69), .Z(n779) );
  MUX2_X1 U802 ( .A(\REGISTERS[14][18] ), .B(\REGISTERS[30][18] ), .S(n120), 
        .Z(n780) );
  MUX2_X1 U803 ( .A(\REGISTERS[6][18] ), .B(\REGISTERS[22][18] ), .S(n120), 
        .Z(n781) );
  MUX2_X1 U804 ( .A(n781), .B(n780), .S(n86), .Z(n782) );
  MUX2_X1 U805 ( .A(\REGISTERS[10][18] ), .B(\REGISTERS[26][18] ), .S(n120), 
        .Z(n783) );
  MUX2_X1 U806 ( .A(\REGISTERS[2][18] ), .B(\REGISTERS[18][18] ), .S(n120), 
        .Z(n784) );
  MUX2_X1 U807 ( .A(n784), .B(n783), .S(n86), .Z(n785) );
  MUX2_X1 U808 ( .A(n785), .B(n782), .S(n69), .Z(n786) );
  MUX2_X1 U809 ( .A(n786), .B(n779), .S(ADD_RD2[0]), .Z(n787) );
  MUX2_X1 U810 ( .A(\REGISTERS[13][18] ), .B(\REGISTERS[29][18] ), .S(n120), 
        .Z(n788) );
  MUX2_X1 U811 ( .A(\REGISTERS[5][18] ), .B(\REGISTERS[21][18] ), .S(n120), 
        .Z(n789) );
  MUX2_X1 U812 ( .A(n789), .B(n788), .S(n86), .Z(n790) );
  MUX2_X1 U813 ( .A(\REGISTERS[9][18] ), .B(\REGISTERS[25][18] ), .S(n120), 
        .Z(n791) );
  MUX2_X1 U814 ( .A(\REGISTERS[1][18] ), .B(\REGISTERS[17][18] ), .S(n120), 
        .Z(n792) );
  MUX2_X1 U815 ( .A(n792), .B(n791), .S(n86), .Z(n793) );
  MUX2_X1 U816 ( .A(n793), .B(n790), .S(n69), .Z(n794) );
  MUX2_X1 U817 ( .A(\REGISTERS[12][18] ), .B(\REGISTERS[28][18] ), .S(n121), 
        .Z(n795) );
  MUX2_X1 U818 ( .A(\REGISTERS[4][18] ), .B(\REGISTERS[20][18] ), .S(n121), 
        .Z(n796) );
  MUX2_X1 U819 ( .A(n796), .B(n795), .S(n86), .Z(n797) );
  MUX2_X1 U820 ( .A(\REGISTERS[8][18] ), .B(\REGISTERS[24][18] ), .S(n121), 
        .Z(n798) );
  MUX2_X1 U821 ( .A(\REGISTERS[0][18] ), .B(\REGISTERS[16][18] ), .S(n121), 
        .Z(n799) );
  MUX2_X1 U822 ( .A(n799), .B(n798), .S(n86), .Z(n800) );
  MUX2_X1 U823 ( .A(n800), .B(n797), .S(n69), .Z(n801) );
  MUX2_X1 U824 ( .A(n801), .B(n794), .S(ADD_RD2[0]), .Z(n802) );
  MUX2_X1 U825 ( .A(n802), .B(n787), .S(ADD_RD2[1]), .Z(N430) );
  MUX2_X1 U826 ( .A(\REGISTERS[15][19] ), .B(\REGISTERS[31][19] ), .S(n121), 
        .Z(n803) );
  MUX2_X1 U827 ( .A(\REGISTERS[7][19] ), .B(\REGISTERS[23][19] ), .S(n121), 
        .Z(n804) );
  MUX2_X1 U828 ( .A(n804), .B(n803), .S(n86), .Z(n805) );
  MUX2_X1 U829 ( .A(\REGISTERS[11][19] ), .B(\REGISTERS[27][19] ), .S(n121), 
        .Z(n806) );
  MUX2_X1 U830 ( .A(\REGISTERS[3][19] ), .B(\REGISTERS[19][19] ), .S(n121), 
        .Z(n807) );
  MUX2_X1 U831 ( .A(n807), .B(n806), .S(n86), .Z(n808) );
  MUX2_X1 U832 ( .A(n808), .B(n805), .S(n69), .Z(n809) );
  MUX2_X1 U833 ( .A(\REGISTERS[14][19] ), .B(\REGISTERS[30][19] ), .S(n121), 
        .Z(n810) );
  MUX2_X1 U834 ( .A(\REGISTERS[6][19] ), .B(\REGISTERS[22][19] ), .S(n121), 
        .Z(n811) );
  MUX2_X1 U835 ( .A(n811), .B(n810), .S(n86), .Z(n812) );
  MUX2_X1 U836 ( .A(\REGISTERS[10][19] ), .B(\REGISTERS[26][19] ), .S(n121), 
        .Z(n813) );
  MUX2_X1 U837 ( .A(\REGISTERS[2][19] ), .B(\REGISTERS[18][19] ), .S(n121), 
        .Z(n814) );
  MUX2_X1 U838 ( .A(n814), .B(n813), .S(n86), .Z(n815) );
  MUX2_X1 U839 ( .A(n815), .B(n812), .S(n69), .Z(n816) );
  MUX2_X1 U840 ( .A(n816), .B(n809), .S(ADD_RD2[0]), .Z(n817) );
  MUX2_X1 U841 ( .A(\REGISTERS[13][19] ), .B(\REGISTERS[29][19] ), .S(n122), 
        .Z(n818) );
  MUX2_X1 U842 ( .A(\REGISTERS[5][19] ), .B(\REGISTERS[21][19] ), .S(n122), 
        .Z(n819) );
  MUX2_X1 U843 ( .A(n819), .B(n818), .S(n87), .Z(n820) );
  MUX2_X1 U844 ( .A(\REGISTERS[9][19] ), .B(\REGISTERS[25][19] ), .S(n122), 
        .Z(n821) );
  MUX2_X1 U845 ( .A(\REGISTERS[1][19] ), .B(\REGISTERS[17][19] ), .S(n122), 
        .Z(n822) );
  MUX2_X1 U846 ( .A(n822), .B(n821), .S(n87), .Z(n823) );
  MUX2_X1 U847 ( .A(n823), .B(n820), .S(n69), .Z(n824) );
  MUX2_X1 U848 ( .A(\REGISTERS[12][19] ), .B(\REGISTERS[28][19] ), .S(n122), 
        .Z(n825) );
  MUX2_X1 U849 ( .A(\REGISTERS[4][19] ), .B(\REGISTERS[20][19] ), .S(n122), 
        .Z(n826) );
  MUX2_X1 U850 ( .A(n826), .B(n825), .S(n87), .Z(n827) );
  MUX2_X1 U851 ( .A(\REGISTERS[8][19] ), .B(\REGISTERS[24][19] ), .S(n122), 
        .Z(n828) );
  MUX2_X1 U852 ( .A(\REGISTERS[0][19] ), .B(\REGISTERS[16][19] ), .S(n122), 
        .Z(n829) );
  MUX2_X1 U853 ( .A(n829), .B(n828), .S(n87), .Z(n830) );
  MUX2_X1 U854 ( .A(n830), .B(n827), .S(n69), .Z(n831) );
  MUX2_X1 U855 ( .A(n831), .B(n824), .S(ADD_RD2[0]), .Z(n832) );
  MUX2_X1 U856 ( .A(n832), .B(n817), .S(ADD_RD2[1]), .Z(N431) );
  MUX2_X1 U857 ( .A(\REGISTERS[15][20] ), .B(\REGISTERS[31][20] ), .S(n122), 
        .Z(n833) );
  MUX2_X1 U858 ( .A(\REGISTERS[7][20] ), .B(\REGISTERS[23][20] ), .S(n122), 
        .Z(n834) );
  MUX2_X1 U859 ( .A(n834), .B(n833), .S(n87), .Z(n835) );
  MUX2_X1 U860 ( .A(\REGISTERS[11][20] ), .B(\REGISTERS[27][20] ), .S(n122), 
        .Z(n836) );
  MUX2_X1 U861 ( .A(\REGISTERS[3][20] ), .B(\REGISTERS[19][20] ), .S(n122), 
        .Z(n837) );
  MUX2_X1 U862 ( .A(n837), .B(n836), .S(n87), .Z(n838) );
  MUX2_X1 U863 ( .A(n838), .B(n835), .S(n69), .Z(n839) );
  MUX2_X1 U864 ( .A(\REGISTERS[14][20] ), .B(\REGISTERS[30][20] ), .S(n123), 
        .Z(n840) );
  MUX2_X1 U865 ( .A(\REGISTERS[6][20] ), .B(\REGISTERS[22][20] ), .S(n123), 
        .Z(n841) );
  MUX2_X1 U866 ( .A(n841), .B(n840), .S(n87), .Z(n842) );
  MUX2_X1 U867 ( .A(\REGISTERS[10][20] ), .B(\REGISTERS[26][20] ), .S(n123), 
        .Z(n843) );
  MUX2_X1 U868 ( .A(\REGISTERS[2][20] ), .B(\REGISTERS[18][20] ), .S(n123), 
        .Z(n844) );
  MUX2_X1 U869 ( .A(n844), .B(n843), .S(n87), .Z(n845) );
  MUX2_X1 U870 ( .A(n845), .B(n842), .S(n69), .Z(n846) );
  MUX2_X1 U871 ( .A(n846), .B(n839), .S(ADD_RD2[0]), .Z(n847) );
  MUX2_X1 U872 ( .A(\REGISTERS[13][20] ), .B(\REGISTERS[29][20] ), .S(n123), 
        .Z(n848) );
  MUX2_X1 U873 ( .A(\REGISTERS[5][20] ), .B(\REGISTERS[21][20] ), .S(n123), 
        .Z(n849) );
  MUX2_X1 U874 ( .A(n849), .B(n848), .S(n87), .Z(n850) );
  MUX2_X1 U875 ( .A(\REGISTERS[9][20] ), .B(\REGISTERS[25][20] ), .S(n123), 
        .Z(n851) );
  MUX2_X1 U876 ( .A(\REGISTERS[1][20] ), .B(\REGISTERS[17][20] ), .S(n123), 
        .Z(n852) );
  MUX2_X1 U877 ( .A(n852), .B(n851), .S(n87), .Z(n853) );
  MUX2_X1 U878 ( .A(n853), .B(n850), .S(n69), .Z(n854) );
  MUX2_X1 U879 ( .A(\REGISTERS[12][20] ), .B(\REGISTERS[28][20] ), .S(n123), 
        .Z(n855) );
  MUX2_X1 U880 ( .A(\REGISTERS[4][20] ), .B(\REGISTERS[20][20] ), .S(n123), 
        .Z(n856) );
  MUX2_X1 U881 ( .A(n856), .B(n855), .S(n87), .Z(n857) );
  MUX2_X1 U882 ( .A(\REGISTERS[8][20] ), .B(\REGISTERS[24][20] ), .S(n123), 
        .Z(n858) );
  MUX2_X1 U883 ( .A(\REGISTERS[0][20] ), .B(\REGISTERS[16][20] ), .S(n123), 
        .Z(n859) );
  MUX2_X1 U884 ( .A(n859), .B(n858), .S(n87), .Z(n860) );
  MUX2_X1 U885 ( .A(n860), .B(n857), .S(n69), .Z(n861) );
  MUX2_X1 U886 ( .A(n861), .B(n854), .S(ADD_RD2[0]), .Z(n862) );
  MUX2_X1 U887 ( .A(n862), .B(n847), .S(ADD_RD2[1]), .Z(N432) );
  MUX2_X1 U888 ( .A(\REGISTERS[15][21] ), .B(\REGISTERS[31][21] ), .S(n124), 
        .Z(n863) );
  MUX2_X1 U889 ( .A(\REGISTERS[7][21] ), .B(\REGISTERS[23][21] ), .S(n124), 
        .Z(n864) );
  MUX2_X1 U890 ( .A(n864), .B(n863), .S(n88), .Z(n865) );
  MUX2_X1 U891 ( .A(\REGISTERS[11][21] ), .B(\REGISTERS[27][21] ), .S(n124), 
        .Z(n866) );
  MUX2_X1 U892 ( .A(\REGISTERS[3][21] ), .B(\REGISTERS[19][21] ), .S(n124), 
        .Z(n867) );
  MUX2_X1 U893 ( .A(n867), .B(n866), .S(n88), .Z(n868) );
  MUX2_X1 U894 ( .A(n868), .B(n865), .S(n70), .Z(n869) );
  MUX2_X1 U895 ( .A(\REGISTERS[14][21] ), .B(\REGISTERS[30][21] ), .S(n124), 
        .Z(n870) );
  MUX2_X1 U896 ( .A(\REGISTERS[6][21] ), .B(\REGISTERS[22][21] ), .S(n124), 
        .Z(n871) );
  MUX2_X1 U897 ( .A(n871), .B(n870), .S(n88), .Z(n872) );
  MUX2_X1 U898 ( .A(\REGISTERS[10][21] ), .B(\REGISTERS[26][21] ), .S(n124), 
        .Z(n873) );
  MUX2_X1 U899 ( .A(\REGISTERS[2][21] ), .B(\REGISTERS[18][21] ), .S(n124), 
        .Z(n874) );
  MUX2_X1 U900 ( .A(n874), .B(n873), .S(n88), .Z(n875) );
  MUX2_X1 U901 ( .A(n875), .B(n872), .S(n70), .Z(n876) );
  MUX2_X1 U902 ( .A(n876), .B(n869), .S(ADD_RD2[0]), .Z(n877) );
  MUX2_X1 U903 ( .A(\REGISTERS[13][21] ), .B(\REGISTERS[29][21] ), .S(n124), 
        .Z(n878) );
  MUX2_X1 U904 ( .A(\REGISTERS[5][21] ), .B(\REGISTERS[21][21] ), .S(n124), 
        .Z(n879) );
  MUX2_X1 U905 ( .A(n879), .B(n878), .S(n88), .Z(n880) );
  MUX2_X1 U906 ( .A(\REGISTERS[9][21] ), .B(\REGISTERS[25][21] ), .S(n124), 
        .Z(n881) );
  MUX2_X1 U907 ( .A(\REGISTERS[1][21] ), .B(\REGISTERS[17][21] ), .S(n124), 
        .Z(n882) );
  MUX2_X1 U908 ( .A(n882), .B(n881), .S(n88), .Z(n883) );
  MUX2_X1 U909 ( .A(n883), .B(n880), .S(n70), .Z(n884) );
  MUX2_X1 U910 ( .A(\REGISTERS[12][21] ), .B(\REGISTERS[28][21] ), .S(n125), 
        .Z(n885) );
  MUX2_X1 U911 ( .A(\REGISTERS[4][21] ), .B(\REGISTERS[20][21] ), .S(n125), 
        .Z(n886) );
  MUX2_X1 U912 ( .A(n886), .B(n885), .S(n88), .Z(n887) );
  MUX2_X1 U913 ( .A(\REGISTERS[8][21] ), .B(\REGISTERS[24][21] ), .S(n125), 
        .Z(n888) );
  MUX2_X1 U914 ( .A(\REGISTERS[0][21] ), .B(\REGISTERS[16][21] ), .S(n125), 
        .Z(n889) );
  MUX2_X1 U915 ( .A(n889), .B(n888), .S(n88), .Z(n890) );
  MUX2_X1 U916 ( .A(n890), .B(n887), .S(n70), .Z(n891) );
  MUX2_X1 U917 ( .A(n891), .B(n884), .S(ADD_RD2[0]), .Z(n892) );
  MUX2_X1 U918 ( .A(n892), .B(n877), .S(ADD_RD2[1]), .Z(N433) );
  MUX2_X1 U919 ( .A(\REGISTERS[15][22] ), .B(\REGISTERS[31][22] ), .S(n125), 
        .Z(n893) );
  MUX2_X1 U920 ( .A(\REGISTERS[7][22] ), .B(\REGISTERS[23][22] ), .S(n125), 
        .Z(n894) );
  MUX2_X1 U921 ( .A(n894), .B(n893), .S(n88), .Z(n895) );
  MUX2_X1 U922 ( .A(\REGISTERS[11][22] ), .B(\REGISTERS[27][22] ), .S(n125), 
        .Z(n896) );
  MUX2_X1 U923 ( .A(\REGISTERS[3][22] ), .B(\REGISTERS[19][22] ), .S(n125), 
        .Z(n897) );
  MUX2_X1 U924 ( .A(n897), .B(n896), .S(n88), .Z(n898) );
  MUX2_X1 U925 ( .A(n898), .B(n895), .S(n70), .Z(n899) );
  MUX2_X1 U926 ( .A(\REGISTERS[14][22] ), .B(\REGISTERS[30][22] ), .S(n125), 
        .Z(n900) );
  MUX2_X1 U927 ( .A(\REGISTERS[6][22] ), .B(\REGISTERS[22][22] ), .S(n125), 
        .Z(n901) );
  MUX2_X1 U928 ( .A(n901), .B(n900), .S(n88), .Z(n902) );
  MUX2_X1 U929 ( .A(\REGISTERS[10][22] ), .B(\REGISTERS[26][22] ), .S(n125), 
        .Z(n903) );
  MUX2_X1 U930 ( .A(\REGISTERS[2][22] ), .B(\REGISTERS[18][22] ), .S(n125), 
        .Z(n904) );
  MUX2_X1 U931 ( .A(n904), .B(n903), .S(n88), .Z(n905) );
  MUX2_X1 U932 ( .A(n905), .B(n902), .S(n70), .Z(n906) );
  MUX2_X1 U933 ( .A(n906), .B(n899), .S(ADD_RD2[0]), .Z(n907) );
  MUX2_X1 U934 ( .A(\REGISTERS[13][22] ), .B(\REGISTERS[29][22] ), .S(n126), 
        .Z(n908) );
  MUX2_X1 U935 ( .A(\REGISTERS[5][22] ), .B(\REGISTERS[21][22] ), .S(n126), 
        .Z(n909) );
  MUX2_X1 U936 ( .A(n909), .B(n908), .S(n89), .Z(n910) );
  MUX2_X1 U937 ( .A(\REGISTERS[9][22] ), .B(\REGISTERS[25][22] ), .S(n126), 
        .Z(n911) );
  MUX2_X1 U938 ( .A(\REGISTERS[1][22] ), .B(\REGISTERS[17][22] ), .S(n126), 
        .Z(n912) );
  MUX2_X1 U939 ( .A(n912), .B(n911), .S(n89), .Z(n913) );
  MUX2_X1 U940 ( .A(n913), .B(n910), .S(n70), .Z(n914) );
  MUX2_X1 U941 ( .A(\REGISTERS[12][22] ), .B(\REGISTERS[28][22] ), .S(n126), 
        .Z(n915) );
  MUX2_X1 U942 ( .A(\REGISTERS[4][22] ), .B(\REGISTERS[20][22] ), .S(n126), 
        .Z(n916) );
  MUX2_X1 U943 ( .A(n916), .B(n915), .S(n89), .Z(n917) );
  MUX2_X1 U944 ( .A(\REGISTERS[8][22] ), .B(\REGISTERS[24][22] ), .S(n126), 
        .Z(n918) );
  MUX2_X1 U945 ( .A(\REGISTERS[0][22] ), .B(\REGISTERS[16][22] ), .S(n126), 
        .Z(n919) );
  MUX2_X1 U946 ( .A(n919), .B(n918), .S(n89), .Z(n920) );
  MUX2_X1 U947 ( .A(n920), .B(n917), .S(n70), .Z(n921) );
  MUX2_X1 U948 ( .A(n921), .B(n914), .S(ADD_RD2[0]), .Z(n922) );
  MUX2_X1 U949 ( .A(n922), .B(n907), .S(ADD_RD2[1]), .Z(N434) );
  MUX2_X1 U950 ( .A(\REGISTERS[15][23] ), .B(\REGISTERS[31][23] ), .S(n126), 
        .Z(n923) );
  MUX2_X1 U951 ( .A(\REGISTERS[7][23] ), .B(\REGISTERS[23][23] ), .S(n126), 
        .Z(n924) );
  MUX2_X1 U952 ( .A(n924), .B(n923), .S(n89), .Z(n925) );
  MUX2_X1 U953 ( .A(\REGISTERS[11][23] ), .B(\REGISTERS[27][23] ), .S(n126), 
        .Z(n926) );
  MUX2_X1 U954 ( .A(\REGISTERS[3][23] ), .B(\REGISTERS[19][23] ), .S(n126), 
        .Z(n927) );
  MUX2_X1 U955 ( .A(n927), .B(n926), .S(n89), .Z(n928) );
  MUX2_X1 U956 ( .A(n928), .B(n925), .S(n70), .Z(n929) );
  MUX2_X1 U957 ( .A(\REGISTERS[14][23] ), .B(\REGISTERS[30][23] ), .S(n127), 
        .Z(n930) );
  MUX2_X1 U958 ( .A(\REGISTERS[6][23] ), .B(\REGISTERS[22][23] ), .S(n127), 
        .Z(n931) );
  MUX2_X1 U959 ( .A(n931), .B(n930), .S(n89), .Z(n932) );
  MUX2_X1 U960 ( .A(\REGISTERS[10][23] ), .B(\REGISTERS[26][23] ), .S(n127), 
        .Z(n933) );
  MUX2_X1 U961 ( .A(\REGISTERS[2][23] ), .B(\REGISTERS[18][23] ), .S(n127), 
        .Z(n934) );
  MUX2_X1 U962 ( .A(n934), .B(n933), .S(n89), .Z(n935) );
  MUX2_X1 U963 ( .A(n935), .B(n932), .S(n70), .Z(n936) );
  MUX2_X1 U964 ( .A(n936), .B(n929), .S(ADD_RD2[0]), .Z(n937) );
  MUX2_X1 U965 ( .A(\REGISTERS[13][23] ), .B(\REGISTERS[29][23] ), .S(n127), 
        .Z(n938) );
  MUX2_X1 U966 ( .A(\REGISTERS[5][23] ), .B(\REGISTERS[21][23] ), .S(n127), 
        .Z(n939) );
  MUX2_X1 U967 ( .A(n939), .B(n938), .S(n89), .Z(n940) );
  MUX2_X1 U968 ( .A(\REGISTERS[9][23] ), .B(\REGISTERS[25][23] ), .S(n127), 
        .Z(n941) );
  MUX2_X1 U969 ( .A(\REGISTERS[1][23] ), .B(\REGISTERS[17][23] ), .S(n127), 
        .Z(n942) );
  MUX2_X1 U970 ( .A(n942), .B(n941), .S(n89), .Z(n943) );
  MUX2_X1 U971 ( .A(n943), .B(n940), .S(n70), .Z(n944) );
  MUX2_X1 U972 ( .A(\REGISTERS[12][23] ), .B(\REGISTERS[28][23] ), .S(n127), 
        .Z(n945) );
  MUX2_X1 U973 ( .A(\REGISTERS[4][23] ), .B(\REGISTERS[20][23] ), .S(n127), 
        .Z(n946) );
  MUX2_X1 U974 ( .A(n946), .B(n945), .S(n89), .Z(n947) );
  MUX2_X1 U975 ( .A(\REGISTERS[8][23] ), .B(\REGISTERS[24][23] ), .S(n127), 
        .Z(n948) );
  MUX2_X1 U976 ( .A(\REGISTERS[0][23] ), .B(\REGISTERS[16][23] ), .S(n127), 
        .Z(n949) );
  MUX2_X1 U977 ( .A(n949), .B(n948), .S(n89), .Z(n950) );
  MUX2_X1 U978 ( .A(n950), .B(n947), .S(n70), .Z(n951) );
  MUX2_X1 U979 ( .A(n951), .B(n944), .S(ADD_RD2[0]), .Z(n952) );
  MUX2_X1 U980 ( .A(n952), .B(n937), .S(ADD_RD2[1]), .Z(N435) );
  MUX2_X1 U981 ( .A(\REGISTERS[15][24] ), .B(\REGISTERS[31][24] ), .S(n128), 
        .Z(n953) );
  MUX2_X1 U982 ( .A(\REGISTERS[7][24] ), .B(\REGISTERS[23][24] ), .S(n128), 
        .Z(n954) );
  MUX2_X1 U983 ( .A(n954), .B(n953), .S(n90), .Z(n955) );
  MUX2_X1 U984 ( .A(\REGISTERS[11][24] ), .B(\REGISTERS[27][24] ), .S(n128), 
        .Z(n956) );
  MUX2_X1 U985 ( .A(\REGISTERS[3][24] ), .B(\REGISTERS[19][24] ), .S(n128), 
        .Z(n957) );
  MUX2_X1 U986 ( .A(n957), .B(n956), .S(n90), .Z(n958) );
  MUX2_X1 U987 ( .A(n958), .B(n955), .S(n71), .Z(n959) );
  MUX2_X1 U988 ( .A(\REGISTERS[14][24] ), .B(\REGISTERS[30][24] ), .S(n128), 
        .Z(n960) );
  MUX2_X1 U989 ( .A(\REGISTERS[6][24] ), .B(\REGISTERS[22][24] ), .S(n128), 
        .Z(n961) );
  MUX2_X1 U990 ( .A(n961), .B(n960), .S(n90), .Z(n962) );
  MUX2_X1 U991 ( .A(\REGISTERS[10][24] ), .B(\REGISTERS[26][24] ), .S(n128), 
        .Z(n963) );
  MUX2_X1 U992 ( .A(\REGISTERS[2][24] ), .B(\REGISTERS[18][24] ), .S(n128), 
        .Z(n964) );
  MUX2_X1 U993 ( .A(n964), .B(n963), .S(n90), .Z(n965) );
  MUX2_X1 U994 ( .A(n965), .B(n962), .S(n71), .Z(n966) );
  MUX2_X1 U995 ( .A(n966), .B(n959), .S(ADD_RD2[0]), .Z(n967) );
  MUX2_X1 U996 ( .A(\REGISTERS[13][24] ), .B(\REGISTERS[29][24] ), .S(n128), 
        .Z(n968) );
  MUX2_X1 U997 ( .A(\REGISTERS[5][24] ), .B(\REGISTERS[21][24] ), .S(n128), 
        .Z(n969) );
  MUX2_X1 U998 ( .A(n969), .B(n968), .S(n90), .Z(n970) );
  MUX2_X1 U999 ( .A(\REGISTERS[9][24] ), .B(\REGISTERS[25][24] ), .S(n128), 
        .Z(n971) );
  MUX2_X1 U1000 ( .A(\REGISTERS[1][24] ), .B(\REGISTERS[17][24] ), .S(n128), 
        .Z(n972) );
  MUX2_X1 U1001 ( .A(n972), .B(n971), .S(n90), .Z(n973) );
  MUX2_X1 U1002 ( .A(n973), .B(n970), .S(n71), .Z(n974) );
  MUX2_X1 U1003 ( .A(\REGISTERS[12][24] ), .B(\REGISTERS[28][24] ), .S(n129), 
        .Z(n975) );
  MUX2_X1 U1004 ( .A(\REGISTERS[4][24] ), .B(\REGISTERS[20][24] ), .S(n129), 
        .Z(n976) );
  MUX2_X1 U1005 ( .A(n976), .B(n975), .S(n90), .Z(n977) );
  MUX2_X1 U1006 ( .A(\REGISTERS[8][24] ), .B(\REGISTERS[24][24] ), .S(n129), 
        .Z(n978) );
  MUX2_X1 U1007 ( .A(\REGISTERS[0][24] ), .B(\REGISTERS[16][24] ), .S(n129), 
        .Z(n979) );
  MUX2_X1 U1008 ( .A(n979), .B(n978), .S(n90), .Z(n980) );
  MUX2_X1 U1009 ( .A(n980), .B(n977), .S(n71), .Z(n981) );
  MUX2_X1 U1010 ( .A(n981), .B(n974), .S(ADD_RD2[0]), .Z(n982) );
  MUX2_X1 U1011 ( .A(n982), .B(n967), .S(ADD_RD2[1]), .Z(N436) );
  MUX2_X1 U1012 ( .A(\REGISTERS[15][25] ), .B(\REGISTERS[31][25] ), .S(n129), 
        .Z(n983) );
  MUX2_X1 U1013 ( .A(\REGISTERS[7][25] ), .B(\REGISTERS[23][25] ), .S(n129), 
        .Z(n984) );
  MUX2_X1 U1014 ( .A(n984), .B(n983), .S(n90), .Z(n985) );
  MUX2_X1 U1015 ( .A(\REGISTERS[11][25] ), .B(\REGISTERS[27][25] ), .S(n129), 
        .Z(n986) );
  MUX2_X1 U1016 ( .A(\REGISTERS[3][25] ), .B(\REGISTERS[19][25] ), .S(n129), 
        .Z(n987) );
  MUX2_X1 U1017 ( .A(n987), .B(n986), .S(n90), .Z(n988) );
  MUX2_X1 U1018 ( .A(n988), .B(n985), .S(n71), .Z(n989) );
  MUX2_X1 U1019 ( .A(\REGISTERS[14][25] ), .B(\REGISTERS[30][25] ), .S(n129), 
        .Z(n990) );
  MUX2_X1 U1020 ( .A(\REGISTERS[6][25] ), .B(\REGISTERS[22][25] ), .S(n129), 
        .Z(n991) );
  MUX2_X1 U1021 ( .A(n991), .B(n990), .S(n90), .Z(n992) );
  MUX2_X1 U1022 ( .A(\REGISTERS[10][25] ), .B(\REGISTERS[26][25] ), .S(n129), 
        .Z(n993) );
  MUX2_X1 U1023 ( .A(\REGISTERS[2][25] ), .B(\REGISTERS[18][25] ), .S(n129), 
        .Z(n994) );
  MUX2_X1 U1024 ( .A(n994), .B(n993), .S(n90), .Z(n995) );
  MUX2_X1 U1025 ( .A(n995), .B(n992), .S(n71), .Z(n996) );
  MUX2_X1 U1026 ( .A(n996), .B(n989), .S(ADD_RD2[0]), .Z(n997) );
  MUX2_X1 U1027 ( .A(\REGISTERS[13][25] ), .B(\REGISTERS[29][25] ), .S(n130), 
        .Z(n998) );
  MUX2_X1 U1028 ( .A(\REGISTERS[5][25] ), .B(\REGISTERS[21][25] ), .S(n130), 
        .Z(n999) );
  MUX2_X1 U1029 ( .A(n999), .B(n998), .S(n91), .Z(n1000) );
  MUX2_X1 U1030 ( .A(\REGISTERS[9][25] ), .B(\REGISTERS[25][25] ), .S(n130), 
        .Z(n1001) );
  MUX2_X1 U1031 ( .A(\REGISTERS[1][25] ), .B(\REGISTERS[17][25] ), .S(n130), 
        .Z(n1002) );
  MUX2_X1 U1032 ( .A(n1002), .B(n1001), .S(n91), .Z(n1003) );
  MUX2_X1 U1033 ( .A(n1003), .B(n1000), .S(n71), .Z(n1004) );
  MUX2_X1 U1034 ( .A(\REGISTERS[12][25] ), .B(\REGISTERS[28][25] ), .S(n130), 
        .Z(n1005) );
  MUX2_X1 U1035 ( .A(\REGISTERS[4][25] ), .B(\REGISTERS[20][25] ), .S(n130), 
        .Z(n1006) );
  MUX2_X1 U1036 ( .A(n1006), .B(n1005), .S(n91), .Z(n1007) );
  MUX2_X1 U1037 ( .A(\REGISTERS[8][25] ), .B(\REGISTERS[24][25] ), .S(n130), 
        .Z(n1008) );
  MUX2_X1 U1038 ( .A(\REGISTERS[0][25] ), .B(\REGISTERS[16][25] ), .S(n130), 
        .Z(n1009) );
  MUX2_X1 U1039 ( .A(n1009), .B(n1008), .S(n91), .Z(n1010) );
  MUX2_X1 U1040 ( .A(n1010), .B(n1007), .S(n71), .Z(n1011) );
  MUX2_X1 U1041 ( .A(n1011), .B(n1004), .S(ADD_RD2[0]), .Z(n1012) );
  MUX2_X1 U1042 ( .A(n1012), .B(n997), .S(ADD_RD2[1]), .Z(N437) );
  MUX2_X1 U1043 ( .A(\REGISTERS[15][26] ), .B(\REGISTERS[31][26] ), .S(n130), 
        .Z(n1013) );
  MUX2_X1 U1044 ( .A(\REGISTERS[7][26] ), .B(\REGISTERS[23][26] ), .S(n130), 
        .Z(n1014) );
  MUX2_X1 U1045 ( .A(n1014), .B(n1013), .S(n91), .Z(n1015) );
  MUX2_X1 U1046 ( .A(\REGISTERS[11][26] ), .B(\REGISTERS[27][26] ), .S(n130), 
        .Z(n1016) );
  MUX2_X1 U1047 ( .A(\REGISTERS[3][26] ), .B(\REGISTERS[19][26] ), .S(n130), 
        .Z(n1017) );
  MUX2_X1 U1048 ( .A(n1017), .B(n1016), .S(n91), .Z(n1018) );
  MUX2_X1 U1049 ( .A(n1018), .B(n1015), .S(n71), .Z(n1019) );
  MUX2_X1 U1050 ( .A(\REGISTERS[14][26] ), .B(\REGISTERS[30][26] ), .S(n131), 
        .Z(n1020) );
  MUX2_X1 U1051 ( .A(\REGISTERS[6][26] ), .B(\REGISTERS[22][26] ), .S(n131), 
        .Z(n1021) );
  MUX2_X1 U1052 ( .A(n1021), .B(n1020), .S(n91), .Z(n1022) );
  MUX2_X1 U1053 ( .A(\REGISTERS[10][26] ), .B(\REGISTERS[26][26] ), .S(n131), 
        .Z(n1023) );
  MUX2_X1 U1054 ( .A(\REGISTERS[2][26] ), .B(\REGISTERS[18][26] ), .S(n131), 
        .Z(n1024) );
  MUX2_X1 U1055 ( .A(n1024), .B(n1023), .S(n91), .Z(n1025) );
  MUX2_X1 U1056 ( .A(n1025), .B(n1022), .S(n71), .Z(n1026) );
  MUX2_X1 U1057 ( .A(n1026), .B(n1019), .S(ADD_RD2[0]), .Z(n1027) );
  MUX2_X1 U1058 ( .A(\REGISTERS[13][26] ), .B(\REGISTERS[29][26] ), .S(n131), 
        .Z(n1028) );
  MUX2_X1 U1059 ( .A(\REGISTERS[5][26] ), .B(\REGISTERS[21][26] ), .S(n131), 
        .Z(n1029) );
  MUX2_X1 U1060 ( .A(n1029), .B(n1028), .S(n91), .Z(n1030) );
  MUX2_X1 U1061 ( .A(\REGISTERS[9][26] ), .B(\REGISTERS[25][26] ), .S(n131), 
        .Z(n1031) );
  MUX2_X1 U1062 ( .A(\REGISTERS[1][26] ), .B(\REGISTERS[17][26] ), .S(n131), 
        .Z(n1032) );
  MUX2_X1 U1063 ( .A(n1032), .B(n1031), .S(n91), .Z(n1033) );
  MUX2_X1 U1064 ( .A(n1033), .B(n1030), .S(n71), .Z(n1034) );
  MUX2_X1 U1065 ( .A(\REGISTERS[12][26] ), .B(\REGISTERS[28][26] ), .S(n131), 
        .Z(n1035) );
  MUX2_X1 U1066 ( .A(\REGISTERS[4][26] ), .B(\REGISTERS[20][26] ), .S(n131), 
        .Z(n1036) );
  MUX2_X1 U1067 ( .A(n1036), .B(n1035), .S(n91), .Z(n1037) );
  MUX2_X1 U1068 ( .A(\REGISTERS[8][26] ), .B(\REGISTERS[24][26] ), .S(n131), 
        .Z(n1038) );
  MUX2_X1 U1069 ( .A(\REGISTERS[0][26] ), .B(\REGISTERS[16][26] ), .S(n131), 
        .Z(n1039) );
  MUX2_X1 U1070 ( .A(n1039), .B(n1038), .S(n91), .Z(n1040) );
  MUX2_X1 U1071 ( .A(n1040), .B(n1037), .S(n71), .Z(n1041) );
  MUX2_X1 U1072 ( .A(n1041), .B(n1034), .S(ADD_RD2[0]), .Z(n1042) );
  MUX2_X1 U1073 ( .A(n1042), .B(n1027), .S(ADD_RD2[1]), .Z(N438) );
  MUX2_X1 U1074 ( .A(\REGISTERS[15][27] ), .B(\REGISTERS[31][27] ), .S(n132), 
        .Z(n1043) );
  MUX2_X1 U1075 ( .A(\REGISTERS[7][27] ), .B(\REGISTERS[23][27] ), .S(n132), 
        .Z(n1044) );
  MUX2_X1 U1076 ( .A(n1044), .B(n1043), .S(n92), .Z(n1045) );
  MUX2_X1 U1077 ( .A(\REGISTERS[11][27] ), .B(\REGISTERS[27][27] ), .S(n132), 
        .Z(n1046) );
  MUX2_X1 U1078 ( .A(\REGISTERS[3][27] ), .B(\REGISTERS[19][27] ), .S(n132), 
        .Z(n1047) );
  MUX2_X1 U1079 ( .A(n1047), .B(n1046), .S(n92), .Z(n1048) );
  MUX2_X1 U1080 ( .A(n1048), .B(n1045), .S(n72), .Z(n1049) );
  MUX2_X1 U1081 ( .A(\REGISTERS[14][27] ), .B(\REGISTERS[30][27] ), .S(n132), 
        .Z(n1050) );
  MUX2_X1 U1082 ( .A(\REGISTERS[6][27] ), .B(\REGISTERS[22][27] ), .S(n132), 
        .Z(n1051) );
  MUX2_X1 U1083 ( .A(n1051), .B(n1050), .S(n92), .Z(n1052) );
  MUX2_X1 U1084 ( .A(\REGISTERS[10][27] ), .B(\REGISTERS[26][27] ), .S(n132), 
        .Z(n1053) );
  MUX2_X1 U1085 ( .A(\REGISTERS[2][27] ), .B(\REGISTERS[18][27] ), .S(n132), 
        .Z(n1054) );
  MUX2_X1 U1086 ( .A(n1054), .B(n1053), .S(n92), .Z(n1055) );
  MUX2_X1 U1087 ( .A(n1055), .B(n1052), .S(n72), .Z(n1056) );
  MUX2_X1 U1088 ( .A(n1056), .B(n1049), .S(ADD_RD2[0]), .Z(n1057) );
  MUX2_X1 U1089 ( .A(\REGISTERS[13][27] ), .B(\REGISTERS[29][27] ), .S(n132), 
        .Z(n1058) );
  MUX2_X1 U1090 ( .A(\REGISTERS[5][27] ), .B(\REGISTERS[21][27] ), .S(n132), 
        .Z(n1059) );
  MUX2_X1 U1091 ( .A(n1059), .B(n1058), .S(n92), .Z(n1060) );
  MUX2_X1 U1092 ( .A(\REGISTERS[9][27] ), .B(\REGISTERS[25][27] ), .S(n132), 
        .Z(n1061) );
  MUX2_X1 U1093 ( .A(\REGISTERS[1][27] ), .B(\REGISTERS[17][27] ), .S(n132), 
        .Z(n1062) );
  MUX2_X1 U1094 ( .A(n1062), .B(n1061), .S(n92), .Z(n1063) );
  MUX2_X1 U1095 ( .A(n1063), .B(n1060), .S(n72), .Z(n1064) );
  MUX2_X1 U1096 ( .A(\REGISTERS[12][27] ), .B(\REGISTERS[28][27] ), .S(n133), 
        .Z(n1065) );
  MUX2_X1 U1097 ( .A(\REGISTERS[4][27] ), .B(\REGISTERS[20][27] ), .S(n133), 
        .Z(n1066) );
  MUX2_X1 U1098 ( .A(n1066), .B(n1065), .S(n92), .Z(n1067) );
  MUX2_X1 U1099 ( .A(\REGISTERS[8][27] ), .B(\REGISTERS[24][27] ), .S(n133), 
        .Z(n1068) );
  MUX2_X1 U1100 ( .A(\REGISTERS[0][27] ), .B(\REGISTERS[16][27] ), .S(n133), 
        .Z(n1069) );
  MUX2_X1 U1101 ( .A(n1069), .B(n1068), .S(n92), .Z(n1070) );
  MUX2_X1 U1102 ( .A(n1070), .B(n1067), .S(n72), .Z(n1071) );
  MUX2_X1 U1103 ( .A(n1071), .B(n1064), .S(ADD_RD2[0]), .Z(n1072) );
  MUX2_X1 U1104 ( .A(n1072), .B(n1057), .S(ADD_RD2[1]), .Z(N439) );
  MUX2_X1 U1105 ( .A(\REGISTERS[15][28] ), .B(\REGISTERS[31][28] ), .S(n133), 
        .Z(n1073) );
  MUX2_X1 U1106 ( .A(\REGISTERS[7][28] ), .B(\REGISTERS[23][28] ), .S(n133), 
        .Z(n1074) );
  MUX2_X1 U1107 ( .A(n1074), .B(n1073), .S(n92), .Z(n1075) );
  MUX2_X1 U1108 ( .A(\REGISTERS[11][28] ), .B(\REGISTERS[27][28] ), .S(n133), 
        .Z(n1076) );
  MUX2_X1 U1109 ( .A(\REGISTERS[3][28] ), .B(\REGISTERS[19][28] ), .S(n133), 
        .Z(n1077) );
  MUX2_X1 U1110 ( .A(n1077), .B(n1076), .S(n92), .Z(n1078) );
  MUX2_X1 U1111 ( .A(n1078), .B(n1075), .S(n72), .Z(n1079) );
  MUX2_X1 U1112 ( .A(\REGISTERS[14][28] ), .B(\REGISTERS[30][28] ), .S(n133), 
        .Z(n1080) );
  MUX2_X1 U1113 ( .A(\REGISTERS[6][28] ), .B(\REGISTERS[22][28] ), .S(n133), 
        .Z(n1081) );
  MUX2_X1 U1114 ( .A(n1081), .B(n1080), .S(n92), .Z(n1082) );
  MUX2_X1 U1115 ( .A(\REGISTERS[10][28] ), .B(\REGISTERS[26][28] ), .S(n133), 
        .Z(n1083) );
  MUX2_X1 U1116 ( .A(\REGISTERS[2][28] ), .B(\REGISTERS[18][28] ), .S(n133), 
        .Z(n1084) );
  MUX2_X1 U1117 ( .A(n1084), .B(n1083), .S(n92), .Z(n1085) );
  MUX2_X1 U1118 ( .A(n1085), .B(n1082), .S(n72), .Z(n1086) );
  MUX2_X1 U1119 ( .A(n1086), .B(n1079), .S(ADD_RD2[0]), .Z(n1087) );
  MUX2_X1 U1120 ( .A(\REGISTERS[13][28] ), .B(\REGISTERS[29][28] ), .S(n134), 
        .Z(n1088) );
  MUX2_X1 U1121 ( .A(\REGISTERS[5][28] ), .B(\REGISTERS[21][28] ), .S(n134), 
        .Z(n1089) );
  MUX2_X1 U1122 ( .A(n1089), .B(n1088), .S(n93), .Z(n1090) );
  MUX2_X1 U1123 ( .A(\REGISTERS[9][28] ), .B(\REGISTERS[25][28] ), .S(n134), 
        .Z(n1091) );
  MUX2_X1 U1124 ( .A(\REGISTERS[1][28] ), .B(\REGISTERS[17][28] ), .S(n134), 
        .Z(n1092) );
  MUX2_X1 U1125 ( .A(n1092), .B(n1091), .S(n93), .Z(n1093) );
  MUX2_X1 U1126 ( .A(n1093), .B(n1090), .S(n72), .Z(n1094) );
  MUX2_X1 U1127 ( .A(\REGISTERS[12][28] ), .B(\REGISTERS[28][28] ), .S(n134), 
        .Z(n1095) );
  MUX2_X1 U1128 ( .A(\REGISTERS[4][28] ), .B(\REGISTERS[20][28] ), .S(n134), 
        .Z(n1096) );
  MUX2_X1 U1129 ( .A(n1096), .B(n1095), .S(n93), .Z(n1097) );
  MUX2_X1 U1130 ( .A(\REGISTERS[8][28] ), .B(\REGISTERS[24][28] ), .S(n134), 
        .Z(n1098) );
  MUX2_X1 U1131 ( .A(\REGISTERS[0][28] ), .B(\REGISTERS[16][28] ), .S(n134), 
        .Z(n1099) );
  MUX2_X1 U1132 ( .A(n1099), .B(n1098), .S(n93), .Z(n1100) );
  MUX2_X1 U1133 ( .A(n1100), .B(n1097), .S(n72), .Z(n1101) );
  MUX2_X1 U1134 ( .A(n1101), .B(n1094), .S(ADD_RD2[0]), .Z(n1102) );
  MUX2_X1 U1135 ( .A(n1102), .B(n1087), .S(ADD_RD2[1]), .Z(N440) );
  MUX2_X1 U1136 ( .A(\REGISTERS[15][29] ), .B(\REGISTERS[31][29] ), .S(n134), 
        .Z(n1103) );
  MUX2_X1 U1137 ( .A(\REGISTERS[7][29] ), .B(\REGISTERS[23][29] ), .S(n134), 
        .Z(n1104) );
  MUX2_X1 U1138 ( .A(n1104), .B(n1103), .S(n93), .Z(n1105) );
  MUX2_X1 U1139 ( .A(\REGISTERS[11][29] ), .B(\REGISTERS[27][29] ), .S(n134), 
        .Z(n1106) );
  MUX2_X1 U1140 ( .A(\REGISTERS[3][29] ), .B(\REGISTERS[19][29] ), .S(n134), 
        .Z(n1107) );
  MUX2_X1 U1141 ( .A(n1107), .B(n1106), .S(n93), .Z(n1108) );
  MUX2_X1 U1142 ( .A(n1108), .B(n1105), .S(n72), .Z(n1109) );
  MUX2_X1 U1143 ( .A(\REGISTERS[14][29] ), .B(\REGISTERS[30][29] ), .S(n135), 
        .Z(n1110) );
  MUX2_X1 U1144 ( .A(\REGISTERS[6][29] ), .B(\REGISTERS[22][29] ), .S(n135), 
        .Z(n1111) );
  MUX2_X1 U1145 ( .A(n1111), .B(n1110), .S(n93), .Z(n1112) );
  MUX2_X1 U1146 ( .A(\REGISTERS[10][29] ), .B(\REGISTERS[26][29] ), .S(n135), 
        .Z(n1113) );
  MUX2_X1 U1147 ( .A(\REGISTERS[2][29] ), .B(\REGISTERS[18][29] ), .S(n135), 
        .Z(n1114) );
  MUX2_X1 U1148 ( .A(n1114), .B(n1113), .S(n93), .Z(n1115) );
  MUX2_X1 U1149 ( .A(n1115), .B(n1112), .S(n72), .Z(n1116) );
  MUX2_X1 U1150 ( .A(n1116), .B(n1109), .S(ADD_RD2[0]), .Z(n1117) );
  MUX2_X1 U1151 ( .A(\REGISTERS[13][29] ), .B(\REGISTERS[29][29] ), .S(n135), 
        .Z(n1118) );
  MUX2_X1 U1152 ( .A(\REGISTERS[5][29] ), .B(\REGISTERS[21][29] ), .S(n135), 
        .Z(n1119) );
  MUX2_X1 U1153 ( .A(n1119), .B(n1118), .S(n93), .Z(n1120) );
  MUX2_X1 U1154 ( .A(\REGISTERS[9][29] ), .B(\REGISTERS[25][29] ), .S(n135), 
        .Z(n1121) );
  MUX2_X1 U1155 ( .A(\REGISTERS[1][29] ), .B(\REGISTERS[17][29] ), .S(n135), 
        .Z(n1122) );
  MUX2_X1 U1156 ( .A(n1122), .B(n1121), .S(n93), .Z(n1123) );
  MUX2_X1 U1157 ( .A(n1123), .B(n1120), .S(n72), .Z(n1124) );
  MUX2_X1 U1158 ( .A(\REGISTERS[12][29] ), .B(\REGISTERS[28][29] ), .S(n135), 
        .Z(n1125) );
  MUX2_X1 U1159 ( .A(\REGISTERS[4][29] ), .B(\REGISTERS[20][29] ), .S(n135), 
        .Z(n1126) );
  MUX2_X1 U1160 ( .A(n1126), .B(n1125), .S(n93), .Z(n1127) );
  MUX2_X1 U1161 ( .A(\REGISTERS[8][29] ), .B(\REGISTERS[24][29] ), .S(n135), 
        .Z(n1128) );
  MUX2_X1 U1162 ( .A(\REGISTERS[0][29] ), .B(\REGISTERS[16][29] ), .S(n135), 
        .Z(n1129) );
  MUX2_X1 U1163 ( .A(n1129), .B(n1128), .S(n93), .Z(n1130) );
  MUX2_X1 U1164 ( .A(n1130), .B(n1127), .S(n72), .Z(n1131) );
  MUX2_X1 U1165 ( .A(n1131), .B(n1124), .S(ADD_RD2[0]), .Z(n1132) );
  MUX2_X1 U1166 ( .A(n1132), .B(n1117), .S(ADD_RD2[1]), .Z(N441) );
  MUX2_X1 U1167 ( .A(\REGISTERS[15][30] ), .B(\REGISTERS[31][30] ), .S(n136), 
        .Z(n1133) );
  MUX2_X1 U1168 ( .A(\REGISTERS[7][30] ), .B(\REGISTERS[23][30] ), .S(n136), 
        .Z(n1134) );
  MUX2_X1 U1169 ( .A(n1134), .B(n1133), .S(n94), .Z(n1135) );
  MUX2_X1 U1170 ( .A(\REGISTERS[11][30] ), .B(\REGISTERS[27][30] ), .S(n136), 
        .Z(n1136) );
  MUX2_X1 U1171 ( .A(\REGISTERS[3][30] ), .B(\REGISTERS[19][30] ), .S(n136), 
        .Z(n1137) );
  MUX2_X1 U1172 ( .A(n1137), .B(n1136), .S(n94), .Z(n1138) );
  MUX2_X1 U1173 ( .A(n1138), .B(n1135), .S(n73), .Z(n1139) );
  MUX2_X1 U1174 ( .A(\REGISTERS[14][30] ), .B(\REGISTERS[30][30] ), .S(n136), 
        .Z(n2164) );
  MUX2_X1 U1175 ( .A(\REGISTERS[6][30] ), .B(\REGISTERS[22][30] ), .S(n136), 
        .Z(n2165) );
  MUX2_X1 U1176 ( .A(n2165), .B(n2164), .S(n94), .Z(n2166) );
  MUX2_X1 U1177 ( .A(\REGISTERS[10][30] ), .B(\REGISTERS[26][30] ), .S(n136), 
        .Z(n2167) );
  MUX2_X1 U1178 ( .A(\REGISTERS[2][30] ), .B(\REGISTERS[18][30] ), .S(n136), 
        .Z(n2168) );
  MUX2_X1 U1179 ( .A(n2168), .B(n2167), .S(n94), .Z(n2169) );
  MUX2_X1 U1180 ( .A(n2169), .B(n2166), .S(n73), .Z(n2170) );
  MUX2_X1 U1181 ( .A(n2170), .B(n1139), .S(ADD_RD2[0]), .Z(n2171) );
  MUX2_X1 U1182 ( .A(\REGISTERS[13][30] ), .B(\REGISTERS[29][30] ), .S(n136), 
        .Z(n2172) );
  MUX2_X1 U1183 ( .A(\REGISTERS[5][30] ), .B(\REGISTERS[21][30] ), .S(n136), 
        .Z(n2173) );
  MUX2_X1 U1184 ( .A(n2173), .B(n2172), .S(n94), .Z(n2174) );
  MUX2_X1 U1185 ( .A(\REGISTERS[9][30] ), .B(\REGISTERS[25][30] ), .S(n136), 
        .Z(n2175) );
  MUX2_X1 U1186 ( .A(\REGISTERS[1][30] ), .B(\REGISTERS[17][30] ), .S(n136), 
        .Z(n2176) );
  MUX2_X1 U1187 ( .A(n2176), .B(n2175), .S(n94), .Z(n2177) );
  MUX2_X1 U1188 ( .A(n2177), .B(n2174), .S(n73), .Z(n2178) );
  MUX2_X1 U1189 ( .A(\REGISTERS[12][30] ), .B(\REGISTERS[28][30] ), .S(n137), 
        .Z(n2179) );
  MUX2_X1 U1190 ( .A(\REGISTERS[4][30] ), .B(\REGISTERS[20][30] ), .S(n137), 
        .Z(n2180) );
  MUX2_X1 U1191 ( .A(n2180), .B(n2179), .S(n94), .Z(n2181) );
  MUX2_X1 U1192 ( .A(\REGISTERS[8][30] ), .B(\REGISTERS[24][30] ), .S(n137), 
        .Z(n2182) );
  MUX2_X1 U1193 ( .A(\REGISTERS[0][30] ), .B(\REGISTERS[16][30] ), .S(n137), 
        .Z(n2183) );
  MUX2_X1 U1194 ( .A(n2183), .B(n2182), .S(n94), .Z(n2184) );
  MUX2_X1 U1195 ( .A(n2184), .B(n2181), .S(n73), .Z(n2185) );
  MUX2_X1 U1196 ( .A(n2185), .B(n2178), .S(ADD_RD2[0]), .Z(n2186) );
  MUX2_X1 U1197 ( .A(n2186), .B(n2171), .S(ADD_RD2[1]), .Z(N442) );
  MUX2_X1 U1198 ( .A(\REGISTERS[15][31] ), .B(\REGISTERS[31][31] ), .S(n137), 
        .Z(n2187) );
  MUX2_X1 U1199 ( .A(\REGISTERS[7][31] ), .B(\REGISTERS[23][31] ), .S(n137), 
        .Z(n2188) );
  MUX2_X1 U1200 ( .A(n2188), .B(n2187), .S(n94), .Z(n2189) );
  MUX2_X1 U1201 ( .A(\REGISTERS[11][31] ), .B(\REGISTERS[27][31] ), .S(n137), 
        .Z(n2190) );
  MUX2_X1 U1202 ( .A(\REGISTERS[3][31] ), .B(\REGISTERS[19][31] ), .S(n137), 
        .Z(n2191) );
  MUX2_X1 U1203 ( .A(n2191), .B(n2190), .S(n94), .Z(n2192) );
  MUX2_X1 U1204 ( .A(n2192), .B(n2189), .S(n73), .Z(n2193) );
  MUX2_X1 U1205 ( .A(\REGISTERS[14][31] ), .B(\REGISTERS[30][31] ), .S(n137), 
        .Z(n2194) );
  MUX2_X1 U1206 ( .A(\REGISTERS[6][31] ), .B(\REGISTERS[22][31] ), .S(n137), 
        .Z(n2195) );
  MUX2_X1 U1207 ( .A(n2195), .B(n2194), .S(n94), .Z(n2196) );
  MUX2_X1 U1208 ( .A(\REGISTERS[10][31] ), .B(\REGISTERS[26][31] ), .S(n137), 
        .Z(n2197) );
  MUX2_X1 U1209 ( .A(\REGISTERS[2][31] ), .B(\REGISTERS[18][31] ), .S(n137), 
        .Z(n2198) );
  MUX2_X1 U1210 ( .A(n2198), .B(n2197), .S(n94), .Z(n2199) );
  MUX2_X1 U1211 ( .A(n2199), .B(n2196), .S(n73), .Z(n2200) );
  MUX2_X1 U1212 ( .A(n2200), .B(n2193), .S(ADD_RD2[0]), .Z(n2201) );
  MUX2_X1 U1213 ( .A(\REGISTERS[13][31] ), .B(\REGISTERS[29][31] ), .S(n138), 
        .Z(n2202) );
  MUX2_X1 U1214 ( .A(\REGISTERS[5][31] ), .B(\REGISTERS[21][31] ), .S(n138), 
        .Z(n2203) );
  MUX2_X1 U1215 ( .A(n2203), .B(n2202), .S(n95), .Z(n2204) );
  MUX2_X1 U1216 ( .A(\REGISTERS[9][31] ), .B(\REGISTERS[25][31] ), .S(n138), 
        .Z(n2205) );
  MUX2_X1 U1217 ( .A(\REGISTERS[1][31] ), .B(\REGISTERS[17][31] ), .S(n138), 
        .Z(n2206) );
  MUX2_X1 U1218 ( .A(n2206), .B(n2205), .S(n95), .Z(n2207) );
  MUX2_X1 U1219 ( .A(n2207), .B(n2204), .S(n73), .Z(n2208) );
  MUX2_X1 U1220 ( .A(\REGISTERS[12][31] ), .B(\REGISTERS[28][31] ), .S(n138), 
        .Z(n2209) );
  MUX2_X1 U1221 ( .A(\REGISTERS[4][31] ), .B(\REGISTERS[20][31] ), .S(n138), 
        .Z(n2210) );
  MUX2_X1 U1222 ( .A(n2210), .B(n2209), .S(n95), .Z(n2211) );
  MUX2_X1 U1223 ( .A(\REGISTERS[8][31] ), .B(\REGISTERS[24][31] ), .S(n138), 
        .Z(n2212) );
  MUX2_X1 U1224 ( .A(\REGISTERS[0][31] ), .B(\REGISTERS[16][31] ), .S(n138), 
        .Z(n2213) );
  MUX2_X1 U1225 ( .A(n2213), .B(n2212), .S(n95), .Z(n2214) );
  MUX2_X1 U1226 ( .A(n2214), .B(n2211), .S(n73), .Z(n2215) );
  MUX2_X1 U1227 ( .A(n2215), .B(n2208), .S(ADD_RD2[0]), .Z(n2216) );
  MUX2_X1 U1228 ( .A(n2216), .B(n2201), .S(ADD_RD2[1]), .Z(N443) );
  MUX2_X1 U1229 ( .A(\REGISTERS[15][0] ), .B(\REGISTERS[31][0] ), .S(n181), 
        .Z(n2217) );
  MUX2_X1 U1230 ( .A(\REGISTERS[7][0] ), .B(\REGISTERS[23][0] ), .S(n181), .Z(
        n2218) );
  MUX2_X1 U1231 ( .A(n2218), .B(n2217), .S(n159), .Z(n2219) );
  MUX2_X1 U1232 ( .A(\REGISTERS[11][0] ), .B(\REGISTERS[27][0] ), .S(n181), 
        .Z(n2220) );
  MUX2_X1 U1233 ( .A(\REGISTERS[3][0] ), .B(\REGISTERS[19][0] ), .S(n181), .Z(
        n2221) );
  MUX2_X1 U1234 ( .A(n2221), .B(n2220), .S(n159), .Z(n2222) );
  MUX2_X1 U1235 ( .A(n2222), .B(n2219), .S(n148), .Z(n2223) );
  MUX2_X1 U1236 ( .A(\REGISTERS[14][0] ), .B(\REGISTERS[30][0] ), .S(n181), 
        .Z(n2224) );
  MUX2_X1 U1237 ( .A(\REGISTERS[6][0] ), .B(\REGISTERS[22][0] ), .S(n181), .Z(
        n2225) );
  MUX2_X1 U1238 ( .A(n2225), .B(n2224), .S(n159), .Z(n2226) );
  MUX2_X1 U1239 ( .A(\REGISTERS[10][0] ), .B(\REGISTERS[26][0] ), .S(n181), 
        .Z(n2227) );
  MUX2_X1 U1240 ( .A(\REGISTERS[2][0] ), .B(\REGISTERS[18][0] ), .S(n181), .Z(
        n2228) );
  MUX2_X1 U1241 ( .A(n2228), .B(n2227), .S(n159), .Z(n2229) );
  MUX2_X1 U1242 ( .A(n2229), .B(n2226), .S(n148), .Z(n2230) );
  MUX2_X1 U1243 ( .A(n2230), .B(n2223), .S(ADD_RD1[0]), .Z(n2231) );
  MUX2_X1 U1244 ( .A(\REGISTERS[13][0] ), .B(\REGISTERS[29][0] ), .S(n181), 
        .Z(n2232) );
  MUX2_X1 U1245 ( .A(\REGISTERS[5][0] ), .B(\REGISTERS[21][0] ), .S(n181), .Z(
        n2233) );
  MUX2_X1 U1246 ( .A(n2233), .B(n2232), .S(n159), .Z(n2234) );
  MUX2_X1 U1247 ( .A(\REGISTERS[9][0] ), .B(\REGISTERS[25][0] ), .S(n181), .Z(
        n2235) );
  MUX2_X1 U1248 ( .A(\REGISTERS[1][0] ), .B(\REGISTERS[17][0] ), .S(n181), .Z(
        n2236) );
  MUX2_X1 U1249 ( .A(n2236), .B(n2235), .S(n159), .Z(n2237) );
  MUX2_X1 U1250 ( .A(n2237), .B(n2234), .S(n148), .Z(n2238) );
  MUX2_X1 U1251 ( .A(\REGISTERS[12][0] ), .B(\REGISTERS[28][0] ), .S(n182), 
        .Z(n2239) );
  MUX2_X1 U1252 ( .A(\REGISTERS[4][0] ), .B(\REGISTERS[20][0] ), .S(n182), .Z(
        n2240) );
  MUX2_X1 U1253 ( .A(n2240), .B(n2239), .S(n159), .Z(n2241) );
  MUX2_X1 U1254 ( .A(\REGISTERS[8][0] ), .B(\REGISTERS[24][0] ), .S(n182), .Z(
        n2242) );
  MUX2_X1 U1255 ( .A(\REGISTERS[0][0] ), .B(\REGISTERS[16][0] ), .S(n182), .Z(
        n2243) );
  MUX2_X1 U1256 ( .A(n2243), .B(n2242), .S(n159), .Z(n2244) );
  MUX2_X1 U1257 ( .A(n2244), .B(n2241), .S(n148), .Z(n2245) );
  MUX2_X1 U1258 ( .A(n2245), .B(n2238), .S(ADD_RD1[0]), .Z(n2246) );
  MUX2_X1 U1259 ( .A(n2246), .B(n2231), .S(ADD_RD1[1]), .Z(N379) );
  MUX2_X1 U1260 ( .A(\REGISTERS[15][1] ), .B(\REGISTERS[31][1] ), .S(n182), 
        .Z(n2247) );
  MUX2_X1 U1261 ( .A(\REGISTERS[7][1] ), .B(\REGISTERS[23][1] ), .S(n182), .Z(
        n2248) );
  MUX2_X1 U1262 ( .A(n2248), .B(n2247), .S(n159), .Z(n2249) );
  MUX2_X1 U1263 ( .A(\REGISTERS[11][1] ), .B(\REGISTERS[27][1] ), .S(n182), 
        .Z(n2250) );
  MUX2_X1 U1264 ( .A(\REGISTERS[3][1] ), .B(\REGISTERS[19][1] ), .S(n182), .Z(
        n2251) );
  MUX2_X1 U1265 ( .A(n2251), .B(n2250), .S(n159), .Z(n2252) );
  MUX2_X1 U1266 ( .A(n2252), .B(n2249), .S(n148), .Z(n2253) );
  MUX2_X1 U1267 ( .A(\REGISTERS[14][1] ), .B(\REGISTERS[30][1] ), .S(n182), 
        .Z(n2254) );
  MUX2_X1 U1268 ( .A(\REGISTERS[6][1] ), .B(\REGISTERS[22][1] ), .S(n182), .Z(
        n2255) );
  MUX2_X1 U1269 ( .A(n2255), .B(n2254), .S(n159), .Z(n2256) );
  MUX2_X1 U1270 ( .A(\REGISTERS[10][1] ), .B(\REGISTERS[26][1] ), .S(n182), 
        .Z(n2257) );
  MUX2_X1 U1271 ( .A(\REGISTERS[2][1] ), .B(\REGISTERS[18][1] ), .S(n182), .Z(
        n2258) );
  MUX2_X1 U1272 ( .A(n2258), .B(n2257), .S(n159), .Z(n2259) );
  MUX2_X1 U1273 ( .A(n2259), .B(n2256), .S(n148), .Z(n2260) );
  MUX2_X1 U1274 ( .A(n2260), .B(n2253), .S(ADD_RD1[0]), .Z(n2261) );
  MUX2_X1 U1275 ( .A(\REGISTERS[13][1] ), .B(\REGISTERS[29][1] ), .S(n183), 
        .Z(n2262) );
  MUX2_X1 U1276 ( .A(\REGISTERS[5][1] ), .B(\REGISTERS[21][1] ), .S(n183), .Z(
        n2263) );
  MUX2_X1 U1277 ( .A(n2263), .B(n2262), .S(n160), .Z(n2264) );
  MUX2_X1 U1278 ( .A(\REGISTERS[9][1] ), .B(\REGISTERS[25][1] ), .S(n183), .Z(
        n2265) );
  MUX2_X1 U1279 ( .A(\REGISTERS[1][1] ), .B(\REGISTERS[17][1] ), .S(n183), .Z(
        n2266) );
  MUX2_X1 U1280 ( .A(n2266), .B(n2265), .S(n160), .Z(n2267) );
  MUX2_X1 U1281 ( .A(n2267), .B(n2264), .S(n148), .Z(n2268) );
  MUX2_X1 U1282 ( .A(\REGISTERS[12][1] ), .B(\REGISTERS[28][1] ), .S(n183), 
        .Z(n2269) );
  MUX2_X1 U1283 ( .A(\REGISTERS[4][1] ), .B(\REGISTERS[20][1] ), .S(n183), .Z(
        n2270) );
  MUX2_X1 U1284 ( .A(n2270), .B(n2269), .S(n160), .Z(n2271) );
  MUX2_X1 U1285 ( .A(\REGISTERS[8][1] ), .B(\REGISTERS[24][1] ), .S(n183), .Z(
        n2272) );
  MUX2_X1 U1286 ( .A(\REGISTERS[0][1] ), .B(\REGISTERS[16][1] ), .S(n183), .Z(
        n2273) );
  MUX2_X1 U1287 ( .A(n2273), .B(n2272), .S(n160), .Z(n2274) );
  MUX2_X1 U1288 ( .A(n2274), .B(n2271), .S(n148), .Z(n2275) );
  MUX2_X1 U1289 ( .A(n2275), .B(n2268), .S(ADD_RD1[0]), .Z(n2276) );
  MUX2_X1 U1290 ( .A(n2276), .B(n2261), .S(ADD_RD1[1]), .Z(N380) );
  MUX2_X1 U1291 ( .A(\REGISTERS[15][2] ), .B(\REGISTERS[31][2] ), .S(n183), 
        .Z(n2277) );
  MUX2_X1 U1292 ( .A(\REGISTERS[7][2] ), .B(\REGISTERS[23][2] ), .S(n183), .Z(
        n2278) );
  MUX2_X1 U1293 ( .A(n2278), .B(n2277), .S(n160), .Z(n2279) );
  MUX2_X1 U1294 ( .A(\REGISTERS[11][2] ), .B(\REGISTERS[27][2] ), .S(n183), 
        .Z(n2280) );
  MUX2_X1 U1295 ( .A(\REGISTERS[3][2] ), .B(\REGISTERS[19][2] ), .S(n183), .Z(
        n2281) );
  MUX2_X1 U1296 ( .A(n2281), .B(n2280), .S(n160), .Z(n2282) );
  MUX2_X1 U1297 ( .A(n2282), .B(n2279), .S(n148), .Z(n2283) );
  MUX2_X1 U1298 ( .A(\REGISTERS[14][2] ), .B(\REGISTERS[30][2] ), .S(n184), 
        .Z(n2284) );
  MUX2_X1 U1299 ( .A(\REGISTERS[6][2] ), .B(\REGISTERS[22][2] ), .S(n184), .Z(
        n2285) );
  MUX2_X1 U1300 ( .A(n2285), .B(n2284), .S(n160), .Z(n2286) );
  MUX2_X1 U1301 ( .A(\REGISTERS[10][2] ), .B(\REGISTERS[26][2] ), .S(n184), 
        .Z(n2287) );
  MUX2_X1 U1302 ( .A(\REGISTERS[2][2] ), .B(\REGISTERS[18][2] ), .S(n184), .Z(
        n2288) );
  MUX2_X1 U1303 ( .A(n2288), .B(n2287), .S(n160), .Z(n2289) );
  MUX2_X1 U1304 ( .A(n2289), .B(n2286), .S(n148), .Z(n2290) );
  MUX2_X1 U1305 ( .A(n2290), .B(n2283), .S(ADD_RD1[0]), .Z(n2291) );
  MUX2_X1 U1306 ( .A(\REGISTERS[13][2] ), .B(\REGISTERS[29][2] ), .S(n184), 
        .Z(n2292) );
  MUX2_X1 U1307 ( .A(\REGISTERS[5][2] ), .B(\REGISTERS[21][2] ), .S(n184), .Z(
        n2293) );
  MUX2_X1 U1308 ( .A(n2293), .B(n2292), .S(n160), .Z(n2294) );
  MUX2_X1 U1309 ( .A(\REGISTERS[9][2] ), .B(\REGISTERS[25][2] ), .S(n184), .Z(
        n2295) );
  MUX2_X1 U1310 ( .A(\REGISTERS[1][2] ), .B(\REGISTERS[17][2] ), .S(n184), .Z(
        n2296) );
  MUX2_X1 U1311 ( .A(n2296), .B(n2295), .S(n160), .Z(n2297) );
  MUX2_X1 U1312 ( .A(n2297), .B(n2294), .S(n148), .Z(n2298) );
  MUX2_X1 U1313 ( .A(\REGISTERS[12][2] ), .B(\REGISTERS[28][2] ), .S(n184), 
        .Z(n2299) );
  MUX2_X1 U1314 ( .A(\REGISTERS[4][2] ), .B(\REGISTERS[20][2] ), .S(n184), .Z(
        n2300) );
  MUX2_X1 U1315 ( .A(n2300), .B(n2299), .S(n160), .Z(n2301) );
  MUX2_X1 U1316 ( .A(\REGISTERS[8][2] ), .B(\REGISTERS[24][2] ), .S(n184), .Z(
        n2302) );
  MUX2_X1 U1317 ( .A(\REGISTERS[0][2] ), .B(\REGISTERS[16][2] ), .S(n184), .Z(
        n2303) );
  MUX2_X1 U1318 ( .A(n2303), .B(n2302), .S(n160), .Z(n2304) );
  MUX2_X1 U1319 ( .A(n2304), .B(n2301), .S(n148), .Z(n2305) );
  MUX2_X1 U1320 ( .A(n2305), .B(n2298), .S(ADD_RD1[0]), .Z(n2306) );
  MUX2_X1 U1321 ( .A(n2306), .B(n2291), .S(ADD_RD1[1]), .Z(N381) );
  MUX2_X1 U1322 ( .A(\REGISTERS[15][3] ), .B(\REGISTERS[31][3] ), .S(n185), 
        .Z(n2307) );
  MUX2_X1 U1323 ( .A(\REGISTERS[7][3] ), .B(\REGISTERS[23][3] ), .S(n185), .Z(
        n2308) );
  MUX2_X1 U1324 ( .A(n2308), .B(n2307), .S(n161), .Z(n2309) );
  MUX2_X1 U1325 ( .A(\REGISTERS[11][3] ), .B(\REGISTERS[27][3] ), .S(n185), 
        .Z(n2310) );
  MUX2_X1 U1326 ( .A(\REGISTERS[3][3] ), .B(\REGISTERS[19][3] ), .S(n185), .Z(
        n2311) );
  MUX2_X1 U1327 ( .A(n2311), .B(n2310), .S(n161), .Z(n2312) );
  MUX2_X1 U1328 ( .A(n2312), .B(n2309), .S(n149), .Z(n2313) );
  MUX2_X1 U1329 ( .A(\REGISTERS[14][3] ), .B(\REGISTERS[30][3] ), .S(n185), 
        .Z(n2314) );
  MUX2_X1 U1330 ( .A(\REGISTERS[6][3] ), .B(\REGISTERS[22][3] ), .S(n185), .Z(
        n2315) );
  MUX2_X1 U1331 ( .A(n2315), .B(n2314), .S(n161), .Z(n2316) );
  MUX2_X1 U1332 ( .A(\REGISTERS[10][3] ), .B(\REGISTERS[26][3] ), .S(n185), 
        .Z(n2317) );
  MUX2_X1 U1333 ( .A(\REGISTERS[2][3] ), .B(\REGISTERS[18][3] ), .S(n185), .Z(
        n2318) );
  MUX2_X1 U1334 ( .A(n2318), .B(n2317), .S(n161), .Z(n2319) );
  MUX2_X1 U1335 ( .A(n2319), .B(n2316), .S(n149), .Z(n2320) );
  MUX2_X1 U1336 ( .A(n2320), .B(n2313), .S(ADD_RD1[0]), .Z(n2321) );
  MUX2_X1 U1337 ( .A(\REGISTERS[13][3] ), .B(\REGISTERS[29][3] ), .S(n185), 
        .Z(n2322) );
  MUX2_X1 U1338 ( .A(\REGISTERS[5][3] ), .B(\REGISTERS[21][3] ), .S(n185), .Z(
        n2323) );
  MUX2_X1 U1339 ( .A(n2323), .B(n2322), .S(n161), .Z(n2324) );
  MUX2_X1 U1340 ( .A(\REGISTERS[9][3] ), .B(\REGISTERS[25][3] ), .S(n185), .Z(
        n2325) );
  MUX2_X1 U1341 ( .A(\REGISTERS[1][3] ), .B(\REGISTERS[17][3] ), .S(n185), .Z(
        n2326) );
  MUX2_X1 U1342 ( .A(n2326), .B(n2325), .S(n161), .Z(n2327) );
  MUX2_X1 U1343 ( .A(n2327), .B(n2324), .S(n149), .Z(n2328) );
  MUX2_X1 U1344 ( .A(\REGISTERS[12][3] ), .B(\REGISTERS[28][3] ), .S(n186), 
        .Z(n2329) );
  MUX2_X1 U1345 ( .A(\REGISTERS[4][3] ), .B(\REGISTERS[20][3] ), .S(n186), .Z(
        n2330) );
  MUX2_X1 U1346 ( .A(n2330), .B(n2329), .S(n161), .Z(n2331) );
  MUX2_X1 U1347 ( .A(\REGISTERS[8][3] ), .B(\REGISTERS[24][3] ), .S(n186), .Z(
        n2332) );
  MUX2_X1 U1348 ( .A(\REGISTERS[0][3] ), .B(\REGISTERS[16][3] ), .S(n186), .Z(
        n2333) );
  MUX2_X1 U1349 ( .A(n2333), .B(n2332), .S(n161), .Z(n2334) );
  MUX2_X1 U1350 ( .A(n2334), .B(n2331), .S(n149), .Z(n2335) );
  MUX2_X1 U1351 ( .A(n2335), .B(n2328), .S(ADD_RD1[0]), .Z(n2336) );
  MUX2_X1 U1352 ( .A(n2336), .B(n2321), .S(ADD_RD1[1]), .Z(N382) );
  MUX2_X1 U1353 ( .A(\REGISTERS[15][4] ), .B(\REGISTERS[31][4] ), .S(n186), 
        .Z(n2337) );
  MUX2_X1 U1354 ( .A(\REGISTERS[7][4] ), .B(\REGISTERS[23][4] ), .S(n186), .Z(
        n2338) );
  MUX2_X1 U1355 ( .A(n2338), .B(n2337), .S(n161), .Z(n2339) );
  MUX2_X1 U1356 ( .A(\REGISTERS[11][4] ), .B(\REGISTERS[27][4] ), .S(n186), 
        .Z(n2340) );
  MUX2_X1 U1357 ( .A(\REGISTERS[3][4] ), .B(\REGISTERS[19][4] ), .S(n186), .Z(
        n2341) );
  MUX2_X1 U1358 ( .A(n2341), .B(n2340), .S(n161), .Z(n2342) );
  MUX2_X1 U1359 ( .A(n2342), .B(n2339), .S(n149), .Z(n2343) );
  MUX2_X1 U1360 ( .A(\REGISTERS[14][4] ), .B(\REGISTERS[30][4] ), .S(n186), 
        .Z(n2344) );
  MUX2_X1 U1361 ( .A(\REGISTERS[6][4] ), .B(\REGISTERS[22][4] ), .S(n186), .Z(
        n2345) );
  MUX2_X1 U1362 ( .A(n2345), .B(n2344), .S(n161), .Z(n2346) );
  MUX2_X1 U1363 ( .A(\REGISTERS[10][4] ), .B(\REGISTERS[26][4] ), .S(n186), 
        .Z(n2347) );
  MUX2_X1 U1364 ( .A(\REGISTERS[2][4] ), .B(\REGISTERS[18][4] ), .S(n186), .Z(
        n2348) );
  MUX2_X1 U1365 ( .A(n2348), .B(n2347), .S(n161), .Z(n2349) );
  MUX2_X1 U1366 ( .A(n2349), .B(n2346), .S(n149), .Z(n2350) );
  MUX2_X1 U1367 ( .A(n2350), .B(n2343), .S(ADD_RD1[0]), .Z(n2351) );
  MUX2_X1 U1368 ( .A(\REGISTERS[13][4] ), .B(\REGISTERS[29][4] ), .S(n187), 
        .Z(n2352) );
  MUX2_X1 U1369 ( .A(\REGISTERS[5][4] ), .B(\REGISTERS[21][4] ), .S(n187), .Z(
        n2353) );
  MUX2_X1 U1370 ( .A(n2353), .B(n2352), .S(n162), .Z(n2354) );
  MUX2_X1 U1371 ( .A(\REGISTERS[9][4] ), .B(\REGISTERS[25][4] ), .S(n187), .Z(
        n2355) );
  MUX2_X1 U1372 ( .A(\REGISTERS[1][4] ), .B(\REGISTERS[17][4] ), .S(n187), .Z(
        n2356) );
  MUX2_X1 U1373 ( .A(n2356), .B(n2355), .S(n162), .Z(n2357) );
  MUX2_X1 U1374 ( .A(n2357), .B(n2354), .S(n149), .Z(n2358) );
  MUX2_X1 U1375 ( .A(\REGISTERS[12][4] ), .B(\REGISTERS[28][4] ), .S(n187), 
        .Z(n2359) );
  MUX2_X1 U1376 ( .A(\REGISTERS[4][4] ), .B(\REGISTERS[20][4] ), .S(n187), .Z(
        n2360) );
  MUX2_X1 U1377 ( .A(n2360), .B(n2359), .S(n162), .Z(n2361) );
  MUX2_X1 U1378 ( .A(\REGISTERS[8][4] ), .B(\REGISTERS[24][4] ), .S(n187), .Z(
        n2362) );
  MUX2_X1 U1379 ( .A(\REGISTERS[0][4] ), .B(\REGISTERS[16][4] ), .S(n187), .Z(
        n2363) );
  MUX2_X1 U1380 ( .A(n2363), .B(n2362), .S(n162), .Z(n2364) );
  MUX2_X1 U1381 ( .A(n2364), .B(n2361), .S(n149), .Z(n2365) );
  MUX2_X1 U1382 ( .A(n2365), .B(n2358), .S(ADD_RD1[0]), .Z(n2366) );
  MUX2_X1 U1383 ( .A(n2366), .B(n2351), .S(ADD_RD1[1]), .Z(N383) );
  MUX2_X1 U1384 ( .A(\REGISTERS[15][5] ), .B(\REGISTERS[31][5] ), .S(n187), 
        .Z(n2367) );
  MUX2_X1 U1385 ( .A(\REGISTERS[7][5] ), .B(\REGISTERS[23][5] ), .S(n187), .Z(
        n2368) );
  MUX2_X1 U1386 ( .A(n2368), .B(n2367), .S(n162), .Z(n2369) );
  MUX2_X1 U1387 ( .A(\REGISTERS[11][5] ), .B(\REGISTERS[27][5] ), .S(n187), 
        .Z(n2370) );
  MUX2_X1 U1388 ( .A(\REGISTERS[3][5] ), .B(\REGISTERS[19][5] ), .S(n187), .Z(
        n2371) );
  MUX2_X1 U1389 ( .A(n2371), .B(n2370), .S(n162), .Z(n2372) );
  MUX2_X1 U1390 ( .A(n2372), .B(n2369), .S(n149), .Z(n2373) );
  MUX2_X1 U1391 ( .A(\REGISTERS[14][5] ), .B(\REGISTERS[30][5] ), .S(n188), 
        .Z(n2374) );
  MUX2_X1 U1392 ( .A(\REGISTERS[6][5] ), .B(\REGISTERS[22][5] ), .S(n188), .Z(
        n2375) );
  MUX2_X1 U1393 ( .A(n2375), .B(n2374), .S(n162), .Z(n2376) );
  MUX2_X1 U1394 ( .A(\REGISTERS[10][5] ), .B(\REGISTERS[26][5] ), .S(n188), 
        .Z(n2377) );
  MUX2_X1 U1395 ( .A(\REGISTERS[2][5] ), .B(\REGISTERS[18][5] ), .S(n188), .Z(
        n2378) );
  MUX2_X1 U1396 ( .A(n2378), .B(n2377), .S(n162), .Z(n2379) );
  MUX2_X1 U1397 ( .A(n2379), .B(n2376), .S(n149), .Z(n2380) );
  MUX2_X1 U1398 ( .A(n2380), .B(n2373), .S(ADD_RD1[0]), .Z(n2381) );
  MUX2_X1 U1399 ( .A(\REGISTERS[13][5] ), .B(\REGISTERS[29][5] ), .S(n188), 
        .Z(n2382) );
  MUX2_X1 U1400 ( .A(\REGISTERS[5][5] ), .B(\REGISTERS[21][5] ), .S(n188), .Z(
        n2383) );
  MUX2_X1 U1401 ( .A(n2383), .B(n2382), .S(n162), .Z(n2384) );
  MUX2_X1 U1402 ( .A(\REGISTERS[9][5] ), .B(\REGISTERS[25][5] ), .S(n188), .Z(
        n2385) );
  MUX2_X1 U1403 ( .A(\REGISTERS[1][5] ), .B(\REGISTERS[17][5] ), .S(n188), .Z(
        n2386) );
  MUX2_X1 U1404 ( .A(n2386), .B(n2385), .S(n162), .Z(n2387) );
  MUX2_X1 U1405 ( .A(n2387), .B(n2384), .S(n149), .Z(n2388) );
  MUX2_X1 U1406 ( .A(\REGISTERS[12][5] ), .B(\REGISTERS[28][5] ), .S(n188), 
        .Z(n2389) );
  MUX2_X1 U1407 ( .A(\REGISTERS[4][5] ), .B(\REGISTERS[20][5] ), .S(n188), .Z(
        n2390) );
  MUX2_X1 U1408 ( .A(n2390), .B(n2389), .S(n162), .Z(n2391) );
  MUX2_X1 U1409 ( .A(\REGISTERS[8][5] ), .B(\REGISTERS[24][5] ), .S(n188), .Z(
        n2392) );
  MUX2_X1 U1410 ( .A(\REGISTERS[0][5] ), .B(\REGISTERS[16][5] ), .S(n188), .Z(
        n2393) );
  MUX2_X1 U1411 ( .A(n2393), .B(n2392), .S(n162), .Z(n2394) );
  MUX2_X1 U1412 ( .A(n2394), .B(n2391), .S(n149), .Z(n2395) );
  MUX2_X1 U1413 ( .A(n2395), .B(n2388), .S(ADD_RD1[0]), .Z(n2396) );
  MUX2_X1 U1414 ( .A(n2396), .B(n2381), .S(ADD_RD1[1]), .Z(N384) );
  MUX2_X1 U1415 ( .A(\REGISTERS[15][6] ), .B(\REGISTERS[31][6] ), .S(n189), 
        .Z(n2397) );
  MUX2_X1 U1416 ( .A(\REGISTERS[7][6] ), .B(\REGISTERS[23][6] ), .S(n189), .Z(
        n2398) );
  MUX2_X1 U1417 ( .A(n2398), .B(n2397), .S(n163), .Z(n2399) );
  MUX2_X1 U1418 ( .A(\REGISTERS[11][6] ), .B(\REGISTERS[27][6] ), .S(n189), 
        .Z(n2400) );
  MUX2_X1 U1419 ( .A(\REGISTERS[3][6] ), .B(\REGISTERS[19][6] ), .S(n189), .Z(
        n2401) );
  MUX2_X1 U1420 ( .A(n2401), .B(n2400), .S(n163), .Z(n2402) );
  MUX2_X1 U1421 ( .A(n2402), .B(n2399), .S(n150), .Z(n2403) );
  MUX2_X1 U1422 ( .A(\REGISTERS[14][6] ), .B(\REGISTERS[30][6] ), .S(n189), 
        .Z(n2404) );
  MUX2_X1 U1423 ( .A(\REGISTERS[6][6] ), .B(\REGISTERS[22][6] ), .S(n189), .Z(
        n2405) );
  MUX2_X1 U1424 ( .A(n2405), .B(n2404), .S(n163), .Z(n2406) );
  MUX2_X1 U1425 ( .A(\REGISTERS[10][6] ), .B(\REGISTERS[26][6] ), .S(n189), 
        .Z(n2407) );
  MUX2_X1 U1426 ( .A(\REGISTERS[2][6] ), .B(\REGISTERS[18][6] ), .S(n189), .Z(
        n2408) );
  MUX2_X1 U1427 ( .A(n2408), .B(n2407), .S(n163), .Z(n2409) );
  MUX2_X1 U1428 ( .A(n2409), .B(n2406), .S(n150), .Z(n2410) );
  MUX2_X1 U1429 ( .A(n2410), .B(n2403), .S(ADD_RD1[0]), .Z(n2411) );
  MUX2_X1 U1430 ( .A(\REGISTERS[13][6] ), .B(\REGISTERS[29][6] ), .S(n189), 
        .Z(n2412) );
  MUX2_X1 U1431 ( .A(\REGISTERS[5][6] ), .B(\REGISTERS[21][6] ), .S(n189), .Z(
        n2413) );
  MUX2_X1 U1432 ( .A(n2413), .B(n2412), .S(n163), .Z(n2414) );
  MUX2_X1 U1433 ( .A(\REGISTERS[9][6] ), .B(\REGISTERS[25][6] ), .S(n189), .Z(
        n2415) );
  MUX2_X1 U1434 ( .A(\REGISTERS[1][6] ), .B(\REGISTERS[17][6] ), .S(n189), .Z(
        n2416) );
  MUX2_X1 U1435 ( .A(n2416), .B(n2415), .S(n163), .Z(n2417) );
  MUX2_X1 U1436 ( .A(n2417), .B(n2414), .S(n150), .Z(n2418) );
  MUX2_X1 U1437 ( .A(\REGISTERS[12][6] ), .B(\REGISTERS[28][6] ), .S(n190), 
        .Z(n2419) );
  MUX2_X1 U1438 ( .A(\REGISTERS[4][6] ), .B(\REGISTERS[20][6] ), .S(n190), .Z(
        n2420) );
  MUX2_X1 U1439 ( .A(n2420), .B(n2419), .S(n163), .Z(n2421) );
  MUX2_X1 U1440 ( .A(\REGISTERS[8][6] ), .B(\REGISTERS[24][6] ), .S(n190), .Z(
        n2422) );
  MUX2_X1 U1441 ( .A(\REGISTERS[0][6] ), .B(\REGISTERS[16][6] ), .S(n190), .Z(
        n2423) );
  MUX2_X1 U1442 ( .A(n2423), .B(n2422), .S(n163), .Z(n2424) );
  MUX2_X1 U1443 ( .A(n2424), .B(n2421), .S(n150), .Z(n2425) );
  MUX2_X1 U1444 ( .A(n2425), .B(n2418), .S(ADD_RD1[0]), .Z(n2426) );
  MUX2_X1 U1445 ( .A(n2426), .B(n2411), .S(ADD_RD1[1]), .Z(N385) );
  MUX2_X1 U1446 ( .A(\REGISTERS[15][7] ), .B(\REGISTERS[31][7] ), .S(n190), 
        .Z(n2427) );
  MUX2_X1 U1447 ( .A(\REGISTERS[7][7] ), .B(\REGISTERS[23][7] ), .S(n190), .Z(
        n2428) );
  MUX2_X1 U1448 ( .A(n2428), .B(n2427), .S(n163), .Z(n2429) );
  MUX2_X1 U1449 ( .A(\REGISTERS[11][7] ), .B(\REGISTERS[27][7] ), .S(n190), 
        .Z(n2430) );
  MUX2_X1 U1450 ( .A(\REGISTERS[3][7] ), .B(\REGISTERS[19][7] ), .S(n190), .Z(
        n2431) );
  MUX2_X1 U1451 ( .A(n2431), .B(n2430), .S(n163), .Z(n2432) );
  MUX2_X1 U1452 ( .A(n2432), .B(n2429), .S(n150), .Z(n2433) );
  MUX2_X1 U1453 ( .A(\REGISTERS[14][7] ), .B(\REGISTERS[30][7] ), .S(n190), 
        .Z(n2434) );
  MUX2_X1 U1454 ( .A(\REGISTERS[6][7] ), .B(\REGISTERS[22][7] ), .S(n190), .Z(
        n2435) );
  MUX2_X1 U1455 ( .A(n2435), .B(n2434), .S(n163), .Z(n2436) );
  MUX2_X1 U1456 ( .A(\REGISTERS[10][7] ), .B(\REGISTERS[26][7] ), .S(n190), 
        .Z(n2437) );
  MUX2_X1 U1457 ( .A(\REGISTERS[2][7] ), .B(\REGISTERS[18][7] ), .S(n190), .Z(
        n2438) );
  MUX2_X1 U1458 ( .A(n2438), .B(n2437), .S(n163), .Z(n2439) );
  MUX2_X1 U1459 ( .A(n2439), .B(n2436), .S(n150), .Z(n2440) );
  MUX2_X1 U1460 ( .A(n2440), .B(n2433), .S(ADD_RD1[0]), .Z(n2441) );
  MUX2_X1 U1461 ( .A(\REGISTERS[13][7] ), .B(\REGISTERS[29][7] ), .S(n191), 
        .Z(n2442) );
  MUX2_X1 U1462 ( .A(\REGISTERS[5][7] ), .B(\REGISTERS[21][7] ), .S(n191), .Z(
        n2443) );
  MUX2_X1 U1463 ( .A(n2443), .B(n2442), .S(n164), .Z(n2444) );
  MUX2_X1 U1464 ( .A(\REGISTERS[9][7] ), .B(\REGISTERS[25][7] ), .S(n191), .Z(
        n2445) );
  MUX2_X1 U1465 ( .A(\REGISTERS[1][7] ), .B(\REGISTERS[17][7] ), .S(n191), .Z(
        n2446) );
  MUX2_X1 U1466 ( .A(n2446), .B(n2445), .S(n164), .Z(n2447) );
  MUX2_X1 U1467 ( .A(n2447), .B(n2444), .S(n150), .Z(n2448) );
  MUX2_X1 U1468 ( .A(\REGISTERS[12][7] ), .B(\REGISTERS[28][7] ), .S(n191), 
        .Z(n2449) );
  MUX2_X1 U1469 ( .A(\REGISTERS[4][7] ), .B(\REGISTERS[20][7] ), .S(n191), .Z(
        n2450) );
  MUX2_X1 U1470 ( .A(n2450), .B(n2449), .S(n164), .Z(n2451) );
  MUX2_X1 U1471 ( .A(\REGISTERS[8][7] ), .B(\REGISTERS[24][7] ), .S(n191), .Z(
        n2452) );
  MUX2_X1 U1472 ( .A(\REGISTERS[0][7] ), .B(\REGISTERS[16][7] ), .S(n191), .Z(
        n2453) );
  MUX2_X1 U1473 ( .A(n2453), .B(n2452), .S(n164), .Z(n2454) );
  MUX2_X1 U1474 ( .A(n2454), .B(n2451), .S(n150), .Z(n2455) );
  MUX2_X1 U1475 ( .A(n2455), .B(n2448), .S(ADD_RD1[0]), .Z(n2456) );
  MUX2_X1 U1476 ( .A(n2456), .B(n2441), .S(ADD_RD1[1]), .Z(N386) );
  MUX2_X1 U1477 ( .A(\REGISTERS[15][8] ), .B(\REGISTERS[31][8] ), .S(n191), 
        .Z(n2457) );
  MUX2_X1 U1478 ( .A(\REGISTERS[7][8] ), .B(\REGISTERS[23][8] ), .S(n191), .Z(
        n2458) );
  MUX2_X1 U1479 ( .A(n2458), .B(n2457), .S(n164), .Z(n2459) );
  MUX2_X1 U1480 ( .A(\REGISTERS[11][8] ), .B(\REGISTERS[27][8] ), .S(n191), 
        .Z(n2460) );
  MUX2_X1 U1481 ( .A(\REGISTERS[3][8] ), .B(\REGISTERS[19][8] ), .S(n191), .Z(
        n2461) );
  MUX2_X1 U1482 ( .A(n2461), .B(n2460), .S(n164), .Z(n2462) );
  MUX2_X1 U1483 ( .A(n2462), .B(n2459), .S(n150), .Z(n2463) );
  MUX2_X1 U1484 ( .A(\REGISTERS[14][8] ), .B(\REGISTERS[30][8] ), .S(n192), 
        .Z(n2464) );
  MUX2_X1 U1485 ( .A(\REGISTERS[6][8] ), .B(\REGISTERS[22][8] ), .S(n192), .Z(
        n2465) );
  MUX2_X1 U1486 ( .A(n2465), .B(n2464), .S(n164), .Z(n2466) );
  MUX2_X1 U1487 ( .A(\REGISTERS[10][8] ), .B(\REGISTERS[26][8] ), .S(n192), 
        .Z(n2467) );
  MUX2_X1 U1488 ( .A(\REGISTERS[2][8] ), .B(\REGISTERS[18][8] ), .S(n192), .Z(
        n2468) );
  MUX2_X1 U1489 ( .A(n2468), .B(n2467), .S(n164), .Z(n2469) );
  MUX2_X1 U1490 ( .A(n2469), .B(n2466), .S(n150), .Z(n2470) );
  MUX2_X1 U1491 ( .A(n2470), .B(n2463), .S(ADD_RD1[0]), .Z(n2471) );
  MUX2_X1 U1492 ( .A(\REGISTERS[13][8] ), .B(\REGISTERS[29][8] ), .S(n192), 
        .Z(n2472) );
  MUX2_X1 U1493 ( .A(\REGISTERS[5][8] ), .B(\REGISTERS[21][8] ), .S(n192), .Z(
        n2473) );
  MUX2_X1 U1494 ( .A(n2473), .B(n2472), .S(n164), .Z(n2474) );
  MUX2_X1 U1495 ( .A(\REGISTERS[9][8] ), .B(\REGISTERS[25][8] ), .S(n192), .Z(
        n2475) );
  MUX2_X1 U1496 ( .A(\REGISTERS[1][8] ), .B(\REGISTERS[17][8] ), .S(n192), .Z(
        n2476) );
  MUX2_X1 U1497 ( .A(n2476), .B(n2475), .S(n164), .Z(n2477) );
  MUX2_X1 U1498 ( .A(n2477), .B(n2474), .S(n150), .Z(n2478) );
  MUX2_X1 U1499 ( .A(\REGISTERS[12][8] ), .B(\REGISTERS[28][8] ), .S(n192), 
        .Z(n2479) );
  MUX2_X1 U1500 ( .A(\REGISTERS[4][8] ), .B(\REGISTERS[20][8] ), .S(n192), .Z(
        n2480) );
  MUX2_X1 U1501 ( .A(n2480), .B(n2479), .S(n164), .Z(n2481) );
  MUX2_X1 U1502 ( .A(\REGISTERS[8][8] ), .B(\REGISTERS[24][8] ), .S(n192), .Z(
        n2482) );
  MUX2_X1 U1503 ( .A(\REGISTERS[0][8] ), .B(\REGISTERS[16][8] ), .S(n192), .Z(
        n2483) );
  MUX2_X1 U1504 ( .A(n2483), .B(n2482), .S(n164), .Z(n2484) );
  MUX2_X1 U1505 ( .A(n2484), .B(n2481), .S(n150), .Z(n2485) );
  MUX2_X1 U1506 ( .A(n2485), .B(n2478), .S(ADD_RD1[0]), .Z(n2486) );
  MUX2_X1 U1507 ( .A(n2486), .B(n2471), .S(ADD_RD1[1]), .Z(N387) );
  MUX2_X1 U1508 ( .A(\REGISTERS[15][9] ), .B(\REGISTERS[31][9] ), .S(n193), 
        .Z(n2487) );
  MUX2_X1 U1509 ( .A(\REGISTERS[7][9] ), .B(\REGISTERS[23][9] ), .S(n193), .Z(
        n2488) );
  MUX2_X1 U1510 ( .A(n2488), .B(n2487), .S(n165), .Z(n2489) );
  MUX2_X1 U1511 ( .A(\REGISTERS[11][9] ), .B(\REGISTERS[27][9] ), .S(n193), 
        .Z(n2490) );
  MUX2_X1 U1512 ( .A(\REGISTERS[3][9] ), .B(\REGISTERS[19][9] ), .S(n193), .Z(
        n2491) );
  MUX2_X1 U1513 ( .A(n2491), .B(n2490), .S(n165), .Z(n2492) );
  MUX2_X1 U1514 ( .A(n2492), .B(n2489), .S(n151), .Z(n2493) );
  MUX2_X1 U1515 ( .A(\REGISTERS[14][9] ), .B(\REGISTERS[30][9] ), .S(n193), 
        .Z(n2494) );
  MUX2_X1 U1516 ( .A(\REGISTERS[6][9] ), .B(\REGISTERS[22][9] ), .S(n193), .Z(
        n2495) );
  MUX2_X1 U1517 ( .A(n2495), .B(n2494), .S(n165), .Z(n2496) );
  MUX2_X1 U1518 ( .A(\REGISTERS[10][9] ), .B(\REGISTERS[26][9] ), .S(n193), 
        .Z(n2497) );
  MUX2_X1 U1519 ( .A(\REGISTERS[2][9] ), .B(\REGISTERS[18][9] ), .S(n193), .Z(
        n2498) );
  MUX2_X1 U1520 ( .A(n2498), .B(n2497), .S(n165), .Z(n2499) );
  MUX2_X1 U1521 ( .A(n2499), .B(n2496), .S(n151), .Z(n2500) );
  MUX2_X1 U1522 ( .A(n2500), .B(n2493), .S(ADD_RD1[0]), .Z(n2501) );
  MUX2_X1 U1523 ( .A(\REGISTERS[13][9] ), .B(\REGISTERS[29][9] ), .S(n193), 
        .Z(n2502) );
  MUX2_X1 U1524 ( .A(\REGISTERS[5][9] ), .B(\REGISTERS[21][9] ), .S(n193), .Z(
        n2503) );
  MUX2_X1 U1525 ( .A(n2503), .B(n2502), .S(n165), .Z(n2504) );
  MUX2_X1 U1526 ( .A(\REGISTERS[9][9] ), .B(\REGISTERS[25][9] ), .S(n193), .Z(
        n2505) );
  MUX2_X1 U1527 ( .A(\REGISTERS[1][9] ), .B(\REGISTERS[17][9] ), .S(n193), .Z(
        n2506) );
  MUX2_X1 U1528 ( .A(n2506), .B(n2505), .S(n165), .Z(n2507) );
  MUX2_X1 U1529 ( .A(n2507), .B(n2504), .S(n151), .Z(n2508) );
  MUX2_X1 U1530 ( .A(\REGISTERS[12][9] ), .B(\REGISTERS[28][9] ), .S(n194), 
        .Z(n2509) );
  MUX2_X1 U1531 ( .A(\REGISTERS[4][9] ), .B(\REGISTERS[20][9] ), .S(n194), .Z(
        n2510) );
  MUX2_X1 U1532 ( .A(n2510), .B(n2509), .S(n165), .Z(n2511) );
  MUX2_X1 U1533 ( .A(\REGISTERS[8][9] ), .B(\REGISTERS[24][9] ), .S(n194), .Z(
        n2512) );
  MUX2_X1 U1534 ( .A(\REGISTERS[0][9] ), .B(\REGISTERS[16][9] ), .S(n194), .Z(
        n2513) );
  MUX2_X1 U1535 ( .A(n2513), .B(n2512), .S(n165), .Z(n2514) );
  MUX2_X1 U1536 ( .A(n2514), .B(n2511), .S(n151), .Z(n2515) );
  MUX2_X1 U1537 ( .A(n2515), .B(n2508), .S(ADD_RD1[0]), .Z(n2516) );
  MUX2_X1 U1538 ( .A(n2516), .B(n2501), .S(ADD_RD1[1]), .Z(N388) );
  MUX2_X1 U1539 ( .A(\REGISTERS[15][10] ), .B(\REGISTERS[31][10] ), .S(n194), 
        .Z(n2517) );
  MUX2_X1 U1540 ( .A(\REGISTERS[7][10] ), .B(\REGISTERS[23][10] ), .S(n194), 
        .Z(n2518) );
  MUX2_X1 U1541 ( .A(n2518), .B(n2517), .S(n165), .Z(n2519) );
  MUX2_X1 U1542 ( .A(\REGISTERS[11][10] ), .B(\REGISTERS[27][10] ), .S(n194), 
        .Z(n2520) );
  MUX2_X1 U1543 ( .A(\REGISTERS[3][10] ), .B(\REGISTERS[19][10] ), .S(n194), 
        .Z(n2521) );
  MUX2_X1 U1544 ( .A(n2521), .B(n2520), .S(n165), .Z(n2522) );
  MUX2_X1 U1545 ( .A(n2522), .B(n2519), .S(n151), .Z(n2523) );
  MUX2_X1 U1546 ( .A(\REGISTERS[14][10] ), .B(\REGISTERS[30][10] ), .S(n194), 
        .Z(n2524) );
  MUX2_X1 U1547 ( .A(\REGISTERS[6][10] ), .B(\REGISTERS[22][10] ), .S(n194), 
        .Z(n2525) );
  MUX2_X1 U1548 ( .A(n2525), .B(n2524), .S(n165), .Z(n2526) );
  MUX2_X1 U1549 ( .A(\REGISTERS[10][10] ), .B(\REGISTERS[26][10] ), .S(n194), 
        .Z(n2527) );
  MUX2_X1 U1550 ( .A(\REGISTERS[2][10] ), .B(\REGISTERS[18][10] ), .S(n194), 
        .Z(n2528) );
  MUX2_X1 U1551 ( .A(n2528), .B(n2527), .S(n165), .Z(n2529) );
  MUX2_X1 U1552 ( .A(n2529), .B(n2526), .S(n151), .Z(n2530) );
  MUX2_X1 U1553 ( .A(n2530), .B(n2523), .S(ADD_RD1[0]), .Z(n2531) );
  MUX2_X1 U1554 ( .A(\REGISTERS[13][10] ), .B(\REGISTERS[29][10] ), .S(n195), 
        .Z(n2532) );
  MUX2_X1 U1555 ( .A(\REGISTERS[5][10] ), .B(\REGISTERS[21][10] ), .S(n195), 
        .Z(n2533) );
  MUX2_X1 U1556 ( .A(n2533), .B(n2532), .S(n166), .Z(n2534) );
  MUX2_X1 U1557 ( .A(\REGISTERS[9][10] ), .B(\REGISTERS[25][10] ), .S(n195), 
        .Z(n2535) );
  MUX2_X1 U1558 ( .A(\REGISTERS[1][10] ), .B(\REGISTERS[17][10] ), .S(n195), 
        .Z(n2536) );
  MUX2_X1 U1559 ( .A(n2536), .B(n2535), .S(n166), .Z(n2537) );
  MUX2_X1 U1560 ( .A(n2537), .B(n2534), .S(n151), .Z(n2538) );
  MUX2_X1 U1561 ( .A(\REGISTERS[12][10] ), .B(\REGISTERS[28][10] ), .S(n195), 
        .Z(n2539) );
  MUX2_X1 U1562 ( .A(\REGISTERS[4][10] ), .B(\REGISTERS[20][10] ), .S(n195), 
        .Z(n2540) );
  MUX2_X1 U1563 ( .A(n2540), .B(n2539), .S(n166), .Z(n2541) );
  MUX2_X1 U1564 ( .A(\REGISTERS[8][10] ), .B(\REGISTERS[24][10] ), .S(n195), 
        .Z(n2542) );
  MUX2_X1 U1565 ( .A(\REGISTERS[0][10] ), .B(\REGISTERS[16][10] ), .S(n195), 
        .Z(n2543) );
  MUX2_X1 U1566 ( .A(n2543), .B(n2542), .S(n166), .Z(n2544) );
  MUX2_X1 U1567 ( .A(n2544), .B(n2541), .S(n151), .Z(n2545) );
  MUX2_X1 U1568 ( .A(n2545), .B(n2538), .S(ADD_RD1[0]), .Z(n2546) );
  MUX2_X1 U1569 ( .A(n2546), .B(n2531), .S(ADD_RD1[1]), .Z(N389) );
  MUX2_X1 U1570 ( .A(\REGISTERS[15][11] ), .B(\REGISTERS[31][11] ), .S(n195), 
        .Z(n2547) );
  MUX2_X1 U1571 ( .A(\REGISTERS[7][11] ), .B(\REGISTERS[23][11] ), .S(n195), 
        .Z(n2548) );
  MUX2_X1 U1572 ( .A(n2548), .B(n2547), .S(n166), .Z(n2549) );
  MUX2_X1 U1573 ( .A(\REGISTERS[11][11] ), .B(\REGISTERS[27][11] ), .S(n195), 
        .Z(n2550) );
  MUX2_X1 U1574 ( .A(\REGISTERS[3][11] ), .B(\REGISTERS[19][11] ), .S(n195), 
        .Z(n2551) );
  MUX2_X1 U1575 ( .A(n2551), .B(n2550), .S(n166), .Z(n2552) );
  MUX2_X1 U1576 ( .A(n2552), .B(n2549), .S(n151), .Z(n2553) );
  MUX2_X1 U1577 ( .A(\REGISTERS[14][11] ), .B(\REGISTERS[30][11] ), .S(n196), 
        .Z(n2554) );
  MUX2_X1 U1578 ( .A(\REGISTERS[6][11] ), .B(\REGISTERS[22][11] ), .S(n196), 
        .Z(n2555) );
  MUX2_X1 U1579 ( .A(n2555), .B(n2554), .S(n166), .Z(n2556) );
  MUX2_X1 U1580 ( .A(\REGISTERS[10][11] ), .B(\REGISTERS[26][11] ), .S(n196), 
        .Z(n2557) );
  MUX2_X1 U1581 ( .A(\REGISTERS[2][11] ), .B(\REGISTERS[18][11] ), .S(n196), 
        .Z(n2558) );
  MUX2_X1 U1582 ( .A(n2558), .B(n2557), .S(n166), .Z(n2559) );
  MUX2_X1 U1583 ( .A(n2559), .B(n2556), .S(n151), .Z(n2560) );
  MUX2_X1 U1584 ( .A(n2560), .B(n2553), .S(ADD_RD1[0]), .Z(n2561) );
  MUX2_X1 U1585 ( .A(\REGISTERS[13][11] ), .B(\REGISTERS[29][11] ), .S(n196), 
        .Z(n2562) );
  MUX2_X1 U1586 ( .A(\REGISTERS[5][11] ), .B(\REGISTERS[21][11] ), .S(n196), 
        .Z(n2563) );
  MUX2_X1 U1587 ( .A(n2563), .B(n2562), .S(n166), .Z(n2564) );
  MUX2_X1 U1588 ( .A(\REGISTERS[9][11] ), .B(\REGISTERS[25][11] ), .S(n196), 
        .Z(n2565) );
  MUX2_X1 U1589 ( .A(\REGISTERS[1][11] ), .B(\REGISTERS[17][11] ), .S(n196), 
        .Z(n2566) );
  MUX2_X1 U1590 ( .A(n2566), .B(n2565), .S(n166), .Z(n2567) );
  MUX2_X1 U1591 ( .A(n2567), .B(n2564), .S(n151), .Z(n2568) );
  MUX2_X1 U1592 ( .A(\REGISTERS[12][11] ), .B(\REGISTERS[28][11] ), .S(n196), 
        .Z(n2569) );
  MUX2_X1 U1593 ( .A(\REGISTERS[4][11] ), .B(\REGISTERS[20][11] ), .S(n196), 
        .Z(n2570) );
  MUX2_X1 U1594 ( .A(n2570), .B(n2569), .S(n166), .Z(n2571) );
  MUX2_X1 U1595 ( .A(\REGISTERS[8][11] ), .B(\REGISTERS[24][11] ), .S(n196), 
        .Z(n2572) );
  MUX2_X1 U1596 ( .A(\REGISTERS[0][11] ), .B(\REGISTERS[16][11] ), .S(n196), 
        .Z(n2573) );
  MUX2_X1 U1597 ( .A(n2573), .B(n2572), .S(n166), .Z(n2574) );
  MUX2_X1 U1598 ( .A(n2574), .B(n2571), .S(n151), .Z(n2575) );
  MUX2_X1 U1599 ( .A(n2575), .B(n2568), .S(ADD_RD1[0]), .Z(n2576) );
  MUX2_X1 U1600 ( .A(n2576), .B(n2561), .S(ADD_RD1[1]), .Z(N390) );
  MUX2_X1 U1601 ( .A(\REGISTERS[15][12] ), .B(\REGISTERS[31][12] ), .S(n197), 
        .Z(n2577) );
  MUX2_X1 U1602 ( .A(\REGISTERS[7][12] ), .B(\REGISTERS[23][12] ), .S(n197), 
        .Z(n2578) );
  MUX2_X1 U1603 ( .A(n2578), .B(n2577), .S(n167), .Z(n2579) );
  MUX2_X1 U1604 ( .A(\REGISTERS[11][12] ), .B(\REGISTERS[27][12] ), .S(n197), 
        .Z(n2580) );
  MUX2_X1 U1605 ( .A(\REGISTERS[3][12] ), .B(\REGISTERS[19][12] ), .S(n197), 
        .Z(n2581) );
  MUX2_X1 U1606 ( .A(n2581), .B(n2580), .S(n167), .Z(n2582) );
  MUX2_X1 U1607 ( .A(n2582), .B(n2579), .S(n152), .Z(n2583) );
  MUX2_X1 U1608 ( .A(\REGISTERS[14][12] ), .B(\REGISTERS[30][12] ), .S(n197), 
        .Z(n2584) );
  MUX2_X1 U1609 ( .A(\REGISTERS[6][12] ), .B(\REGISTERS[22][12] ), .S(n197), 
        .Z(n2585) );
  MUX2_X1 U1610 ( .A(n2585), .B(n2584), .S(n167), .Z(n2586) );
  MUX2_X1 U1611 ( .A(\REGISTERS[10][12] ), .B(\REGISTERS[26][12] ), .S(n197), 
        .Z(n2587) );
  MUX2_X1 U1612 ( .A(\REGISTERS[2][12] ), .B(\REGISTERS[18][12] ), .S(n197), 
        .Z(n2588) );
  MUX2_X1 U1613 ( .A(n2588), .B(n2587), .S(n167), .Z(n2589) );
  MUX2_X1 U1614 ( .A(n2589), .B(n2586), .S(n152), .Z(n2590) );
  MUX2_X1 U1615 ( .A(n2590), .B(n2583), .S(ADD_RD1[0]), .Z(n2591) );
  MUX2_X1 U1616 ( .A(\REGISTERS[13][12] ), .B(\REGISTERS[29][12] ), .S(n197), 
        .Z(n2592) );
  MUX2_X1 U1617 ( .A(\REGISTERS[5][12] ), .B(\REGISTERS[21][12] ), .S(n197), 
        .Z(n2593) );
  MUX2_X1 U1618 ( .A(n2593), .B(n2592), .S(n167), .Z(n2594) );
  MUX2_X1 U1619 ( .A(\REGISTERS[9][12] ), .B(\REGISTERS[25][12] ), .S(n197), 
        .Z(n2595) );
  MUX2_X1 U1620 ( .A(\REGISTERS[1][12] ), .B(\REGISTERS[17][12] ), .S(n197), 
        .Z(n2596) );
  MUX2_X1 U1621 ( .A(n2596), .B(n2595), .S(n167), .Z(n2597) );
  MUX2_X1 U1622 ( .A(n2597), .B(n2594), .S(n152), .Z(n2598) );
  MUX2_X1 U1623 ( .A(\REGISTERS[12][12] ), .B(\REGISTERS[28][12] ), .S(n198), 
        .Z(n2599) );
  MUX2_X1 U1624 ( .A(\REGISTERS[4][12] ), .B(\REGISTERS[20][12] ), .S(n198), 
        .Z(n2600) );
  MUX2_X1 U1625 ( .A(n2600), .B(n2599), .S(n167), .Z(n2601) );
  MUX2_X1 U1626 ( .A(\REGISTERS[8][12] ), .B(\REGISTERS[24][12] ), .S(n198), 
        .Z(n2602) );
  MUX2_X1 U1627 ( .A(\REGISTERS[0][12] ), .B(\REGISTERS[16][12] ), .S(n198), 
        .Z(n2603) );
  MUX2_X1 U1628 ( .A(n2603), .B(n2602), .S(n167), .Z(n2604) );
  MUX2_X1 U1629 ( .A(n2604), .B(n2601), .S(n152), .Z(n2605) );
  MUX2_X1 U1630 ( .A(n2605), .B(n2598), .S(ADD_RD1[0]), .Z(n2606) );
  MUX2_X1 U1631 ( .A(n2606), .B(n2591), .S(ADD_RD1[1]), .Z(N391) );
  MUX2_X1 U1632 ( .A(\REGISTERS[15][13] ), .B(\REGISTERS[31][13] ), .S(n198), 
        .Z(n2607) );
  MUX2_X1 U1633 ( .A(\REGISTERS[7][13] ), .B(\REGISTERS[23][13] ), .S(n198), 
        .Z(n2608) );
  MUX2_X1 U1634 ( .A(n2608), .B(n2607), .S(n167), .Z(n2609) );
  MUX2_X1 U1635 ( .A(\REGISTERS[11][13] ), .B(\REGISTERS[27][13] ), .S(n198), 
        .Z(n2610) );
  MUX2_X1 U1636 ( .A(\REGISTERS[3][13] ), .B(\REGISTERS[19][13] ), .S(n198), 
        .Z(n2611) );
  MUX2_X1 U1637 ( .A(n2611), .B(n2610), .S(n167), .Z(n2612) );
  MUX2_X1 U1638 ( .A(n2612), .B(n2609), .S(n152), .Z(n2613) );
  MUX2_X1 U1639 ( .A(\REGISTERS[14][13] ), .B(\REGISTERS[30][13] ), .S(n198), 
        .Z(n2614) );
  MUX2_X1 U1640 ( .A(\REGISTERS[6][13] ), .B(\REGISTERS[22][13] ), .S(n198), 
        .Z(n2615) );
  MUX2_X1 U1641 ( .A(n2615), .B(n2614), .S(n167), .Z(n2616) );
  MUX2_X1 U1642 ( .A(\REGISTERS[10][13] ), .B(\REGISTERS[26][13] ), .S(n198), 
        .Z(n2617) );
  MUX2_X1 U1643 ( .A(\REGISTERS[2][13] ), .B(\REGISTERS[18][13] ), .S(n198), 
        .Z(n2618) );
  MUX2_X1 U1644 ( .A(n2618), .B(n2617), .S(n167), .Z(n2619) );
  MUX2_X1 U1645 ( .A(n2619), .B(n2616), .S(n152), .Z(n2620) );
  MUX2_X1 U1646 ( .A(n2620), .B(n2613), .S(ADD_RD1[0]), .Z(n2621) );
  MUX2_X1 U1647 ( .A(\REGISTERS[13][13] ), .B(\REGISTERS[29][13] ), .S(n199), 
        .Z(n2622) );
  MUX2_X1 U1648 ( .A(\REGISTERS[5][13] ), .B(\REGISTERS[21][13] ), .S(n199), 
        .Z(n2623) );
  MUX2_X1 U1649 ( .A(n2623), .B(n2622), .S(n168), .Z(n2624) );
  MUX2_X1 U1650 ( .A(\REGISTERS[9][13] ), .B(\REGISTERS[25][13] ), .S(n199), 
        .Z(n2625) );
  MUX2_X1 U1651 ( .A(\REGISTERS[1][13] ), .B(\REGISTERS[17][13] ), .S(n199), 
        .Z(n2626) );
  MUX2_X1 U1652 ( .A(n2626), .B(n2625), .S(n168), .Z(n2627) );
  MUX2_X1 U1653 ( .A(n2627), .B(n2624), .S(n152), .Z(n2628) );
  MUX2_X1 U1654 ( .A(\REGISTERS[12][13] ), .B(\REGISTERS[28][13] ), .S(n199), 
        .Z(n2629) );
  MUX2_X1 U1655 ( .A(\REGISTERS[4][13] ), .B(\REGISTERS[20][13] ), .S(n199), 
        .Z(n2630) );
  MUX2_X1 U1656 ( .A(n2630), .B(n2629), .S(n168), .Z(n2631) );
  MUX2_X1 U1657 ( .A(\REGISTERS[8][13] ), .B(\REGISTERS[24][13] ), .S(n199), 
        .Z(n2632) );
  MUX2_X1 U1658 ( .A(\REGISTERS[0][13] ), .B(\REGISTERS[16][13] ), .S(n199), 
        .Z(n2633) );
  MUX2_X1 U1659 ( .A(n2633), .B(n2632), .S(n168), .Z(n2634) );
  MUX2_X1 U1660 ( .A(n2634), .B(n2631), .S(n152), .Z(n2635) );
  MUX2_X1 U1661 ( .A(n2635), .B(n2628), .S(ADD_RD1[0]), .Z(n2636) );
  MUX2_X1 U1662 ( .A(n2636), .B(n2621), .S(ADD_RD1[1]), .Z(N392) );
  MUX2_X1 U1663 ( .A(\REGISTERS[15][14] ), .B(\REGISTERS[31][14] ), .S(n199), 
        .Z(n2637) );
  MUX2_X1 U1664 ( .A(\REGISTERS[7][14] ), .B(\REGISTERS[23][14] ), .S(n199), 
        .Z(n2638) );
  MUX2_X1 U1665 ( .A(n2638), .B(n2637), .S(n168), .Z(n2639) );
  MUX2_X1 U1666 ( .A(\REGISTERS[11][14] ), .B(\REGISTERS[27][14] ), .S(n199), 
        .Z(n2640) );
  MUX2_X1 U1667 ( .A(\REGISTERS[3][14] ), .B(\REGISTERS[19][14] ), .S(n199), 
        .Z(n2641) );
  MUX2_X1 U1668 ( .A(n2641), .B(n2640), .S(n168), .Z(n2642) );
  MUX2_X1 U1669 ( .A(n2642), .B(n2639), .S(n152), .Z(n2643) );
  MUX2_X1 U1670 ( .A(\REGISTERS[14][14] ), .B(\REGISTERS[30][14] ), .S(n200), 
        .Z(n2644) );
  MUX2_X1 U1671 ( .A(\REGISTERS[6][14] ), .B(\REGISTERS[22][14] ), .S(n200), 
        .Z(n2645) );
  MUX2_X1 U1672 ( .A(n2645), .B(n2644), .S(n168), .Z(n2646) );
  MUX2_X1 U1673 ( .A(\REGISTERS[10][14] ), .B(\REGISTERS[26][14] ), .S(n200), 
        .Z(n2647) );
  MUX2_X1 U1674 ( .A(\REGISTERS[2][14] ), .B(\REGISTERS[18][14] ), .S(n200), 
        .Z(n2648) );
  MUX2_X1 U1675 ( .A(n2648), .B(n2647), .S(n168), .Z(n2649) );
  MUX2_X1 U1676 ( .A(n2649), .B(n2646), .S(n152), .Z(n2650) );
  MUX2_X1 U1677 ( .A(n2650), .B(n2643), .S(ADD_RD1[0]), .Z(n2651) );
  MUX2_X1 U1678 ( .A(\REGISTERS[13][14] ), .B(\REGISTERS[29][14] ), .S(n200), 
        .Z(n2652) );
  MUX2_X1 U1679 ( .A(\REGISTERS[5][14] ), .B(\REGISTERS[21][14] ), .S(n200), 
        .Z(n2653) );
  MUX2_X1 U1680 ( .A(n2653), .B(n2652), .S(n168), .Z(n2654) );
  MUX2_X1 U1681 ( .A(\REGISTERS[9][14] ), .B(\REGISTERS[25][14] ), .S(n200), 
        .Z(n2655) );
  MUX2_X1 U1682 ( .A(\REGISTERS[1][14] ), .B(\REGISTERS[17][14] ), .S(n200), 
        .Z(n2656) );
  MUX2_X1 U1683 ( .A(n2656), .B(n2655), .S(n168), .Z(n2657) );
  MUX2_X1 U1684 ( .A(n2657), .B(n2654), .S(n152), .Z(n2658) );
  MUX2_X1 U1685 ( .A(\REGISTERS[12][14] ), .B(\REGISTERS[28][14] ), .S(n200), 
        .Z(n2659) );
  MUX2_X1 U1686 ( .A(\REGISTERS[4][14] ), .B(\REGISTERS[20][14] ), .S(n200), 
        .Z(n2660) );
  MUX2_X1 U1687 ( .A(n2660), .B(n2659), .S(n168), .Z(n2661) );
  MUX2_X1 U1688 ( .A(\REGISTERS[8][14] ), .B(\REGISTERS[24][14] ), .S(n200), 
        .Z(n2662) );
  MUX2_X1 U1689 ( .A(\REGISTERS[0][14] ), .B(\REGISTERS[16][14] ), .S(n200), 
        .Z(n2663) );
  MUX2_X1 U1690 ( .A(n2663), .B(n2662), .S(n168), .Z(n2664) );
  MUX2_X1 U1691 ( .A(n2664), .B(n2661), .S(n152), .Z(n2665) );
  MUX2_X1 U1692 ( .A(n2665), .B(n2658), .S(ADD_RD1[0]), .Z(n2666) );
  MUX2_X1 U1693 ( .A(n2666), .B(n2651), .S(ADD_RD1[1]), .Z(N393) );
  MUX2_X1 U1694 ( .A(\REGISTERS[15][15] ), .B(\REGISTERS[31][15] ), .S(n201), 
        .Z(n2667) );
  MUX2_X1 U1695 ( .A(\REGISTERS[7][15] ), .B(\REGISTERS[23][15] ), .S(n201), 
        .Z(n2668) );
  MUX2_X1 U1696 ( .A(n2668), .B(n2667), .S(n169), .Z(n2669) );
  MUX2_X1 U1697 ( .A(\REGISTERS[11][15] ), .B(\REGISTERS[27][15] ), .S(n201), 
        .Z(n2670) );
  MUX2_X1 U1698 ( .A(\REGISTERS[3][15] ), .B(\REGISTERS[19][15] ), .S(n201), 
        .Z(n2671) );
  MUX2_X1 U1699 ( .A(n2671), .B(n2670), .S(n169), .Z(n2672) );
  MUX2_X1 U1700 ( .A(n2672), .B(n2669), .S(n153), .Z(n2673) );
  MUX2_X1 U1701 ( .A(\REGISTERS[14][15] ), .B(\REGISTERS[30][15] ), .S(n201), 
        .Z(n2674) );
  MUX2_X1 U1702 ( .A(\REGISTERS[6][15] ), .B(\REGISTERS[22][15] ), .S(n201), 
        .Z(n2675) );
  MUX2_X1 U1703 ( .A(n2675), .B(n2674), .S(n169), .Z(n2676) );
  MUX2_X1 U1704 ( .A(\REGISTERS[10][15] ), .B(\REGISTERS[26][15] ), .S(n201), 
        .Z(n2677) );
  MUX2_X1 U1705 ( .A(\REGISTERS[2][15] ), .B(\REGISTERS[18][15] ), .S(n201), 
        .Z(n2678) );
  MUX2_X1 U1706 ( .A(n2678), .B(n2677), .S(n169), .Z(n2679) );
  MUX2_X1 U1707 ( .A(n2679), .B(n2676), .S(n153), .Z(n2680) );
  MUX2_X1 U1708 ( .A(n2680), .B(n2673), .S(ADD_RD1[0]), .Z(n2681) );
  MUX2_X1 U1709 ( .A(\REGISTERS[13][15] ), .B(\REGISTERS[29][15] ), .S(n201), 
        .Z(n2682) );
  MUX2_X1 U1710 ( .A(\REGISTERS[5][15] ), .B(\REGISTERS[21][15] ), .S(n201), 
        .Z(n2683) );
  MUX2_X1 U1711 ( .A(n2683), .B(n2682), .S(n169), .Z(n2684) );
  MUX2_X1 U1712 ( .A(\REGISTERS[9][15] ), .B(\REGISTERS[25][15] ), .S(n201), 
        .Z(n2685) );
  MUX2_X1 U1713 ( .A(\REGISTERS[1][15] ), .B(\REGISTERS[17][15] ), .S(n201), 
        .Z(n2686) );
  MUX2_X1 U1714 ( .A(n2686), .B(n2685), .S(n169), .Z(n2687) );
  MUX2_X1 U1715 ( .A(n2687), .B(n2684), .S(n153), .Z(n2688) );
  MUX2_X1 U1716 ( .A(\REGISTERS[12][15] ), .B(\REGISTERS[28][15] ), .S(n202), 
        .Z(n2689) );
  MUX2_X1 U1717 ( .A(\REGISTERS[4][15] ), .B(\REGISTERS[20][15] ), .S(n202), 
        .Z(n2690) );
  MUX2_X1 U1718 ( .A(n2690), .B(n2689), .S(n169), .Z(n2691) );
  MUX2_X1 U1719 ( .A(\REGISTERS[8][15] ), .B(\REGISTERS[24][15] ), .S(n202), 
        .Z(n2692) );
  MUX2_X1 U1720 ( .A(\REGISTERS[0][15] ), .B(\REGISTERS[16][15] ), .S(n202), 
        .Z(n2693) );
  MUX2_X1 U1721 ( .A(n2693), .B(n2692), .S(n169), .Z(n2694) );
  MUX2_X1 U1722 ( .A(n2694), .B(n2691), .S(n153), .Z(n2695) );
  MUX2_X1 U1723 ( .A(n2695), .B(n2688), .S(ADD_RD1[0]), .Z(n2696) );
  MUX2_X1 U1724 ( .A(n2696), .B(n2681), .S(ADD_RD1[1]), .Z(N394) );
  MUX2_X1 U1725 ( .A(\REGISTERS[15][16] ), .B(\REGISTERS[31][16] ), .S(n202), 
        .Z(n2697) );
  MUX2_X1 U1726 ( .A(\REGISTERS[7][16] ), .B(\REGISTERS[23][16] ), .S(n202), 
        .Z(n2698) );
  MUX2_X1 U1727 ( .A(n2698), .B(n2697), .S(n169), .Z(n2699) );
  MUX2_X1 U1728 ( .A(\REGISTERS[11][16] ), .B(\REGISTERS[27][16] ), .S(n202), 
        .Z(n2700) );
  MUX2_X1 U1729 ( .A(\REGISTERS[3][16] ), .B(\REGISTERS[19][16] ), .S(n202), 
        .Z(n2701) );
  MUX2_X1 U1730 ( .A(n2701), .B(n2700), .S(n169), .Z(n2702) );
  MUX2_X1 U1731 ( .A(n2702), .B(n2699), .S(n153), .Z(n2703) );
  MUX2_X1 U1732 ( .A(\REGISTERS[14][16] ), .B(\REGISTERS[30][16] ), .S(n202), 
        .Z(n2704) );
  MUX2_X1 U1733 ( .A(\REGISTERS[6][16] ), .B(\REGISTERS[22][16] ), .S(n202), 
        .Z(n2705) );
  MUX2_X1 U1734 ( .A(n2705), .B(n2704), .S(n169), .Z(n2706) );
  MUX2_X1 U1735 ( .A(\REGISTERS[10][16] ), .B(\REGISTERS[26][16] ), .S(n202), 
        .Z(n2707) );
  MUX2_X1 U1736 ( .A(\REGISTERS[2][16] ), .B(\REGISTERS[18][16] ), .S(n202), 
        .Z(n2708) );
  MUX2_X1 U1737 ( .A(n2708), .B(n2707), .S(n169), .Z(n2709) );
  MUX2_X1 U1738 ( .A(n2709), .B(n2706), .S(n153), .Z(n2710) );
  MUX2_X1 U1739 ( .A(n2710), .B(n2703), .S(ADD_RD1[0]), .Z(n2711) );
  MUX2_X1 U1740 ( .A(\REGISTERS[13][16] ), .B(\REGISTERS[29][16] ), .S(n203), 
        .Z(n2712) );
  MUX2_X1 U1741 ( .A(\REGISTERS[5][16] ), .B(\REGISTERS[21][16] ), .S(n203), 
        .Z(n2713) );
  MUX2_X1 U1742 ( .A(n2713), .B(n2712), .S(n170), .Z(n2714) );
  MUX2_X1 U1743 ( .A(\REGISTERS[9][16] ), .B(\REGISTERS[25][16] ), .S(n203), 
        .Z(n2715) );
  MUX2_X1 U1744 ( .A(\REGISTERS[1][16] ), .B(\REGISTERS[17][16] ), .S(n203), 
        .Z(n2716) );
  MUX2_X1 U1745 ( .A(n2716), .B(n2715), .S(n170), .Z(n2717) );
  MUX2_X1 U1746 ( .A(n2717), .B(n2714), .S(n153), .Z(n2718) );
  MUX2_X1 U1747 ( .A(\REGISTERS[12][16] ), .B(\REGISTERS[28][16] ), .S(n203), 
        .Z(n2719) );
  MUX2_X1 U1748 ( .A(\REGISTERS[4][16] ), .B(\REGISTERS[20][16] ), .S(n203), 
        .Z(n2720) );
  MUX2_X1 U1749 ( .A(n2720), .B(n2719), .S(n170), .Z(n2721) );
  MUX2_X1 U1750 ( .A(\REGISTERS[8][16] ), .B(\REGISTERS[24][16] ), .S(n203), 
        .Z(n2722) );
  MUX2_X1 U1751 ( .A(\REGISTERS[0][16] ), .B(\REGISTERS[16][16] ), .S(n203), 
        .Z(n2723) );
  MUX2_X1 U1752 ( .A(n2723), .B(n2722), .S(n170), .Z(n2724) );
  MUX2_X1 U1753 ( .A(n2724), .B(n2721), .S(n153), .Z(n2725) );
  MUX2_X1 U1754 ( .A(n2725), .B(n2718), .S(ADD_RD1[0]), .Z(n2726) );
  MUX2_X1 U1755 ( .A(n2726), .B(n2711), .S(ADD_RD1[1]), .Z(N395) );
  MUX2_X1 U1756 ( .A(\REGISTERS[15][17] ), .B(\REGISTERS[31][17] ), .S(n203), 
        .Z(n2727) );
  MUX2_X1 U1757 ( .A(\REGISTERS[7][17] ), .B(\REGISTERS[23][17] ), .S(n203), 
        .Z(n2728) );
  MUX2_X1 U1758 ( .A(n2728), .B(n2727), .S(n170), .Z(n2729) );
  MUX2_X1 U1759 ( .A(\REGISTERS[11][17] ), .B(\REGISTERS[27][17] ), .S(n203), 
        .Z(n2730) );
  MUX2_X1 U1760 ( .A(\REGISTERS[3][17] ), .B(\REGISTERS[19][17] ), .S(n203), 
        .Z(n2731) );
  MUX2_X1 U1761 ( .A(n2731), .B(n2730), .S(n170), .Z(n2732) );
  MUX2_X1 U1762 ( .A(n2732), .B(n2729), .S(n153), .Z(n2733) );
  MUX2_X1 U1763 ( .A(\REGISTERS[14][17] ), .B(\REGISTERS[30][17] ), .S(n204), 
        .Z(n2734) );
  MUX2_X1 U1764 ( .A(\REGISTERS[6][17] ), .B(\REGISTERS[22][17] ), .S(n204), 
        .Z(n2735) );
  MUX2_X1 U1765 ( .A(n2735), .B(n2734), .S(n170), .Z(n2736) );
  MUX2_X1 U1766 ( .A(\REGISTERS[10][17] ), .B(\REGISTERS[26][17] ), .S(n204), 
        .Z(n2737) );
  MUX2_X1 U1767 ( .A(\REGISTERS[2][17] ), .B(\REGISTERS[18][17] ), .S(n204), 
        .Z(n2738) );
  MUX2_X1 U1768 ( .A(n2738), .B(n2737), .S(n170), .Z(n2739) );
  MUX2_X1 U1769 ( .A(n2739), .B(n2736), .S(n153), .Z(n2740) );
  MUX2_X1 U1770 ( .A(n2740), .B(n2733), .S(ADD_RD1[0]), .Z(n2741) );
  MUX2_X1 U1771 ( .A(\REGISTERS[13][17] ), .B(\REGISTERS[29][17] ), .S(n204), 
        .Z(n2742) );
  MUX2_X1 U1772 ( .A(\REGISTERS[5][17] ), .B(\REGISTERS[21][17] ), .S(n204), 
        .Z(n2743) );
  MUX2_X1 U1773 ( .A(n2743), .B(n2742), .S(n170), .Z(n2744) );
  MUX2_X1 U1774 ( .A(\REGISTERS[9][17] ), .B(\REGISTERS[25][17] ), .S(n204), 
        .Z(n2745) );
  MUX2_X1 U1775 ( .A(\REGISTERS[1][17] ), .B(\REGISTERS[17][17] ), .S(n204), 
        .Z(n2746) );
  MUX2_X1 U1776 ( .A(n2746), .B(n2745), .S(n170), .Z(n2747) );
  MUX2_X1 U1777 ( .A(n2747), .B(n2744), .S(n153), .Z(n2748) );
  MUX2_X1 U1778 ( .A(\REGISTERS[12][17] ), .B(\REGISTERS[28][17] ), .S(n204), 
        .Z(n2749) );
  MUX2_X1 U1779 ( .A(\REGISTERS[4][17] ), .B(\REGISTERS[20][17] ), .S(n204), 
        .Z(n2750) );
  MUX2_X1 U1780 ( .A(n2750), .B(n2749), .S(n170), .Z(n2751) );
  MUX2_X1 U1781 ( .A(\REGISTERS[8][17] ), .B(\REGISTERS[24][17] ), .S(n204), 
        .Z(n2752) );
  MUX2_X1 U1782 ( .A(\REGISTERS[0][17] ), .B(\REGISTERS[16][17] ), .S(n204), 
        .Z(n2753) );
  MUX2_X1 U1783 ( .A(n2753), .B(n2752), .S(n170), .Z(n2754) );
  MUX2_X1 U1784 ( .A(n2754), .B(n2751), .S(n153), .Z(n2755) );
  MUX2_X1 U1785 ( .A(n2755), .B(n2748), .S(ADD_RD1[0]), .Z(n2756) );
  MUX2_X1 U1786 ( .A(n2756), .B(n2741), .S(ADD_RD1[1]), .Z(N396) );
  MUX2_X1 U1787 ( .A(\REGISTERS[15][18] ), .B(\REGISTERS[31][18] ), .S(n205), 
        .Z(n2757) );
  MUX2_X1 U1788 ( .A(\REGISTERS[7][18] ), .B(\REGISTERS[23][18] ), .S(n205), 
        .Z(n2758) );
  MUX2_X1 U1789 ( .A(n2758), .B(n2757), .S(n171), .Z(n2759) );
  MUX2_X1 U1790 ( .A(\REGISTERS[11][18] ), .B(\REGISTERS[27][18] ), .S(n205), 
        .Z(n2760) );
  MUX2_X1 U1791 ( .A(\REGISTERS[3][18] ), .B(\REGISTERS[19][18] ), .S(n205), 
        .Z(n2761) );
  MUX2_X1 U1792 ( .A(n2761), .B(n2760), .S(n171), .Z(n2762) );
  MUX2_X1 U1793 ( .A(n2762), .B(n2759), .S(n154), .Z(n2763) );
  MUX2_X1 U1794 ( .A(\REGISTERS[14][18] ), .B(\REGISTERS[30][18] ), .S(n205), 
        .Z(n2764) );
  MUX2_X1 U1795 ( .A(\REGISTERS[6][18] ), .B(\REGISTERS[22][18] ), .S(n205), 
        .Z(n2765) );
  MUX2_X1 U1796 ( .A(n2765), .B(n2764), .S(n171), .Z(n2766) );
  MUX2_X1 U1797 ( .A(\REGISTERS[10][18] ), .B(\REGISTERS[26][18] ), .S(n205), 
        .Z(n2767) );
  MUX2_X1 U1798 ( .A(\REGISTERS[2][18] ), .B(\REGISTERS[18][18] ), .S(n205), 
        .Z(n2768) );
  MUX2_X1 U1799 ( .A(n2768), .B(n2767), .S(n171), .Z(n2769) );
  MUX2_X1 U1800 ( .A(n2769), .B(n2766), .S(n154), .Z(n2770) );
  MUX2_X1 U1801 ( .A(n2770), .B(n2763), .S(ADD_RD1[0]), .Z(n2771) );
  MUX2_X1 U1802 ( .A(\REGISTERS[13][18] ), .B(\REGISTERS[29][18] ), .S(n205), 
        .Z(n2772) );
  MUX2_X1 U1803 ( .A(\REGISTERS[5][18] ), .B(\REGISTERS[21][18] ), .S(n205), 
        .Z(n2773) );
  MUX2_X1 U1804 ( .A(n2773), .B(n2772), .S(n171), .Z(n2774) );
  MUX2_X1 U1805 ( .A(\REGISTERS[9][18] ), .B(\REGISTERS[25][18] ), .S(n205), 
        .Z(n2775) );
  MUX2_X1 U1806 ( .A(\REGISTERS[1][18] ), .B(\REGISTERS[17][18] ), .S(n205), 
        .Z(n2776) );
  MUX2_X1 U1807 ( .A(n2776), .B(n2775), .S(n171), .Z(n2777) );
  MUX2_X1 U1808 ( .A(n2777), .B(n2774), .S(n154), .Z(n2778) );
  MUX2_X1 U1809 ( .A(\REGISTERS[12][18] ), .B(\REGISTERS[28][18] ), .S(n206), 
        .Z(n2779) );
  MUX2_X1 U1810 ( .A(\REGISTERS[4][18] ), .B(\REGISTERS[20][18] ), .S(n206), 
        .Z(n2780) );
  MUX2_X1 U1811 ( .A(n2780), .B(n2779), .S(n171), .Z(n2781) );
  MUX2_X1 U1812 ( .A(\REGISTERS[8][18] ), .B(\REGISTERS[24][18] ), .S(n206), 
        .Z(n2782) );
  MUX2_X1 U1813 ( .A(\REGISTERS[0][18] ), .B(\REGISTERS[16][18] ), .S(n206), 
        .Z(n2783) );
  MUX2_X1 U1814 ( .A(n2783), .B(n2782), .S(n171), .Z(n2784) );
  MUX2_X1 U1815 ( .A(n2784), .B(n2781), .S(n154), .Z(n2785) );
  MUX2_X1 U1816 ( .A(n2785), .B(n2778), .S(ADD_RD1[0]), .Z(n2786) );
  MUX2_X1 U1817 ( .A(n2786), .B(n2771), .S(ADD_RD1[1]), .Z(N397) );
  MUX2_X1 U1818 ( .A(\REGISTERS[15][19] ), .B(\REGISTERS[31][19] ), .S(n206), 
        .Z(n2787) );
  MUX2_X1 U1819 ( .A(\REGISTERS[7][19] ), .B(\REGISTERS[23][19] ), .S(n206), 
        .Z(n2788) );
  MUX2_X1 U1820 ( .A(n2788), .B(n2787), .S(n171), .Z(n2789) );
  MUX2_X1 U1821 ( .A(\REGISTERS[11][19] ), .B(\REGISTERS[27][19] ), .S(n206), 
        .Z(n2790) );
  MUX2_X1 U1822 ( .A(\REGISTERS[3][19] ), .B(\REGISTERS[19][19] ), .S(n206), 
        .Z(n2791) );
  MUX2_X1 U1823 ( .A(n2791), .B(n2790), .S(n171), .Z(n2792) );
  MUX2_X1 U1824 ( .A(n2792), .B(n2789), .S(n154), .Z(n2793) );
  MUX2_X1 U1825 ( .A(\REGISTERS[14][19] ), .B(\REGISTERS[30][19] ), .S(n206), 
        .Z(n2794) );
  MUX2_X1 U1826 ( .A(\REGISTERS[6][19] ), .B(\REGISTERS[22][19] ), .S(n206), 
        .Z(n2795) );
  MUX2_X1 U1827 ( .A(n2795), .B(n2794), .S(n171), .Z(n2796) );
  MUX2_X1 U1828 ( .A(\REGISTERS[10][19] ), .B(\REGISTERS[26][19] ), .S(n206), 
        .Z(n2797) );
  MUX2_X1 U1829 ( .A(\REGISTERS[2][19] ), .B(\REGISTERS[18][19] ), .S(n206), 
        .Z(n2798) );
  MUX2_X1 U1830 ( .A(n2798), .B(n2797), .S(n171), .Z(n2799) );
  MUX2_X1 U1831 ( .A(n2799), .B(n2796), .S(n154), .Z(n2800) );
  MUX2_X1 U1832 ( .A(n2800), .B(n2793), .S(ADD_RD1[0]), .Z(n2801) );
  MUX2_X1 U1833 ( .A(\REGISTERS[13][19] ), .B(\REGISTERS[29][19] ), .S(n207), 
        .Z(n2802) );
  MUX2_X1 U1834 ( .A(\REGISTERS[5][19] ), .B(\REGISTERS[21][19] ), .S(n207), 
        .Z(n2803) );
  MUX2_X1 U1835 ( .A(n2803), .B(n2802), .S(n172), .Z(n2804) );
  MUX2_X1 U1836 ( .A(\REGISTERS[9][19] ), .B(\REGISTERS[25][19] ), .S(n207), 
        .Z(n2805) );
  MUX2_X1 U1837 ( .A(\REGISTERS[1][19] ), .B(\REGISTERS[17][19] ), .S(n207), 
        .Z(n2806) );
  MUX2_X1 U1838 ( .A(n2806), .B(n2805), .S(n172), .Z(n2807) );
  MUX2_X1 U1839 ( .A(n2807), .B(n2804), .S(n154), .Z(n2808) );
  MUX2_X1 U1840 ( .A(\REGISTERS[12][19] ), .B(\REGISTERS[28][19] ), .S(n207), 
        .Z(n2809) );
  MUX2_X1 U1841 ( .A(\REGISTERS[4][19] ), .B(\REGISTERS[20][19] ), .S(n207), 
        .Z(n2810) );
  MUX2_X1 U1842 ( .A(n2810), .B(n2809), .S(n172), .Z(n2811) );
  MUX2_X1 U1843 ( .A(\REGISTERS[8][19] ), .B(\REGISTERS[24][19] ), .S(n207), 
        .Z(n2812) );
  MUX2_X1 U1844 ( .A(\REGISTERS[0][19] ), .B(\REGISTERS[16][19] ), .S(n207), 
        .Z(n2813) );
  MUX2_X1 U1845 ( .A(n2813), .B(n2812), .S(n172), .Z(n2814) );
  MUX2_X1 U1846 ( .A(n2814), .B(n2811), .S(n154), .Z(n2815) );
  MUX2_X1 U1847 ( .A(n2815), .B(n2808), .S(ADD_RD1[0]), .Z(n2816) );
  MUX2_X1 U1848 ( .A(n2816), .B(n2801), .S(ADD_RD1[1]), .Z(N398) );
  MUX2_X1 U1849 ( .A(\REGISTERS[15][20] ), .B(\REGISTERS[31][20] ), .S(n207), 
        .Z(n2817) );
  MUX2_X1 U1850 ( .A(\REGISTERS[7][20] ), .B(\REGISTERS[23][20] ), .S(n207), 
        .Z(n2818) );
  MUX2_X1 U1851 ( .A(n2818), .B(n2817), .S(n172), .Z(n2819) );
  MUX2_X1 U1852 ( .A(\REGISTERS[11][20] ), .B(\REGISTERS[27][20] ), .S(n207), 
        .Z(n2820) );
  MUX2_X1 U1853 ( .A(\REGISTERS[3][20] ), .B(\REGISTERS[19][20] ), .S(n207), 
        .Z(n2821) );
  MUX2_X1 U1854 ( .A(n2821), .B(n2820), .S(n172), .Z(n2822) );
  MUX2_X1 U1855 ( .A(n2822), .B(n2819), .S(n154), .Z(n2823) );
  MUX2_X1 U1856 ( .A(\REGISTERS[14][20] ), .B(\REGISTERS[30][20] ), .S(n208), 
        .Z(n2824) );
  MUX2_X1 U1857 ( .A(\REGISTERS[6][20] ), .B(\REGISTERS[22][20] ), .S(n208), 
        .Z(n2825) );
  MUX2_X1 U1858 ( .A(n2825), .B(n2824), .S(n172), .Z(n2826) );
  MUX2_X1 U1859 ( .A(\REGISTERS[10][20] ), .B(\REGISTERS[26][20] ), .S(n208), 
        .Z(n2827) );
  MUX2_X1 U1860 ( .A(\REGISTERS[2][20] ), .B(\REGISTERS[18][20] ), .S(n208), 
        .Z(n2828) );
  MUX2_X1 U1861 ( .A(n2828), .B(n2827), .S(n172), .Z(n2829) );
  MUX2_X1 U1862 ( .A(n2829), .B(n2826), .S(n154), .Z(n2830) );
  MUX2_X1 U1863 ( .A(n2830), .B(n2823), .S(ADD_RD1[0]), .Z(n2831) );
  MUX2_X1 U1864 ( .A(\REGISTERS[13][20] ), .B(\REGISTERS[29][20] ), .S(n208), 
        .Z(n2832) );
  MUX2_X1 U1865 ( .A(\REGISTERS[5][20] ), .B(\REGISTERS[21][20] ), .S(n208), 
        .Z(n2833) );
  MUX2_X1 U1866 ( .A(n2833), .B(n2832), .S(n172), .Z(n2834) );
  MUX2_X1 U1867 ( .A(\REGISTERS[9][20] ), .B(\REGISTERS[25][20] ), .S(n208), 
        .Z(n2835) );
  MUX2_X1 U1868 ( .A(\REGISTERS[1][20] ), .B(\REGISTERS[17][20] ), .S(n208), 
        .Z(n2836) );
  MUX2_X1 U1869 ( .A(n2836), .B(n2835), .S(n172), .Z(n2837) );
  MUX2_X1 U1870 ( .A(n2837), .B(n2834), .S(n154), .Z(n2838) );
  MUX2_X1 U1871 ( .A(\REGISTERS[12][20] ), .B(\REGISTERS[28][20] ), .S(n208), 
        .Z(n2839) );
  MUX2_X1 U1872 ( .A(\REGISTERS[4][20] ), .B(\REGISTERS[20][20] ), .S(n208), 
        .Z(n2840) );
  MUX2_X1 U1873 ( .A(n2840), .B(n2839), .S(n172), .Z(n2841) );
  MUX2_X1 U1874 ( .A(\REGISTERS[8][20] ), .B(\REGISTERS[24][20] ), .S(n208), 
        .Z(n2842) );
  MUX2_X1 U1875 ( .A(\REGISTERS[0][20] ), .B(\REGISTERS[16][20] ), .S(n208), 
        .Z(n2843) );
  MUX2_X1 U1876 ( .A(n2843), .B(n2842), .S(n172), .Z(n2844) );
  MUX2_X1 U1877 ( .A(n2844), .B(n2841), .S(n154), .Z(n2845) );
  MUX2_X1 U1878 ( .A(n2845), .B(n2838), .S(ADD_RD1[0]), .Z(n2846) );
  MUX2_X1 U1879 ( .A(n2846), .B(n2831), .S(ADD_RD1[1]), .Z(N399) );
  MUX2_X1 U1880 ( .A(\REGISTERS[15][21] ), .B(\REGISTERS[31][21] ), .S(n209), 
        .Z(n2847) );
  MUX2_X1 U1881 ( .A(\REGISTERS[7][21] ), .B(\REGISTERS[23][21] ), .S(n209), 
        .Z(n2848) );
  MUX2_X1 U1882 ( .A(n2848), .B(n2847), .S(n173), .Z(n2849) );
  MUX2_X1 U1883 ( .A(\REGISTERS[11][21] ), .B(\REGISTERS[27][21] ), .S(n209), 
        .Z(n2850) );
  MUX2_X1 U1884 ( .A(\REGISTERS[3][21] ), .B(\REGISTERS[19][21] ), .S(n209), 
        .Z(n2851) );
  MUX2_X1 U1885 ( .A(n2851), .B(n2850), .S(n173), .Z(n2852) );
  MUX2_X1 U1886 ( .A(n2852), .B(n2849), .S(n155), .Z(n2853) );
  MUX2_X1 U1887 ( .A(\REGISTERS[14][21] ), .B(\REGISTERS[30][21] ), .S(n209), 
        .Z(n2854) );
  MUX2_X1 U1888 ( .A(\REGISTERS[6][21] ), .B(\REGISTERS[22][21] ), .S(n209), 
        .Z(n2855) );
  MUX2_X1 U1889 ( .A(n2855), .B(n2854), .S(n173), .Z(n2856) );
  MUX2_X1 U1890 ( .A(\REGISTERS[10][21] ), .B(\REGISTERS[26][21] ), .S(n209), 
        .Z(n2857) );
  MUX2_X1 U1891 ( .A(\REGISTERS[2][21] ), .B(\REGISTERS[18][21] ), .S(n209), 
        .Z(n2858) );
  MUX2_X1 U1892 ( .A(n2858), .B(n2857), .S(n173), .Z(n2859) );
  MUX2_X1 U1893 ( .A(n2859), .B(n2856), .S(n155), .Z(n2860) );
  MUX2_X1 U1894 ( .A(n2860), .B(n2853), .S(ADD_RD1[0]), .Z(n2861) );
  MUX2_X1 U1895 ( .A(\REGISTERS[13][21] ), .B(\REGISTERS[29][21] ), .S(n209), 
        .Z(n2862) );
  MUX2_X1 U1896 ( .A(\REGISTERS[5][21] ), .B(\REGISTERS[21][21] ), .S(n209), 
        .Z(n2863) );
  MUX2_X1 U1897 ( .A(n2863), .B(n2862), .S(n173), .Z(n2864) );
  MUX2_X1 U1898 ( .A(\REGISTERS[9][21] ), .B(\REGISTERS[25][21] ), .S(n209), 
        .Z(n2865) );
  MUX2_X1 U1899 ( .A(\REGISTERS[1][21] ), .B(\REGISTERS[17][21] ), .S(n209), 
        .Z(n2866) );
  MUX2_X1 U1900 ( .A(n2866), .B(n2865), .S(n173), .Z(n2867) );
  MUX2_X1 U1901 ( .A(n2867), .B(n2864), .S(n155), .Z(n2868) );
  MUX2_X1 U1902 ( .A(\REGISTERS[12][21] ), .B(\REGISTERS[28][21] ), .S(n210), 
        .Z(n2869) );
  MUX2_X1 U1903 ( .A(\REGISTERS[4][21] ), .B(\REGISTERS[20][21] ), .S(n210), 
        .Z(n2870) );
  MUX2_X1 U1904 ( .A(n2870), .B(n2869), .S(n173), .Z(n2871) );
  MUX2_X1 U1905 ( .A(\REGISTERS[8][21] ), .B(\REGISTERS[24][21] ), .S(n210), 
        .Z(n2872) );
  MUX2_X1 U1906 ( .A(\REGISTERS[0][21] ), .B(\REGISTERS[16][21] ), .S(n210), 
        .Z(n2873) );
  MUX2_X1 U1907 ( .A(n2873), .B(n2872), .S(n173), .Z(n2874) );
  MUX2_X1 U1908 ( .A(n2874), .B(n2871), .S(n155), .Z(n2875) );
  MUX2_X1 U1909 ( .A(n2875), .B(n2868), .S(ADD_RD1[0]), .Z(n2876) );
  MUX2_X1 U1910 ( .A(n2876), .B(n2861), .S(ADD_RD1[1]), .Z(N400) );
  MUX2_X1 U1911 ( .A(\REGISTERS[15][22] ), .B(\REGISTERS[31][22] ), .S(n210), 
        .Z(n2877) );
  MUX2_X1 U1912 ( .A(\REGISTERS[7][22] ), .B(\REGISTERS[23][22] ), .S(n210), 
        .Z(n2878) );
  MUX2_X1 U1913 ( .A(n2878), .B(n2877), .S(n173), .Z(n2879) );
  MUX2_X1 U1914 ( .A(\REGISTERS[11][22] ), .B(\REGISTERS[27][22] ), .S(n210), 
        .Z(n2880) );
  MUX2_X1 U1915 ( .A(\REGISTERS[3][22] ), .B(\REGISTERS[19][22] ), .S(n210), 
        .Z(n2881) );
  MUX2_X1 U1916 ( .A(n2881), .B(n2880), .S(n173), .Z(n2882) );
  MUX2_X1 U1917 ( .A(n2882), .B(n2879), .S(n155), .Z(n2883) );
  MUX2_X1 U1918 ( .A(\REGISTERS[14][22] ), .B(\REGISTERS[30][22] ), .S(n210), 
        .Z(n2884) );
  MUX2_X1 U1919 ( .A(\REGISTERS[6][22] ), .B(\REGISTERS[22][22] ), .S(n210), 
        .Z(n2885) );
  MUX2_X1 U1920 ( .A(n2885), .B(n2884), .S(n173), .Z(n2886) );
  MUX2_X1 U1921 ( .A(\REGISTERS[10][22] ), .B(\REGISTERS[26][22] ), .S(n210), 
        .Z(n2887) );
  MUX2_X1 U1922 ( .A(\REGISTERS[2][22] ), .B(\REGISTERS[18][22] ), .S(n210), 
        .Z(n2888) );
  MUX2_X1 U1923 ( .A(n2888), .B(n2887), .S(n173), .Z(n2889) );
  MUX2_X1 U1924 ( .A(n2889), .B(n2886), .S(n155), .Z(n2890) );
  MUX2_X1 U1925 ( .A(n2890), .B(n2883), .S(ADD_RD1[0]), .Z(n2891) );
  MUX2_X1 U1926 ( .A(\REGISTERS[13][22] ), .B(\REGISTERS[29][22] ), .S(n211), 
        .Z(n2892) );
  MUX2_X1 U1927 ( .A(\REGISTERS[5][22] ), .B(\REGISTERS[21][22] ), .S(n211), 
        .Z(n2893) );
  MUX2_X1 U1928 ( .A(n2893), .B(n2892), .S(n174), .Z(n2894) );
  MUX2_X1 U1929 ( .A(\REGISTERS[9][22] ), .B(\REGISTERS[25][22] ), .S(n211), 
        .Z(n2895) );
  MUX2_X1 U1930 ( .A(\REGISTERS[1][22] ), .B(\REGISTERS[17][22] ), .S(n211), 
        .Z(n2896) );
  MUX2_X1 U1931 ( .A(n2896), .B(n2895), .S(n174), .Z(n2897) );
  MUX2_X1 U1932 ( .A(n2897), .B(n2894), .S(n155), .Z(n2898) );
  MUX2_X1 U1933 ( .A(\REGISTERS[12][22] ), .B(\REGISTERS[28][22] ), .S(n211), 
        .Z(n2899) );
  MUX2_X1 U1934 ( .A(\REGISTERS[4][22] ), .B(\REGISTERS[20][22] ), .S(n211), 
        .Z(n2900) );
  MUX2_X1 U1935 ( .A(n2900), .B(n2899), .S(n174), .Z(n2901) );
  MUX2_X1 U1936 ( .A(\REGISTERS[8][22] ), .B(\REGISTERS[24][22] ), .S(n211), 
        .Z(n2902) );
  MUX2_X1 U1937 ( .A(\REGISTERS[0][22] ), .B(\REGISTERS[16][22] ), .S(n211), 
        .Z(n2903) );
  MUX2_X1 U1938 ( .A(n2903), .B(n2902), .S(n174), .Z(n2904) );
  MUX2_X1 U1939 ( .A(n2904), .B(n2901), .S(n155), .Z(n2905) );
  MUX2_X1 U1940 ( .A(n2905), .B(n2898), .S(ADD_RD1[0]), .Z(n2906) );
  MUX2_X1 U1941 ( .A(n2906), .B(n2891), .S(ADD_RD1[1]), .Z(N401) );
  MUX2_X1 U1942 ( .A(\REGISTERS[15][23] ), .B(\REGISTERS[31][23] ), .S(n211), 
        .Z(n2907) );
  MUX2_X1 U1943 ( .A(\REGISTERS[7][23] ), .B(\REGISTERS[23][23] ), .S(n211), 
        .Z(n2908) );
  MUX2_X1 U1944 ( .A(n2908), .B(n2907), .S(n174), .Z(n2909) );
  MUX2_X1 U1945 ( .A(\REGISTERS[11][23] ), .B(\REGISTERS[27][23] ), .S(n211), 
        .Z(n2910) );
  MUX2_X1 U1946 ( .A(\REGISTERS[3][23] ), .B(\REGISTERS[19][23] ), .S(n211), 
        .Z(n2911) );
  MUX2_X1 U1947 ( .A(n2911), .B(n2910), .S(n174), .Z(n2912) );
  MUX2_X1 U1948 ( .A(n2912), .B(n2909), .S(n155), .Z(n2913) );
  MUX2_X1 U1949 ( .A(\REGISTERS[14][23] ), .B(\REGISTERS[30][23] ), .S(n212), 
        .Z(n2914) );
  MUX2_X1 U1950 ( .A(\REGISTERS[6][23] ), .B(\REGISTERS[22][23] ), .S(n212), 
        .Z(n2915) );
  MUX2_X1 U1951 ( .A(n2915), .B(n2914), .S(n174), .Z(n2916) );
  MUX2_X1 U1952 ( .A(\REGISTERS[10][23] ), .B(\REGISTERS[26][23] ), .S(n212), 
        .Z(n2917) );
  MUX2_X1 U1953 ( .A(\REGISTERS[2][23] ), .B(\REGISTERS[18][23] ), .S(n212), 
        .Z(n2918) );
  MUX2_X1 U1954 ( .A(n2918), .B(n2917), .S(n174), .Z(n2919) );
  MUX2_X1 U1955 ( .A(n2919), .B(n2916), .S(n155), .Z(n2920) );
  MUX2_X1 U1956 ( .A(n2920), .B(n2913), .S(ADD_RD1[0]), .Z(n2921) );
  MUX2_X1 U1957 ( .A(\REGISTERS[13][23] ), .B(\REGISTERS[29][23] ), .S(n212), 
        .Z(n2922) );
  MUX2_X1 U1958 ( .A(\REGISTERS[5][23] ), .B(\REGISTERS[21][23] ), .S(n212), 
        .Z(n2923) );
  MUX2_X1 U1959 ( .A(n2923), .B(n2922), .S(n174), .Z(n2924) );
  MUX2_X1 U1960 ( .A(\REGISTERS[9][23] ), .B(\REGISTERS[25][23] ), .S(n212), 
        .Z(n2925) );
  MUX2_X1 U1961 ( .A(\REGISTERS[1][23] ), .B(\REGISTERS[17][23] ), .S(n212), 
        .Z(n2926) );
  MUX2_X1 U1962 ( .A(n2926), .B(n2925), .S(n174), .Z(n2927) );
  MUX2_X1 U1963 ( .A(n2927), .B(n2924), .S(n155), .Z(n2928) );
  MUX2_X1 U1964 ( .A(\REGISTERS[12][23] ), .B(\REGISTERS[28][23] ), .S(n212), 
        .Z(n2929) );
  MUX2_X1 U1965 ( .A(\REGISTERS[4][23] ), .B(\REGISTERS[20][23] ), .S(n212), 
        .Z(n2930) );
  MUX2_X1 U1966 ( .A(n2930), .B(n2929), .S(n174), .Z(n2931) );
  MUX2_X1 U1967 ( .A(\REGISTERS[8][23] ), .B(\REGISTERS[24][23] ), .S(n212), 
        .Z(n2932) );
  MUX2_X1 U1968 ( .A(\REGISTERS[0][23] ), .B(\REGISTERS[16][23] ), .S(n212), 
        .Z(n2933) );
  MUX2_X1 U1969 ( .A(n2933), .B(n2932), .S(n174), .Z(n2934) );
  MUX2_X1 U1970 ( .A(n2934), .B(n2931), .S(n155), .Z(n2935) );
  MUX2_X1 U1971 ( .A(n2935), .B(n2928), .S(ADD_RD1[0]), .Z(n2936) );
  MUX2_X1 U1972 ( .A(n2936), .B(n2921), .S(ADD_RD1[1]), .Z(N402) );
  MUX2_X1 U1973 ( .A(\REGISTERS[15][24] ), .B(\REGISTERS[31][24] ), .S(n213), 
        .Z(n2937) );
  MUX2_X1 U1974 ( .A(\REGISTERS[7][24] ), .B(\REGISTERS[23][24] ), .S(n213), 
        .Z(n2938) );
  MUX2_X1 U1975 ( .A(n2938), .B(n2937), .S(n175), .Z(n2939) );
  MUX2_X1 U1976 ( .A(\REGISTERS[11][24] ), .B(\REGISTERS[27][24] ), .S(n213), 
        .Z(n2940) );
  MUX2_X1 U1977 ( .A(\REGISTERS[3][24] ), .B(\REGISTERS[19][24] ), .S(n213), 
        .Z(n2941) );
  MUX2_X1 U1978 ( .A(n2941), .B(n2940), .S(n175), .Z(n2942) );
  MUX2_X1 U1979 ( .A(n2942), .B(n2939), .S(n156), .Z(n2943) );
  MUX2_X1 U1980 ( .A(\REGISTERS[14][24] ), .B(\REGISTERS[30][24] ), .S(n213), 
        .Z(n2944) );
  MUX2_X1 U1981 ( .A(\REGISTERS[6][24] ), .B(\REGISTERS[22][24] ), .S(n213), 
        .Z(n2945) );
  MUX2_X1 U1982 ( .A(n2945), .B(n2944), .S(n175), .Z(n2946) );
  MUX2_X1 U1983 ( .A(\REGISTERS[10][24] ), .B(\REGISTERS[26][24] ), .S(n213), 
        .Z(n2947) );
  MUX2_X1 U1984 ( .A(\REGISTERS[2][24] ), .B(\REGISTERS[18][24] ), .S(n213), 
        .Z(n2948) );
  MUX2_X1 U1985 ( .A(n2948), .B(n2947), .S(n175), .Z(n2949) );
  MUX2_X1 U1986 ( .A(n2949), .B(n2946), .S(n156), .Z(n2950) );
  MUX2_X1 U1987 ( .A(n2950), .B(n2943), .S(ADD_RD1[0]), .Z(n2951) );
  MUX2_X1 U1988 ( .A(\REGISTERS[13][24] ), .B(\REGISTERS[29][24] ), .S(n213), 
        .Z(n2952) );
  MUX2_X1 U1989 ( .A(\REGISTERS[5][24] ), .B(\REGISTERS[21][24] ), .S(n213), 
        .Z(n2953) );
  MUX2_X1 U1990 ( .A(n2953), .B(n2952), .S(n175), .Z(n2954) );
  MUX2_X1 U1991 ( .A(\REGISTERS[9][24] ), .B(\REGISTERS[25][24] ), .S(n213), 
        .Z(n2955) );
  MUX2_X1 U1992 ( .A(\REGISTERS[1][24] ), .B(\REGISTERS[17][24] ), .S(n213), 
        .Z(n2956) );
  MUX2_X1 U1993 ( .A(n2956), .B(n2955), .S(n175), .Z(n2957) );
  MUX2_X1 U1994 ( .A(n2957), .B(n2954), .S(n156), .Z(n2958) );
  MUX2_X1 U1995 ( .A(\REGISTERS[12][24] ), .B(\REGISTERS[28][24] ), .S(n214), 
        .Z(n2959) );
  MUX2_X1 U1996 ( .A(\REGISTERS[4][24] ), .B(\REGISTERS[20][24] ), .S(n214), 
        .Z(n2960) );
  MUX2_X1 U1997 ( .A(n2960), .B(n2959), .S(n175), .Z(n2961) );
  MUX2_X1 U1998 ( .A(\REGISTERS[8][24] ), .B(\REGISTERS[24][24] ), .S(n214), 
        .Z(n2962) );
  MUX2_X1 U1999 ( .A(\REGISTERS[0][24] ), .B(\REGISTERS[16][24] ), .S(n214), 
        .Z(n2963) );
  MUX2_X1 U2000 ( .A(n2963), .B(n2962), .S(n175), .Z(n2964) );
  MUX2_X1 U2001 ( .A(n2964), .B(n2961), .S(n156), .Z(n2965) );
  MUX2_X1 U2002 ( .A(n2965), .B(n2958), .S(ADD_RD1[0]), .Z(n2966) );
  MUX2_X1 U2003 ( .A(n2966), .B(n2951), .S(ADD_RD1[1]), .Z(N403) );
  MUX2_X1 U2004 ( .A(\REGISTERS[15][25] ), .B(\REGISTERS[31][25] ), .S(n214), 
        .Z(n2967) );
  MUX2_X1 U2005 ( .A(\REGISTERS[7][25] ), .B(\REGISTERS[23][25] ), .S(n214), 
        .Z(n2968) );
  MUX2_X1 U2006 ( .A(n2968), .B(n2967), .S(n175), .Z(n2969) );
  MUX2_X1 U2007 ( .A(\REGISTERS[11][25] ), .B(\REGISTERS[27][25] ), .S(n214), 
        .Z(n2970) );
  MUX2_X1 U2008 ( .A(\REGISTERS[3][25] ), .B(\REGISTERS[19][25] ), .S(n214), 
        .Z(n2971) );
  MUX2_X1 U2009 ( .A(n2971), .B(n2970), .S(n175), .Z(n2972) );
  MUX2_X1 U2010 ( .A(n2972), .B(n2969), .S(n156), .Z(n2973) );
  MUX2_X1 U2011 ( .A(\REGISTERS[14][25] ), .B(\REGISTERS[30][25] ), .S(n214), 
        .Z(n2974) );
  MUX2_X1 U2012 ( .A(\REGISTERS[6][25] ), .B(\REGISTERS[22][25] ), .S(n214), 
        .Z(n2975) );
  MUX2_X1 U2013 ( .A(n2975), .B(n2974), .S(n175), .Z(n2976) );
  MUX2_X1 U2014 ( .A(\REGISTERS[10][25] ), .B(\REGISTERS[26][25] ), .S(n214), 
        .Z(n2977) );
  MUX2_X1 U2015 ( .A(\REGISTERS[2][25] ), .B(\REGISTERS[18][25] ), .S(n214), 
        .Z(n2978) );
  MUX2_X1 U2016 ( .A(n2978), .B(n2977), .S(n175), .Z(n2979) );
  MUX2_X1 U2017 ( .A(n2979), .B(n2976), .S(n156), .Z(n2980) );
  MUX2_X1 U2018 ( .A(n2980), .B(n2973), .S(ADD_RD1[0]), .Z(n2981) );
  MUX2_X1 U2019 ( .A(\REGISTERS[13][25] ), .B(\REGISTERS[29][25] ), .S(n215), 
        .Z(n2982) );
  MUX2_X1 U2020 ( .A(\REGISTERS[5][25] ), .B(\REGISTERS[21][25] ), .S(n215), 
        .Z(n2983) );
  MUX2_X1 U2021 ( .A(n2983), .B(n2982), .S(n176), .Z(n2984) );
  MUX2_X1 U2022 ( .A(\REGISTERS[9][25] ), .B(\REGISTERS[25][25] ), .S(n215), 
        .Z(n2985) );
  MUX2_X1 U2023 ( .A(\REGISTERS[1][25] ), .B(\REGISTERS[17][25] ), .S(n215), 
        .Z(n2986) );
  MUX2_X1 U2024 ( .A(n2986), .B(n2985), .S(n176), .Z(n2987) );
  MUX2_X1 U2025 ( .A(n2987), .B(n2984), .S(n156), .Z(n2988) );
  MUX2_X1 U2026 ( .A(\REGISTERS[12][25] ), .B(\REGISTERS[28][25] ), .S(n215), 
        .Z(n2989) );
  MUX2_X1 U2027 ( .A(\REGISTERS[4][25] ), .B(\REGISTERS[20][25] ), .S(n215), 
        .Z(n2990) );
  MUX2_X1 U2028 ( .A(n2990), .B(n2989), .S(n176), .Z(n2991) );
  MUX2_X1 U2029 ( .A(\REGISTERS[8][25] ), .B(\REGISTERS[24][25] ), .S(n215), 
        .Z(n2992) );
  MUX2_X1 U2030 ( .A(\REGISTERS[0][25] ), .B(\REGISTERS[16][25] ), .S(n215), 
        .Z(n2993) );
  MUX2_X1 U2031 ( .A(n2993), .B(n2992), .S(n176), .Z(n2994) );
  MUX2_X1 U2032 ( .A(n2994), .B(n2991), .S(n156), .Z(n2995) );
  MUX2_X1 U2033 ( .A(n2995), .B(n2988), .S(ADD_RD1[0]), .Z(n2996) );
  MUX2_X1 U2034 ( .A(n2996), .B(n2981), .S(ADD_RD1[1]), .Z(N404) );
  MUX2_X1 U2035 ( .A(\REGISTERS[15][26] ), .B(\REGISTERS[31][26] ), .S(n215), 
        .Z(n2997) );
  MUX2_X1 U2036 ( .A(\REGISTERS[7][26] ), .B(\REGISTERS[23][26] ), .S(n215), 
        .Z(n2998) );
  MUX2_X1 U2037 ( .A(n2998), .B(n2997), .S(n176), .Z(n2999) );
  MUX2_X1 U2038 ( .A(\REGISTERS[11][26] ), .B(\REGISTERS[27][26] ), .S(n215), 
        .Z(n3000) );
  MUX2_X1 U2039 ( .A(\REGISTERS[3][26] ), .B(\REGISTERS[19][26] ), .S(n215), 
        .Z(n3001) );
  MUX2_X1 U2040 ( .A(n3001), .B(n3000), .S(n176), .Z(n3002) );
  MUX2_X1 U2041 ( .A(n3002), .B(n2999), .S(n156), .Z(n3003) );
  MUX2_X1 U2042 ( .A(\REGISTERS[14][26] ), .B(\REGISTERS[30][26] ), .S(n216), 
        .Z(n3004) );
  MUX2_X1 U2043 ( .A(\REGISTERS[6][26] ), .B(\REGISTERS[22][26] ), .S(n216), 
        .Z(n3005) );
  MUX2_X1 U2044 ( .A(n3005), .B(n3004), .S(n176), .Z(n3006) );
  MUX2_X1 U2045 ( .A(\REGISTERS[10][26] ), .B(\REGISTERS[26][26] ), .S(n216), 
        .Z(n3007) );
  MUX2_X1 U2046 ( .A(\REGISTERS[2][26] ), .B(\REGISTERS[18][26] ), .S(n216), 
        .Z(n3008) );
  MUX2_X1 U2047 ( .A(n3008), .B(n3007), .S(n176), .Z(n3009) );
  MUX2_X1 U2048 ( .A(n3009), .B(n3006), .S(n156), .Z(n3010) );
  MUX2_X1 U2049 ( .A(n3010), .B(n3003), .S(ADD_RD1[0]), .Z(n3011) );
  MUX2_X1 U2050 ( .A(\REGISTERS[13][26] ), .B(\REGISTERS[29][26] ), .S(n216), 
        .Z(n3012) );
  MUX2_X1 U2051 ( .A(\REGISTERS[5][26] ), .B(\REGISTERS[21][26] ), .S(n216), 
        .Z(n3013) );
  MUX2_X1 U2052 ( .A(n3013), .B(n3012), .S(n176), .Z(n3014) );
  MUX2_X1 U2053 ( .A(\REGISTERS[9][26] ), .B(\REGISTERS[25][26] ), .S(n216), 
        .Z(n3015) );
  MUX2_X1 U2054 ( .A(\REGISTERS[1][26] ), .B(\REGISTERS[17][26] ), .S(n216), 
        .Z(n3016) );
  MUX2_X1 U2055 ( .A(n3016), .B(n3015), .S(n176), .Z(n3017) );
  MUX2_X1 U2056 ( .A(n3017), .B(n3014), .S(n156), .Z(n3018) );
  MUX2_X1 U2057 ( .A(\REGISTERS[12][26] ), .B(\REGISTERS[28][26] ), .S(n216), 
        .Z(n3019) );
  MUX2_X1 U2058 ( .A(\REGISTERS[4][26] ), .B(\REGISTERS[20][26] ), .S(n216), 
        .Z(n3020) );
  MUX2_X1 U2059 ( .A(n3020), .B(n3019), .S(n176), .Z(n3021) );
  MUX2_X1 U2060 ( .A(\REGISTERS[8][26] ), .B(\REGISTERS[24][26] ), .S(n216), 
        .Z(n3022) );
  MUX2_X1 U2061 ( .A(\REGISTERS[0][26] ), .B(\REGISTERS[16][26] ), .S(n216), 
        .Z(n3023) );
  MUX2_X1 U2062 ( .A(n3023), .B(n3022), .S(n176), .Z(n3024) );
  MUX2_X1 U2063 ( .A(n3024), .B(n3021), .S(n156), .Z(n3025) );
  MUX2_X1 U2064 ( .A(n3025), .B(n3018), .S(ADD_RD1[0]), .Z(n3026) );
  MUX2_X1 U2065 ( .A(n3026), .B(n3011), .S(ADD_RD1[1]), .Z(N405) );
  MUX2_X1 U2066 ( .A(\REGISTERS[15][27] ), .B(\REGISTERS[31][27] ), .S(n217), 
        .Z(n3027) );
  MUX2_X1 U2067 ( .A(\REGISTERS[7][27] ), .B(\REGISTERS[23][27] ), .S(n217), 
        .Z(n3028) );
  MUX2_X1 U2068 ( .A(n3028), .B(n3027), .S(n177), .Z(n3029) );
  MUX2_X1 U2069 ( .A(\REGISTERS[11][27] ), .B(\REGISTERS[27][27] ), .S(n217), 
        .Z(n3030) );
  MUX2_X1 U2070 ( .A(\REGISTERS[3][27] ), .B(\REGISTERS[19][27] ), .S(n217), 
        .Z(n3031) );
  MUX2_X1 U2071 ( .A(n3031), .B(n3030), .S(n177), .Z(n3032) );
  MUX2_X1 U2072 ( .A(n3032), .B(n3029), .S(n157), .Z(n3033) );
  MUX2_X1 U2073 ( .A(\REGISTERS[14][27] ), .B(\REGISTERS[30][27] ), .S(n217), 
        .Z(n3034) );
  MUX2_X1 U2074 ( .A(\REGISTERS[6][27] ), .B(\REGISTERS[22][27] ), .S(n217), 
        .Z(n3035) );
  MUX2_X1 U2075 ( .A(n3035), .B(n3034), .S(n177), .Z(n3036) );
  MUX2_X1 U2076 ( .A(\REGISTERS[10][27] ), .B(\REGISTERS[26][27] ), .S(n217), 
        .Z(n3037) );
  MUX2_X1 U2077 ( .A(\REGISTERS[2][27] ), .B(\REGISTERS[18][27] ), .S(n217), 
        .Z(n3038) );
  MUX2_X1 U2078 ( .A(n3038), .B(n3037), .S(n177), .Z(n3039) );
  MUX2_X1 U2079 ( .A(n3039), .B(n3036), .S(n157), .Z(n3040) );
  MUX2_X1 U2080 ( .A(n3040), .B(n3033), .S(ADD_RD1[0]), .Z(n3041) );
  MUX2_X1 U2081 ( .A(\REGISTERS[13][27] ), .B(\REGISTERS[29][27] ), .S(n217), 
        .Z(n3042) );
  MUX2_X1 U2082 ( .A(\REGISTERS[5][27] ), .B(\REGISTERS[21][27] ), .S(n217), 
        .Z(n3043) );
  MUX2_X1 U2083 ( .A(n3043), .B(n3042), .S(n177), .Z(n3044) );
  MUX2_X1 U2084 ( .A(\REGISTERS[9][27] ), .B(\REGISTERS[25][27] ), .S(n217), 
        .Z(n3045) );
  MUX2_X1 U2085 ( .A(\REGISTERS[1][27] ), .B(\REGISTERS[17][27] ), .S(n217), 
        .Z(n3046) );
  MUX2_X1 U2086 ( .A(n3046), .B(n3045), .S(n177), .Z(n3047) );
  MUX2_X1 U2087 ( .A(n3047), .B(n3044), .S(n157), .Z(n3048) );
  MUX2_X1 U2088 ( .A(\REGISTERS[12][27] ), .B(\REGISTERS[28][27] ), .S(n218), 
        .Z(n3049) );
  MUX2_X1 U2089 ( .A(\REGISTERS[4][27] ), .B(\REGISTERS[20][27] ), .S(n218), 
        .Z(n3050) );
  MUX2_X1 U2090 ( .A(n3050), .B(n3049), .S(n177), .Z(n3051) );
  MUX2_X1 U2091 ( .A(\REGISTERS[8][27] ), .B(\REGISTERS[24][27] ), .S(n218), 
        .Z(n3052) );
  MUX2_X1 U2092 ( .A(\REGISTERS[0][27] ), .B(\REGISTERS[16][27] ), .S(n218), 
        .Z(n3053) );
  MUX2_X1 U2093 ( .A(n3053), .B(n3052), .S(n177), .Z(n3054) );
  MUX2_X1 U2094 ( .A(n3054), .B(n3051), .S(n157), .Z(n3055) );
  MUX2_X1 U2095 ( .A(n3055), .B(n3048), .S(ADD_RD1[0]), .Z(n3056) );
  MUX2_X1 U2096 ( .A(n3056), .B(n3041), .S(ADD_RD1[1]), .Z(N406) );
  MUX2_X1 U2097 ( .A(\REGISTERS[15][28] ), .B(\REGISTERS[31][28] ), .S(n218), 
        .Z(n3057) );
  MUX2_X1 U2098 ( .A(\REGISTERS[7][28] ), .B(\REGISTERS[23][28] ), .S(n218), 
        .Z(n3058) );
  MUX2_X1 U2099 ( .A(n3058), .B(n3057), .S(n177), .Z(n3059) );
  MUX2_X1 U2100 ( .A(\REGISTERS[11][28] ), .B(\REGISTERS[27][28] ), .S(n218), 
        .Z(n3060) );
  MUX2_X1 U2101 ( .A(\REGISTERS[3][28] ), .B(\REGISTERS[19][28] ), .S(n218), 
        .Z(n3061) );
  MUX2_X1 U2102 ( .A(n3061), .B(n3060), .S(n177), .Z(n3062) );
  MUX2_X1 U2103 ( .A(n3062), .B(n3059), .S(n157), .Z(n3063) );
  MUX2_X1 U2104 ( .A(\REGISTERS[14][28] ), .B(\REGISTERS[30][28] ), .S(n218), 
        .Z(n3064) );
  MUX2_X1 U2105 ( .A(\REGISTERS[6][28] ), .B(\REGISTERS[22][28] ), .S(n218), 
        .Z(n3065) );
  MUX2_X1 U2106 ( .A(n3065), .B(n3064), .S(n177), .Z(n3066) );
  MUX2_X1 U2107 ( .A(\REGISTERS[10][28] ), .B(\REGISTERS[26][28] ), .S(n218), 
        .Z(n3067) );
  MUX2_X1 U2108 ( .A(\REGISTERS[2][28] ), .B(\REGISTERS[18][28] ), .S(n218), 
        .Z(n3068) );
  MUX2_X1 U2109 ( .A(n3068), .B(n3067), .S(n177), .Z(n3069) );
  MUX2_X1 U2110 ( .A(n3069), .B(n3066), .S(n157), .Z(n3070) );
  MUX2_X1 U2111 ( .A(n3070), .B(n3063), .S(ADD_RD1[0]), .Z(n3071) );
  MUX2_X1 U2112 ( .A(\REGISTERS[13][28] ), .B(\REGISTERS[29][28] ), .S(n219), 
        .Z(n3072) );
  MUX2_X1 U2113 ( .A(\REGISTERS[5][28] ), .B(\REGISTERS[21][28] ), .S(n219), 
        .Z(n3073) );
  MUX2_X1 U2114 ( .A(n3073), .B(n3072), .S(n178), .Z(n3074) );
  MUX2_X1 U2115 ( .A(\REGISTERS[9][28] ), .B(\REGISTERS[25][28] ), .S(n219), 
        .Z(n3075) );
  MUX2_X1 U2116 ( .A(\REGISTERS[1][28] ), .B(\REGISTERS[17][28] ), .S(n219), 
        .Z(n3076) );
  MUX2_X1 U2117 ( .A(n3076), .B(n3075), .S(n178), .Z(n3077) );
  MUX2_X1 U2118 ( .A(n3077), .B(n3074), .S(n157), .Z(n3078) );
  MUX2_X1 U2119 ( .A(\REGISTERS[12][28] ), .B(\REGISTERS[28][28] ), .S(n219), 
        .Z(n3079) );
  MUX2_X1 U2120 ( .A(\REGISTERS[4][28] ), .B(\REGISTERS[20][28] ), .S(n219), 
        .Z(n3080) );
  MUX2_X1 U2121 ( .A(n3080), .B(n3079), .S(n178), .Z(n3081) );
  MUX2_X1 U2122 ( .A(\REGISTERS[8][28] ), .B(\REGISTERS[24][28] ), .S(n219), 
        .Z(n3082) );
  MUX2_X1 U2123 ( .A(\REGISTERS[0][28] ), .B(\REGISTERS[16][28] ), .S(n219), 
        .Z(n3083) );
  MUX2_X1 U2124 ( .A(n3083), .B(n3082), .S(n178), .Z(n3084) );
  MUX2_X1 U2125 ( .A(n3084), .B(n3081), .S(n157), .Z(n3085) );
  MUX2_X1 U2126 ( .A(n3085), .B(n3078), .S(ADD_RD1[0]), .Z(n3086) );
  MUX2_X1 U2127 ( .A(n3086), .B(n3071), .S(ADD_RD1[1]), .Z(N407) );
  MUX2_X1 U2128 ( .A(\REGISTERS[15][29] ), .B(\REGISTERS[31][29] ), .S(n219), 
        .Z(n3087) );
  MUX2_X1 U2129 ( .A(\REGISTERS[7][29] ), .B(\REGISTERS[23][29] ), .S(n219), 
        .Z(n3088) );
  MUX2_X1 U2130 ( .A(n3088), .B(n3087), .S(n178), .Z(n3089) );
  MUX2_X1 U2131 ( .A(\REGISTERS[11][29] ), .B(\REGISTERS[27][29] ), .S(n219), 
        .Z(n3090) );
  MUX2_X1 U2132 ( .A(\REGISTERS[3][29] ), .B(\REGISTERS[19][29] ), .S(n219), 
        .Z(n3091) );
  MUX2_X1 U2133 ( .A(n3091), .B(n3090), .S(n178), .Z(n3092) );
  MUX2_X1 U2134 ( .A(n3092), .B(n3089), .S(n157), .Z(n3093) );
  MUX2_X1 U2135 ( .A(\REGISTERS[14][29] ), .B(\REGISTERS[30][29] ), .S(n220), 
        .Z(n3094) );
  MUX2_X1 U2136 ( .A(\REGISTERS[6][29] ), .B(\REGISTERS[22][29] ), .S(n220), 
        .Z(n3095) );
  MUX2_X1 U2137 ( .A(n3095), .B(n3094), .S(n178), .Z(n3096) );
  MUX2_X1 U2138 ( .A(\REGISTERS[10][29] ), .B(\REGISTERS[26][29] ), .S(n220), 
        .Z(n3097) );
  MUX2_X1 U2139 ( .A(\REGISTERS[2][29] ), .B(\REGISTERS[18][29] ), .S(n220), 
        .Z(n3098) );
  MUX2_X1 U2140 ( .A(n3098), .B(n3097), .S(n178), .Z(n3099) );
  MUX2_X1 U2141 ( .A(n3099), .B(n3096), .S(n157), .Z(n3100) );
  MUX2_X1 U2142 ( .A(n3100), .B(n3093), .S(ADD_RD1[0]), .Z(n3101) );
  MUX2_X1 U2143 ( .A(\REGISTERS[13][29] ), .B(\REGISTERS[29][29] ), .S(n220), 
        .Z(n3102) );
  MUX2_X1 U2144 ( .A(\REGISTERS[5][29] ), .B(\REGISTERS[21][29] ), .S(n220), 
        .Z(n3103) );
  MUX2_X1 U2145 ( .A(n3103), .B(n3102), .S(n178), .Z(n3104) );
  MUX2_X1 U2146 ( .A(\REGISTERS[9][29] ), .B(\REGISTERS[25][29] ), .S(n220), 
        .Z(n3105) );
  MUX2_X1 U2147 ( .A(\REGISTERS[1][29] ), .B(\REGISTERS[17][29] ), .S(n220), 
        .Z(n3106) );
  MUX2_X1 U2148 ( .A(n3106), .B(n3105), .S(n178), .Z(n3107) );
  MUX2_X1 U2149 ( .A(n3107), .B(n3104), .S(n157), .Z(n3108) );
  MUX2_X1 U2150 ( .A(\REGISTERS[12][29] ), .B(\REGISTERS[28][29] ), .S(n220), 
        .Z(n3109) );
  MUX2_X1 U2151 ( .A(\REGISTERS[4][29] ), .B(\REGISTERS[20][29] ), .S(n220), 
        .Z(n3110) );
  MUX2_X1 U2152 ( .A(n3110), .B(n3109), .S(n178), .Z(n3111) );
  MUX2_X1 U2153 ( .A(\REGISTERS[8][29] ), .B(\REGISTERS[24][29] ), .S(n220), 
        .Z(n3112) );
  MUX2_X1 U2154 ( .A(\REGISTERS[0][29] ), .B(\REGISTERS[16][29] ), .S(n220), 
        .Z(n3113) );
  MUX2_X1 U2155 ( .A(n3113), .B(n3112), .S(n178), .Z(n3114) );
  MUX2_X1 U2156 ( .A(n3114), .B(n3111), .S(n157), .Z(n3115) );
  MUX2_X1 U2157 ( .A(n3115), .B(n3108), .S(ADD_RD1[0]), .Z(n3116) );
  MUX2_X1 U2158 ( .A(n3116), .B(n3101), .S(ADD_RD1[1]), .Z(N408) );
  MUX2_X1 U2159 ( .A(\REGISTERS[15][30] ), .B(\REGISTERS[31][30] ), .S(n221), 
        .Z(n3117) );
  MUX2_X1 U2160 ( .A(\REGISTERS[7][30] ), .B(\REGISTERS[23][30] ), .S(n221), 
        .Z(n3118) );
  MUX2_X1 U2161 ( .A(n3118), .B(n3117), .S(n179), .Z(n3119) );
  MUX2_X1 U2162 ( .A(\REGISTERS[11][30] ), .B(\REGISTERS[27][30] ), .S(n221), 
        .Z(n3120) );
  MUX2_X1 U2163 ( .A(\REGISTERS[3][30] ), .B(\REGISTERS[19][30] ), .S(n221), 
        .Z(n3121) );
  MUX2_X1 U2164 ( .A(n3121), .B(n3120), .S(n179), .Z(n3122) );
  MUX2_X1 U2165 ( .A(n3122), .B(n3119), .S(n158), .Z(n3123) );
  MUX2_X1 U2166 ( .A(\REGISTERS[14][30] ), .B(\REGISTERS[30][30] ), .S(n221), 
        .Z(n3124) );
  MUX2_X1 U2167 ( .A(\REGISTERS[6][30] ), .B(\REGISTERS[22][30] ), .S(n221), 
        .Z(n3125) );
  MUX2_X1 U2168 ( .A(n3125), .B(n3124), .S(n179), .Z(n3126) );
  MUX2_X1 U2169 ( .A(\REGISTERS[10][30] ), .B(\REGISTERS[26][30] ), .S(n221), 
        .Z(n3127) );
  MUX2_X1 U2170 ( .A(\REGISTERS[2][30] ), .B(\REGISTERS[18][30] ), .S(n221), 
        .Z(n3128) );
  MUX2_X1 U2171 ( .A(n3128), .B(n3127), .S(n179), .Z(n3129) );
  MUX2_X1 U2172 ( .A(n3129), .B(n3126), .S(n158), .Z(n3130) );
  MUX2_X1 U2173 ( .A(n3130), .B(n3123), .S(ADD_RD1[0]), .Z(n3131) );
  MUX2_X1 U2174 ( .A(\REGISTERS[13][30] ), .B(\REGISTERS[29][30] ), .S(n221), 
        .Z(n3132) );
  MUX2_X1 U2175 ( .A(\REGISTERS[5][30] ), .B(\REGISTERS[21][30] ), .S(n221), 
        .Z(n3133) );
  MUX2_X1 U2176 ( .A(n3133), .B(n3132), .S(n179), .Z(n3134) );
  MUX2_X1 U2177 ( .A(\REGISTERS[9][30] ), .B(\REGISTERS[25][30] ), .S(n221), 
        .Z(n3135) );
  MUX2_X1 U2178 ( .A(\REGISTERS[1][30] ), .B(\REGISTERS[17][30] ), .S(n221), 
        .Z(n3136) );
  MUX2_X1 U2179 ( .A(n3136), .B(n3135), .S(n179), .Z(n3137) );
  MUX2_X1 U2180 ( .A(n3137), .B(n3134), .S(n158), .Z(n3138) );
  MUX2_X1 U2181 ( .A(\REGISTERS[12][30] ), .B(\REGISTERS[28][30] ), .S(n222), 
        .Z(n3139) );
  MUX2_X1 U2182 ( .A(\REGISTERS[4][30] ), .B(\REGISTERS[20][30] ), .S(n222), 
        .Z(n3140) );
  MUX2_X1 U2183 ( .A(n3140), .B(n3139), .S(n179), .Z(n3141) );
  MUX2_X1 U2184 ( .A(\REGISTERS[8][30] ), .B(\REGISTERS[24][30] ), .S(n222), 
        .Z(n3142) );
  MUX2_X1 U2185 ( .A(\REGISTERS[0][30] ), .B(\REGISTERS[16][30] ), .S(n222), 
        .Z(n3143) );
  MUX2_X1 U2186 ( .A(n3143), .B(n3142), .S(n179), .Z(n3144) );
  MUX2_X1 U2187 ( .A(n3144), .B(n3141), .S(n158), .Z(n3145) );
  MUX2_X1 U2188 ( .A(n3145), .B(n3138), .S(ADD_RD1[0]), .Z(n3146) );
  MUX2_X1 U2189 ( .A(n3146), .B(n3131), .S(ADD_RD1[1]), .Z(N409) );
  MUX2_X1 U2190 ( .A(\REGISTERS[15][31] ), .B(\REGISTERS[31][31] ), .S(n222), 
        .Z(n3147) );
  MUX2_X1 U2191 ( .A(\REGISTERS[7][31] ), .B(\REGISTERS[23][31] ), .S(n222), 
        .Z(n3148) );
  MUX2_X1 U2192 ( .A(n3148), .B(n3147), .S(n179), .Z(n3149) );
  MUX2_X1 U2193 ( .A(\REGISTERS[11][31] ), .B(\REGISTERS[27][31] ), .S(n222), 
        .Z(n3150) );
  MUX2_X1 U2194 ( .A(\REGISTERS[3][31] ), .B(\REGISTERS[19][31] ), .S(n222), 
        .Z(n3151) );
  MUX2_X1 U2195 ( .A(n3151), .B(n3150), .S(n179), .Z(n3152) );
  MUX2_X1 U2196 ( .A(n3152), .B(n3149), .S(n158), .Z(n3153) );
  MUX2_X1 U2197 ( .A(\REGISTERS[14][31] ), .B(\REGISTERS[30][31] ), .S(n222), 
        .Z(n3154) );
  MUX2_X1 U2198 ( .A(\REGISTERS[6][31] ), .B(\REGISTERS[22][31] ), .S(n222), 
        .Z(n3155) );
  MUX2_X1 U2199 ( .A(n3155), .B(n3154), .S(n179), .Z(n3156) );
  MUX2_X1 U2200 ( .A(\REGISTERS[10][31] ), .B(\REGISTERS[26][31] ), .S(n222), 
        .Z(n3157) );
  MUX2_X1 U2201 ( .A(\REGISTERS[2][31] ), .B(\REGISTERS[18][31] ), .S(n222), 
        .Z(n3158) );
  MUX2_X1 U2202 ( .A(n3158), .B(n3157), .S(n179), .Z(n3159) );
  MUX2_X1 U2203 ( .A(n3159), .B(n3156), .S(n158), .Z(n3160) );
  MUX2_X1 U2204 ( .A(n3160), .B(n3153), .S(ADD_RD1[0]), .Z(n3161) );
  MUX2_X1 U2205 ( .A(\REGISTERS[13][31] ), .B(\REGISTERS[29][31] ), .S(n223), 
        .Z(n3162) );
  MUX2_X1 U2206 ( .A(\REGISTERS[5][31] ), .B(\REGISTERS[21][31] ), .S(n223), 
        .Z(n3163) );
  MUX2_X1 U2207 ( .A(n3163), .B(n3162), .S(n180), .Z(n3164) );
  MUX2_X1 U2208 ( .A(\REGISTERS[9][31] ), .B(\REGISTERS[25][31] ), .S(n223), 
        .Z(n3165) );
  MUX2_X1 U2209 ( .A(\REGISTERS[1][31] ), .B(\REGISTERS[17][31] ), .S(n223), 
        .Z(n3166) );
  MUX2_X1 U2210 ( .A(n3166), .B(n3165), .S(n180), .Z(n3167) );
  MUX2_X1 U2211 ( .A(n3167), .B(n3164), .S(n158), .Z(n3168) );
  MUX2_X1 U2212 ( .A(\REGISTERS[12][31] ), .B(\REGISTERS[28][31] ), .S(n223), 
        .Z(n3169) );
  MUX2_X1 U2213 ( .A(\REGISTERS[4][31] ), .B(\REGISTERS[20][31] ), .S(n223), 
        .Z(n3170) );
  MUX2_X1 U2214 ( .A(n3170), .B(n3169), .S(n180), .Z(n3171) );
  MUX2_X1 U2215 ( .A(\REGISTERS[8][31] ), .B(\REGISTERS[24][31] ), .S(n223), 
        .Z(n3172) );
  MUX2_X1 U2216 ( .A(\REGISTERS[0][31] ), .B(\REGISTERS[16][31] ), .S(n223), 
        .Z(n3173) );
  MUX2_X1 U2217 ( .A(n3173), .B(n3172), .S(n180), .Z(n3174) );
  MUX2_X1 U2218 ( .A(n3174), .B(n3171), .S(n158), .Z(n3175) );
  MUX2_X1 U2219 ( .A(n3175), .B(n3168), .S(ADD_RD1[0]), .Z(n3176) );
  MUX2_X1 U2220 ( .A(n3176), .B(n3161), .S(ADD_RD1[1]), .Z(N410) );
  MUX2_X1 U2221 ( .A(\REGISTERS[0][31] ), .B(n3177), .S(n3178), .Z(n2163) );
  MUX2_X1 U2222 ( .A(\REGISTERS[0][30] ), .B(n3179), .S(n3178), .Z(n2162) );
  MUX2_X1 U2223 ( .A(\REGISTERS[0][29] ), .B(n3180), .S(n3178), .Z(n2161) );
  MUX2_X1 U2224 ( .A(\REGISTERS[0][28] ), .B(n3181), .S(n3178), .Z(n2160) );
  MUX2_X1 U2225 ( .A(\REGISTERS[0][27] ), .B(n3182), .S(n3178), .Z(n2159) );
  MUX2_X1 U2226 ( .A(\REGISTERS[0][26] ), .B(n3183), .S(n3178), .Z(n2158) );
  MUX2_X1 U2227 ( .A(\REGISTERS[0][25] ), .B(n3184), .S(n3178), .Z(n2157) );
  MUX2_X1 U2228 ( .A(\REGISTERS[0][24] ), .B(n3185), .S(n3178), .Z(n2156) );
  MUX2_X1 U2229 ( .A(\REGISTERS[0][23] ), .B(n3186), .S(n3178), .Z(n2155) );
  MUX2_X1 U2230 ( .A(\REGISTERS[0][22] ), .B(n3187), .S(n3178), .Z(n2154) );
  MUX2_X1 U2231 ( .A(\REGISTERS[0][21] ), .B(n3188), .S(n3178), .Z(n2153) );
  MUX2_X1 U2232 ( .A(\REGISTERS[0][20] ), .B(n3189), .S(n3178), .Z(n2152) );
  MUX2_X1 U2233 ( .A(\REGISTERS[0][19] ), .B(n3190), .S(n3178), .Z(n2151) );
  MUX2_X1 U2234 ( .A(\REGISTERS[0][18] ), .B(n3191), .S(n3178), .Z(n2150) );
  MUX2_X1 U2235 ( .A(\REGISTERS[0][17] ), .B(n3192), .S(n3178), .Z(n2149) );
  MUX2_X1 U2236 ( .A(\REGISTERS[0][16] ), .B(n3193), .S(n3178), .Z(n2148) );
  MUX2_X1 U2237 ( .A(\REGISTERS[0][15] ), .B(n3194), .S(n3178), .Z(n2147) );
  MUX2_X1 U2238 ( .A(\REGISTERS[0][14] ), .B(n3195), .S(n3178), .Z(n2146) );
  MUX2_X1 U2239 ( .A(\REGISTERS[0][13] ), .B(n3196), .S(n3178), .Z(n2145) );
  MUX2_X1 U2240 ( .A(\REGISTERS[0][12] ), .B(n3197), .S(n3178), .Z(n2144) );
  MUX2_X1 U2241 ( .A(\REGISTERS[0][11] ), .B(n3198), .S(n3178), .Z(n2143) );
  MUX2_X1 U2242 ( .A(\REGISTERS[0][10] ), .B(n3199), .S(n3178), .Z(n2142) );
  MUX2_X1 U2243 ( .A(\REGISTERS[0][9] ), .B(n3200), .S(n3178), .Z(n2141) );
  MUX2_X1 U2244 ( .A(\REGISTERS[0][8] ), .B(n3201), .S(n3178), .Z(n2140) );
  MUX2_X1 U2245 ( .A(\REGISTERS[0][7] ), .B(n3202), .S(n3178), .Z(n2139) );
  MUX2_X1 U2246 ( .A(\REGISTERS[0][6] ), .B(n3203), .S(n3178), .Z(n2138) );
  MUX2_X1 U2247 ( .A(\REGISTERS[0][5] ), .B(n3204), .S(n3178), .Z(n2137) );
  MUX2_X1 U2248 ( .A(\REGISTERS[0][4] ), .B(n3205), .S(n3178), .Z(n2136) );
  MUX2_X1 U2249 ( .A(\REGISTERS[0][3] ), .B(n3206), .S(n3178), .Z(n2135) );
  MUX2_X1 U2250 ( .A(\REGISTERS[0][2] ), .B(n3207), .S(n3178), .Z(n2134) );
  MUX2_X1 U2251 ( .A(\REGISTERS[0][1] ), .B(n3208), .S(n3178), .Z(n2133) );
  MUX2_X1 U2252 ( .A(\REGISTERS[0][0] ), .B(n3209), .S(n3178), .Z(n2132) );
  MUX2_X1 U2253 ( .A(\REGISTERS[1][31] ), .B(n3177), .S(n60), .Z(n2131) );
  MUX2_X1 U2254 ( .A(\REGISTERS[1][30] ), .B(n3179), .S(n60), .Z(n2130) );
  MUX2_X1 U2255 ( .A(\REGISTERS[1][29] ), .B(n3180), .S(n60), .Z(n2129) );
  MUX2_X1 U2256 ( .A(\REGISTERS[1][28] ), .B(n3181), .S(n60), .Z(n2128) );
  MUX2_X1 U2257 ( .A(\REGISTERS[1][27] ), .B(n3182), .S(n60), .Z(n2127) );
  MUX2_X1 U2258 ( .A(\REGISTERS[1][26] ), .B(n3183), .S(n60), .Z(n2126) );
  MUX2_X1 U2259 ( .A(\REGISTERS[1][25] ), .B(n3184), .S(n60), .Z(n2125) );
  MUX2_X1 U2260 ( .A(\REGISTERS[1][24] ), .B(n3185), .S(n60), .Z(n2124) );
  MUX2_X1 U2261 ( .A(\REGISTERS[1][23] ), .B(n3186), .S(n60), .Z(n2123) );
  MUX2_X1 U2262 ( .A(\REGISTERS[1][22] ), .B(n3187), .S(n60), .Z(n2122) );
  MUX2_X1 U2263 ( .A(\REGISTERS[1][21] ), .B(n3188), .S(n60), .Z(n2121) );
  MUX2_X1 U2264 ( .A(\REGISTERS[1][20] ), .B(n3189), .S(n60), .Z(n2120) );
  MUX2_X1 U2265 ( .A(\REGISTERS[1][19] ), .B(n3190), .S(n60), .Z(n2119) );
  MUX2_X1 U2266 ( .A(\REGISTERS[1][18] ), .B(n3191), .S(n60), .Z(n2118) );
  MUX2_X1 U2267 ( .A(\REGISTERS[1][17] ), .B(n3192), .S(n60), .Z(n2117) );
  MUX2_X1 U2268 ( .A(\REGISTERS[1][16] ), .B(n3193), .S(n60), .Z(n2116) );
  MUX2_X1 U2269 ( .A(\REGISTERS[1][15] ), .B(n3194), .S(n60), .Z(n2115) );
  MUX2_X1 U2270 ( .A(\REGISTERS[1][14] ), .B(n3195), .S(n60), .Z(n2114) );
  MUX2_X1 U2271 ( .A(\REGISTERS[1][13] ), .B(n3196), .S(n60), .Z(n2113) );
  MUX2_X1 U2272 ( .A(\REGISTERS[1][12] ), .B(n3197), .S(n60), .Z(n2112) );
  MUX2_X1 U2273 ( .A(\REGISTERS[1][11] ), .B(n3198), .S(n60), .Z(n2111) );
  MUX2_X1 U2274 ( .A(\REGISTERS[1][10] ), .B(n3199), .S(n60), .Z(n2110) );
  MUX2_X1 U2275 ( .A(\REGISTERS[1][9] ), .B(n3200), .S(n60), .Z(n2109) );
  MUX2_X1 U2276 ( .A(\REGISTERS[1][8] ), .B(n3201), .S(n60), .Z(n2108) );
  MUX2_X1 U2277 ( .A(\REGISTERS[1][7] ), .B(n3202), .S(n60), .Z(n2107) );
  MUX2_X1 U2278 ( .A(\REGISTERS[1][6] ), .B(n3203), .S(n60), .Z(n2106) );
  MUX2_X1 U2279 ( .A(\REGISTERS[1][5] ), .B(n3204), .S(n60), .Z(n2105) );
  MUX2_X1 U2280 ( .A(\REGISTERS[1][4] ), .B(n3205), .S(n60), .Z(n2104) );
  MUX2_X1 U2281 ( .A(\REGISTERS[1][3] ), .B(n3206), .S(n60), .Z(n2103) );
  MUX2_X1 U2282 ( .A(\REGISTERS[1][2] ), .B(n3207), .S(n60), .Z(n2102) );
  MUX2_X1 U2283 ( .A(\REGISTERS[1][1] ), .B(n3208), .S(n60), .Z(n2101) );
  MUX2_X1 U2284 ( .A(\REGISTERS[1][0] ), .B(n3209), .S(n60), .Z(n2100) );
  OAI21_X1 U2285 ( .B1(n3210), .B2(n3214), .A(n3212), .ZN(n3213) );
  MUX2_X1 U2286 ( .A(\REGISTERS[2][31] ), .B(n3177), .S(n62), .Z(n2099) );
  MUX2_X1 U2287 ( .A(\REGISTERS[2][30] ), .B(n3179), .S(n62), .Z(n2098) );
  MUX2_X1 U2288 ( .A(\REGISTERS[2][29] ), .B(n3180), .S(n62), .Z(n2097) );
  MUX2_X1 U2289 ( .A(\REGISTERS[2][28] ), .B(n3181), .S(n62), .Z(n2096) );
  MUX2_X1 U2290 ( .A(\REGISTERS[2][27] ), .B(n3182), .S(n62), .Z(n2095) );
  MUX2_X1 U2291 ( .A(\REGISTERS[2][26] ), .B(n3183), .S(n62), .Z(n2094) );
  MUX2_X1 U2292 ( .A(\REGISTERS[2][25] ), .B(n3184), .S(n62), .Z(n2093) );
  MUX2_X1 U2293 ( .A(\REGISTERS[2][24] ), .B(n3185), .S(n62), .Z(n2092) );
  MUX2_X1 U2294 ( .A(\REGISTERS[2][23] ), .B(n3186), .S(n62), .Z(n2091) );
  MUX2_X1 U2295 ( .A(\REGISTERS[2][22] ), .B(n3187), .S(n62), .Z(n2090) );
  MUX2_X1 U2296 ( .A(\REGISTERS[2][21] ), .B(n3188), .S(n62), .Z(n2089) );
  MUX2_X1 U2297 ( .A(\REGISTERS[2][20] ), .B(n3189), .S(n62), .Z(n2088) );
  MUX2_X1 U2298 ( .A(\REGISTERS[2][19] ), .B(n3190), .S(n62), .Z(n2087) );
  MUX2_X1 U2299 ( .A(\REGISTERS[2][18] ), .B(n3191), .S(n62), .Z(n2086) );
  MUX2_X1 U2300 ( .A(\REGISTERS[2][17] ), .B(n3192), .S(n62), .Z(n2085) );
  MUX2_X1 U2301 ( .A(\REGISTERS[2][16] ), .B(n3193), .S(n62), .Z(n2084) );
  MUX2_X1 U2302 ( .A(\REGISTERS[2][15] ), .B(n3194), .S(n62), .Z(n2083) );
  MUX2_X1 U2303 ( .A(\REGISTERS[2][14] ), .B(n3195), .S(n62), .Z(n2082) );
  MUX2_X1 U2304 ( .A(\REGISTERS[2][13] ), .B(n3196), .S(n62), .Z(n2081) );
  MUX2_X1 U2305 ( .A(\REGISTERS[2][12] ), .B(n3197), .S(n62), .Z(n2080) );
  MUX2_X1 U2306 ( .A(\REGISTERS[2][11] ), .B(n3198), .S(n62), .Z(n2079) );
  MUX2_X1 U2307 ( .A(\REGISTERS[2][10] ), .B(n3199), .S(n62), .Z(n2078) );
  MUX2_X1 U2308 ( .A(\REGISTERS[2][9] ), .B(n3200), .S(n62), .Z(n2077) );
  MUX2_X1 U2309 ( .A(\REGISTERS[2][8] ), .B(n3201), .S(n62), .Z(n2076) );
  MUX2_X1 U2310 ( .A(\REGISTERS[2][7] ), .B(n3202), .S(n62), .Z(n2075) );
  MUX2_X1 U2311 ( .A(\REGISTERS[2][6] ), .B(n3203), .S(n62), .Z(n2074) );
  MUX2_X1 U2312 ( .A(\REGISTERS[2][5] ), .B(n3204), .S(n62), .Z(n2073) );
  MUX2_X1 U2313 ( .A(\REGISTERS[2][4] ), .B(n3205), .S(n62), .Z(n2072) );
  MUX2_X1 U2314 ( .A(\REGISTERS[2][3] ), .B(n3206), .S(n62), .Z(n2071) );
  MUX2_X1 U2315 ( .A(\REGISTERS[2][2] ), .B(n3207), .S(n62), .Z(n2070) );
  MUX2_X1 U2316 ( .A(\REGISTERS[2][1] ), .B(n3208), .S(n62), .Z(n2069) );
  MUX2_X1 U2317 ( .A(\REGISTERS[2][0] ), .B(n3209), .S(n62), .Z(n2068) );
  OAI21_X1 U2318 ( .B1(n3210), .B2(n3216), .A(n3212), .ZN(n3215) );
  MUX2_X1 U2319 ( .A(\REGISTERS[3][31] ), .B(n3177), .S(n56), .Z(n2067) );
  MUX2_X1 U2320 ( .A(\REGISTERS[3][30] ), .B(n3179), .S(n56), .Z(n2066) );
  MUX2_X1 U2321 ( .A(\REGISTERS[3][29] ), .B(n3180), .S(n56), .Z(n2065) );
  MUX2_X1 U2322 ( .A(\REGISTERS[3][28] ), .B(n3181), .S(n56), .Z(n2064) );
  MUX2_X1 U2323 ( .A(\REGISTERS[3][27] ), .B(n3182), .S(n56), .Z(n2063) );
  MUX2_X1 U2324 ( .A(\REGISTERS[3][26] ), .B(n3183), .S(n56), .Z(n2062) );
  MUX2_X1 U2325 ( .A(\REGISTERS[3][25] ), .B(n3184), .S(n56), .Z(n2061) );
  MUX2_X1 U2326 ( .A(\REGISTERS[3][24] ), .B(n3185), .S(n56), .Z(n2060) );
  MUX2_X1 U2327 ( .A(\REGISTERS[3][23] ), .B(n3186), .S(n56), .Z(n2059) );
  MUX2_X1 U2328 ( .A(\REGISTERS[3][22] ), .B(n3187), .S(n56), .Z(n2058) );
  MUX2_X1 U2329 ( .A(\REGISTERS[3][21] ), .B(n3188), .S(n56), .Z(n2057) );
  MUX2_X1 U2330 ( .A(\REGISTERS[3][20] ), .B(n3189), .S(n56), .Z(n2056) );
  MUX2_X1 U2331 ( .A(\REGISTERS[3][19] ), .B(n3190), .S(n56), .Z(n2055) );
  MUX2_X1 U2332 ( .A(\REGISTERS[3][18] ), .B(n3191), .S(n56), .Z(n2054) );
  MUX2_X1 U2333 ( .A(\REGISTERS[3][17] ), .B(n3192), .S(n56), .Z(n2053) );
  MUX2_X1 U2334 ( .A(\REGISTERS[3][16] ), .B(n3193), .S(n56), .Z(n2052) );
  MUX2_X1 U2335 ( .A(\REGISTERS[3][15] ), .B(n3194), .S(n56), .Z(n2051) );
  MUX2_X1 U2336 ( .A(\REGISTERS[3][14] ), .B(n3195), .S(n56), .Z(n2050) );
  MUX2_X1 U2337 ( .A(\REGISTERS[3][13] ), .B(n3196), .S(n56), .Z(n2049) );
  MUX2_X1 U2338 ( .A(\REGISTERS[3][12] ), .B(n3197), .S(n56), .Z(n2048) );
  MUX2_X1 U2339 ( .A(\REGISTERS[3][11] ), .B(n3198), .S(n56), .Z(n2047) );
  MUX2_X1 U2340 ( .A(\REGISTERS[3][10] ), .B(n3199), .S(n56), .Z(n2046) );
  MUX2_X1 U2341 ( .A(\REGISTERS[3][9] ), .B(n3200), .S(n56), .Z(n2045) );
  MUX2_X1 U2342 ( .A(\REGISTERS[3][8] ), .B(n3201), .S(n56), .Z(n2044) );
  MUX2_X1 U2343 ( .A(\REGISTERS[3][7] ), .B(n3202), .S(n56), .Z(n2043) );
  MUX2_X1 U2344 ( .A(\REGISTERS[3][6] ), .B(n3203), .S(n56), .Z(n2042) );
  MUX2_X1 U2345 ( .A(\REGISTERS[3][5] ), .B(n3204), .S(n56), .Z(n2041) );
  MUX2_X1 U2346 ( .A(\REGISTERS[3][4] ), .B(n3205), .S(n56), .Z(n2040) );
  MUX2_X1 U2347 ( .A(\REGISTERS[3][3] ), .B(n3206), .S(n56), .Z(n2039) );
  MUX2_X1 U2348 ( .A(\REGISTERS[3][2] ), .B(n3207), .S(n56), .Z(n2038) );
  MUX2_X1 U2349 ( .A(\REGISTERS[3][1] ), .B(n3208), .S(n56), .Z(n2037) );
  MUX2_X1 U2350 ( .A(\REGISTERS[3][0] ), .B(n3209), .S(n56), .Z(n2036) );
  OAI21_X1 U2351 ( .B1(n3210), .B2(n3218), .A(n3212), .ZN(n3217) );
  MUX2_X1 U2352 ( .A(\REGISTERS[4][31] ), .B(n3177), .S(n58), .Z(n2035) );
  MUX2_X1 U2353 ( .A(\REGISTERS[4][30] ), .B(n3179), .S(n58), .Z(n2034) );
  MUX2_X1 U2354 ( .A(\REGISTERS[4][29] ), .B(n3180), .S(n58), .Z(n2033) );
  MUX2_X1 U2355 ( .A(\REGISTERS[4][28] ), .B(n3181), .S(n58), .Z(n2032) );
  MUX2_X1 U2356 ( .A(\REGISTERS[4][27] ), .B(n3182), .S(n58), .Z(n2031) );
  MUX2_X1 U2357 ( .A(\REGISTERS[4][26] ), .B(n3183), .S(n58), .Z(n2030) );
  MUX2_X1 U2358 ( .A(\REGISTERS[4][25] ), .B(n3184), .S(n58), .Z(n2029) );
  MUX2_X1 U2359 ( .A(\REGISTERS[4][24] ), .B(n3185), .S(n58), .Z(n2028) );
  MUX2_X1 U2360 ( .A(\REGISTERS[4][23] ), .B(n3186), .S(n58), .Z(n2027) );
  MUX2_X1 U2361 ( .A(\REGISTERS[4][22] ), .B(n3187), .S(n58), .Z(n2026) );
  MUX2_X1 U2362 ( .A(\REGISTERS[4][21] ), .B(n3188), .S(n58), .Z(n2025) );
  MUX2_X1 U2363 ( .A(\REGISTERS[4][20] ), .B(n3189), .S(n58), .Z(n2024) );
  MUX2_X1 U2364 ( .A(\REGISTERS[4][19] ), .B(n3190), .S(n58), .Z(n2023) );
  MUX2_X1 U2365 ( .A(\REGISTERS[4][18] ), .B(n3191), .S(n58), .Z(n2022) );
  MUX2_X1 U2366 ( .A(\REGISTERS[4][17] ), .B(n3192), .S(n58), .Z(n2021) );
  MUX2_X1 U2367 ( .A(\REGISTERS[4][16] ), .B(n3193), .S(n58), .Z(n2020) );
  MUX2_X1 U2368 ( .A(\REGISTERS[4][15] ), .B(n3194), .S(n58), .Z(n2019) );
  MUX2_X1 U2369 ( .A(\REGISTERS[4][14] ), .B(n3195), .S(n58), .Z(n2018) );
  MUX2_X1 U2370 ( .A(\REGISTERS[4][13] ), .B(n3196), .S(n58), .Z(n2017) );
  MUX2_X1 U2371 ( .A(\REGISTERS[4][12] ), .B(n3197), .S(n58), .Z(n2016) );
  MUX2_X1 U2372 ( .A(\REGISTERS[4][11] ), .B(n3198), .S(n58), .Z(n2015) );
  MUX2_X1 U2373 ( .A(\REGISTERS[4][10] ), .B(n3199), .S(n58), .Z(n2014) );
  MUX2_X1 U2374 ( .A(\REGISTERS[4][9] ), .B(n3200), .S(n58), .Z(n2013) );
  MUX2_X1 U2375 ( .A(\REGISTERS[4][8] ), .B(n3201), .S(n58), .Z(n2012) );
  MUX2_X1 U2376 ( .A(\REGISTERS[4][7] ), .B(n3202), .S(n58), .Z(n2011) );
  MUX2_X1 U2377 ( .A(\REGISTERS[4][6] ), .B(n3203), .S(n58), .Z(n2010) );
  MUX2_X1 U2378 ( .A(\REGISTERS[4][5] ), .B(n3204), .S(n58), .Z(n2009) );
  MUX2_X1 U2379 ( .A(\REGISTERS[4][4] ), .B(n3205), .S(n58), .Z(n2008) );
  MUX2_X1 U2380 ( .A(\REGISTERS[4][3] ), .B(n3206), .S(n58), .Z(n2007) );
  MUX2_X1 U2381 ( .A(\REGISTERS[4][2] ), .B(n3207), .S(n58), .Z(n2006) );
  MUX2_X1 U2382 ( .A(\REGISTERS[4][1] ), .B(n3208), .S(n58), .Z(n2005) );
  MUX2_X1 U2383 ( .A(\REGISTERS[4][0] ), .B(n3209), .S(n58), .Z(n2004) );
  OAI21_X1 U2384 ( .B1(n3210), .B2(n3220), .A(n3212), .ZN(n3219) );
  MUX2_X1 U2385 ( .A(\REGISTERS[5][31] ), .B(n3177), .S(n52), .Z(n2003) );
  MUX2_X1 U2386 ( .A(\REGISTERS[5][30] ), .B(n3179), .S(n52), .Z(n2002) );
  MUX2_X1 U2387 ( .A(\REGISTERS[5][29] ), .B(n3180), .S(n52), .Z(n2001) );
  MUX2_X1 U2388 ( .A(\REGISTERS[5][28] ), .B(n3181), .S(n52), .Z(n2000) );
  MUX2_X1 U2389 ( .A(\REGISTERS[5][27] ), .B(n3182), .S(n52), .Z(n1999) );
  MUX2_X1 U2390 ( .A(\REGISTERS[5][26] ), .B(n3183), .S(n52), .Z(n1998) );
  MUX2_X1 U2391 ( .A(\REGISTERS[5][25] ), .B(n3184), .S(n52), .Z(n1997) );
  MUX2_X1 U2392 ( .A(\REGISTERS[5][24] ), .B(n3185), .S(n52), .Z(n1996) );
  MUX2_X1 U2393 ( .A(\REGISTERS[5][23] ), .B(n3186), .S(n52), .Z(n1995) );
  MUX2_X1 U2394 ( .A(\REGISTERS[5][22] ), .B(n3187), .S(n52), .Z(n1994) );
  MUX2_X1 U2395 ( .A(\REGISTERS[5][21] ), .B(n3188), .S(n52), .Z(n1993) );
  MUX2_X1 U2396 ( .A(\REGISTERS[5][20] ), .B(n3189), .S(n52), .Z(n1992) );
  MUX2_X1 U2397 ( .A(\REGISTERS[5][19] ), .B(n3190), .S(n52), .Z(n1991) );
  MUX2_X1 U2398 ( .A(\REGISTERS[5][18] ), .B(n3191), .S(n52), .Z(n1990) );
  MUX2_X1 U2399 ( .A(\REGISTERS[5][17] ), .B(n3192), .S(n52), .Z(n1989) );
  MUX2_X1 U2400 ( .A(\REGISTERS[5][16] ), .B(n3193), .S(n52), .Z(n1988) );
  MUX2_X1 U2401 ( .A(\REGISTERS[5][15] ), .B(n3194), .S(n52), .Z(n1987) );
  MUX2_X1 U2402 ( .A(\REGISTERS[5][14] ), .B(n3195), .S(n52), .Z(n1986) );
  MUX2_X1 U2403 ( .A(\REGISTERS[5][13] ), .B(n3196), .S(n52), .Z(n1985) );
  MUX2_X1 U2404 ( .A(\REGISTERS[5][12] ), .B(n3197), .S(n52), .Z(n1984) );
  MUX2_X1 U2405 ( .A(\REGISTERS[5][11] ), .B(n3198), .S(n52), .Z(n1983) );
  MUX2_X1 U2406 ( .A(\REGISTERS[5][10] ), .B(n3199), .S(n52), .Z(n1982) );
  MUX2_X1 U2407 ( .A(\REGISTERS[5][9] ), .B(n3200), .S(n52), .Z(n1981) );
  MUX2_X1 U2408 ( .A(\REGISTERS[5][8] ), .B(n3201), .S(n52), .Z(n1980) );
  MUX2_X1 U2409 ( .A(\REGISTERS[5][7] ), .B(n3202), .S(n52), .Z(n1979) );
  MUX2_X1 U2410 ( .A(\REGISTERS[5][6] ), .B(n3203), .S(n52), .Z(n1978) );
  MUX2_X1 U2411 ( .A(\REGISTERS[5][5] ), .B(n3204), .S(n52), .Z(n1977) );
  MUX2_X1 U2412 ( .A(\REGISTERS[5][4] ), .B(n3205), .S(n52), .Z(n1976) );
  MUX2_X1 U2413 ( .A(\REGISTERS[5][3] ), .B(n3206), .S(n52), .Z(n1975) );
  MUX2_X1 U2414 ( .A(\REGISTERS[5][2] ), .B(n3207), .S(n52), .Z(n1974) );
  MUX2_X1 U2415 ( .A(\REGISTERS[5][1] ), .B(n3208), .S(n52), .Z(n1973) );
  MUX2_X1 U2416 ( .A(\REGISTERS[5][0] ), .B(n3209), .S(n52), .Z(n1972) );
  OAI21_X1 U2417 ( .B1(n3210), .B2(n3222), .A(n3212), .ZN(n3221) );
  MUX2_X1 U2418 ( .A(\REGISTERS[6][31] ), .B(n3177), .S(n54), .Z(n1971) );
  MUX2_X1 U2419 ( .A(\REGISTERS[6][30] ), .B(n3179), .S(n54), .Z(n1970) );
  MUX2_X1 U2420 ( .A(\REGISTERS[6][29] ), .B(n3180), .S(n54), .Z(n1969) );
  MUX2_X1 U2421 ( .A(\REGISTERS[6][28] ), .B(n3181), .S(n54), .Z(n1968) );
  MUX2_X1 U2422 ( .A(\REGISTERS[6][27] ), .B(n3182), .S(n54), .Z(n1967) );
  MUX2_X1 U2423 ( .A(\REGISTERS[6][26] ), .B(n3183), .S(n54), .Z(n1966) );
  MUX2_X1 U2424 ( .A(\REGISTERS[6][25] ), .B(n3184), .S(n54), .Z(n1965) );
  MUX2_X1 U2425 ( .A(\REGISTERS[6][24] ), .B(n3185), .S(n54), .Z(n1964) );
  MUX2_X1 U2426 ( .A(\REGISTERS[6][23] ), .B(n3186), .S(n54), .Z(n1963) );
  MUX2_X1 U2427 ( .A(\REGISTERS[6][22] ), .B(n3187), .S(n54), .Z(n1962) );
  MUX2_X1 U2428 ( .A(\REGISTERS[6][21] ), .B(n3188), .S(n54), .Z(n1961) );
  MUX2_X1 U2429 ( .A(\REGISTERS[6][20] ), .B(n3189), .S(n54), .Z(n1960) );
  MUX2_X1 U2430 ( .A(\REGISTERS[6][19] ), .B(n3190), .S(n54), .Z(n1959) );
  MUX2_X1 U2431 ( .A(\REGISTERS[6][18] ), .B(n3191), .S(n54), .Z(n1958) );
  MUX2_X1 U2432 ( .A(\REGISTERS[6][17] ), .B(n3192), .S(n54), .Z(n1957) );
  MUX2_X1 U2433 ( .A(\REGISTERS[6][16] ), .B(n3193), .S(n54), .Z(n1956) );
  MUX2_X1 U2434 ( .A(\REGISTERS[6][15] ), .B(n3194), .S(n54), .Z(n1955) );
  MUX2_X1 U2435 ( .A(\REGISTERS[6][14] ), .B(n3195), .S(n54), .Z(n1954) );
  MUX2_X1 U2436 ( .A(\REGISTERS[6][13] ), .B(n3196), .S(n54), .Z(n1953) );
  MUX2_X1 U2437 ( .A(\REGISTERS[6][12] ), .B(n3197), .S(n54), .Z(n1952) );
  MUX2_X1 U2438 ( .A(\REGISTERS[6][11] ), .B(n3198), .S(n54), .Z(n1951) );
  MUX2_X1 U2439 ( .A(\REGISTERS[6][10] ), .B(n3199), .S(n54), .Z(n1950) );
  MUX2_X1 U2440 ( .A(\REGISTERS[6][9] ), .B(n3200), .S(n54), .Z(n1949) );
  MUX2_X1 U2441 ( .A(\REGISTERS[6][8] ), .B(n3201), .S(n54), .Z(n1948) );
  MUX2_X1 U2442 ( .A(\REGISTERS[6][7] ), .B(n3202), .S(n54), .Z(n1947) );
  MUX2_X1 U2443 ( .A(\REGISTERS[6][6] ), .B(n3203), .S(n54), .Z(n1946) );
  MUX2_X1 U2444 ( .A(\REGISTERS[6][5] ), .B(n3204), .S(n54), .Z(n1945) );
  MUX2_X1 U2445 ( .A(\REGISTERS[6][4] ), .B(n3205), .S(n54), .Z(n1944) );
  MUX2_X1 U2446 ( .A(\REGISTERS[6][3] ), .B(n3206), .S(n54), .Z(n1943) );
  MUX2_X1 U2447 ( .A(\REGISTERS[6][2] ), .B(n3207), .S(n54), .Z(n1942) );
  MUX2_X1 U2448 ( .A(\REGISTERS[6][1] ), .B(n3208), .S(n54), .Z(n1941) );
  MUX2_X1 U2449 ( .A(\REGISTERS[6][0] ), .B(n3209), .S(n54), .Z(n1940) );
  OAI21_X1 U2450 ( .B1(n3210), .B2(n3224), .A(n3212), .ZN(n3223) );
  MUX2_X1 U2451 ( .A(\REGISTERS[7][31] ), .B(n3177), .S(n48), .Z(n1939) );
  MUX2_X1 U2452 ( .A(\REGISTERS[7][30] ), .B(n3179), .S(n48), .Z(n1938) );
  MUX2_X1 U2453 ( .A(\REGISTERS[7][29] ), .B(n3180), .S(n48), .Z(n1937) );
  MUX2_X1 U2454 ( .A(\REGISTERS[7][28] ), .B(n3181), .S(n48), .Z(n1936) );
  MUX2_X1 U2455 ( .A(\REGISTERS[7][27] ), .B(n3182), .S(n48), .Z(n1935) );
  MUX2_X1 U2456 ( .A(\REGISTERS[7][26] ), .B(n3183), .S(n48), .Z(n1934) );
  MUX2_X1 U2457 ( .A(\REGISTERS[7][25] ), .B(n3184), .S(n48), .Z(n1933) );
  MUX2_X1 U2458 ( .A(\REGISTERS[7][24] ), .B(n3185), .S(n48), .Z(n1932) );
  MUX2_X1 U2459 ( .A(\REGISTERS[7][23] ), .B(n3186), .S(n48), .Z(n1931) );
  MUX2_X1 U2460 ( .A(\REGISTERS[7][22] ), .B(n3187), .S(n48), .Z(n1930) );
  MUX2_X1 U2461 ( .A(\REGISTERS[7][21] ), .B(n3188), .S(n48), .Z(n1929) );
  MUX2_X1 U2462 ( .A(\REGISTERS[7][20] ), .B(n3189), .S(n48), .Z(n1928) );
  MUX2_X1 U2463 ( .A(\REGISTERS[7][19] ), .B(n3190), .S(n48), .Z(n1927) );
  MUX2_X1 U2464 ( .A(\REGISTERS[7][18] ), .B(n3191), .S(n48), .Z(n1926) );
  MUX2_X1 U2465 ( .A(\REGISTERS[7][17] ), .B(n3192), .S(n48), .Z(n1925) );
  MUX2_X1 U2466 ( .A(\REGISTERS[7][16] ), .B(n3193), .S(n48), .Z(n1924) );
  MUX2_X1 U2467 ( .A(\REGISTERS[7][15] ), .B(n3194), .S(n48), .Z(n1923) );
  MUX2_X1 U2468 ( .A(\REGISTERS[7][14] ), .B(n3195), .S(n48), .Z(n1922) );
  MUX2_X1 U2469 ( .A(\REGISTERS[7][13] ), .B(n3196), .S(n48), .Z(n1921) );
  MUX2_X1 U2470 ( .A(\REGISTERS[7][12] ), .B(n3197), .S(n48), .Z(n1920) );
  MUX2_X1 U2471 ( .A(\REGISTERS[7][11] ), .B(n3198), .S(n48), .Z(n1919) );
  MUX2_X1 U2472 ( .A(\REGISTERS[7][10] ), .B(n3199), .S(n48), .Z(n1918) );
  MUX2_X1 U2473 ( .A(\REGISTERS[7][9] ), .B(n3200), .S(n48), .Z(n1917) );
  MUX2_X1 U2474 ( .A(\REGISTERS[7][8] ), .B(n3201), .S(n48), .Z(n1916) );
  MUX2_X1 U2475 ( .A(\REGISTERS[7][7] ), .B(n3202), .S(n48), .Z(n1915) );
  MUX2_X1 U2476 ( .A(\REGISTERS[7][6] ), .B(n3203), .S(n48), .Z(n1914) );
  MUX2_X1 U2477 ( .A(\REGISTERS[7][5] ), .B(n3204), .S(n48), .Z(n1913) );
  MUX2_X1 U2478 ( .A(\REGISTERS[7][4] ), .B(n3205), .S(n48), .Z(n1912) );
  MUX2_X1 U2479 ( .A(\REGISTERS[7][3] ), .B(n3206), .S(n48), .Z(n1911) );
  MUX2_X1 U2480 ( .A(\REGISTERS[7][2] ), .B(n3207), .S(n48), .Z(n1910) );
  MUX2_X1 U2481 ( .A(\REGISTERS[7][1] ), .B(n3208), .S(n48), .Z(n1909) );
  MUX2_X1 U2482 ( .A(\REGISTERS[7][0] ), .B(n3209), .S(n48), .Z(n1908) );
  OAI21_X1 U2483 ( .B1(n3210), .B2(n3226), .A(n3212), .ZN(n3225) );
  NAND3_X1 U2484 ( .A1(n3227), .A2(n3228), .A3(n3229), .ZN(n3210) );
  MUX2_X1 U2485 ( .A(\REGISTERS[8][31] ), .B(n3177), .S(n50), .Z(n1907) );
  MUX2_X1 U2486 ( .A(\REGISTERS[8][30] ), .B(n3179), .S(n50), .Z(n1906) );
  MUX2_X1 U2487 ( .A(\REGISTERS[8][29] ), .B(n3180), .S(n50), .Z(n1905) );
  MUX2_X1 U2488 ( .A(\REGISTERS[8][28] ), .B(n3181), .S(n50), .Z(n1904) );
  MUX2_X1 U2489 ( .A(\REGISTERS[8][27] ), .B(n3182), .S(n50), .Z(n1903) );
  MUX2_X1 U2490 ( .A(\REGISTERS[8][26] ), .B(n3183), .S(n50), .Z(n1902) );
  MUX2_X1 U2491 ( .A(\REGISTERS[8][25] ), .B(n3184), .S(n50), .Z(n1901) );
  MUX2_X1 U2492 ( .A(\REGISTERS[8][24] ), .B(n3185), .S(n50), .Z(n1900) );
  MUX2_X1 U2493 ( .A(\REGISTERS[8][23] ), .B(n3186), .S(n50), .Z(n1899) );
  MUX2_X1 U2494 ( .A(\REGISTERS[8][22] ), .B(n3187), .S(n50), .Z(n1898) );
  MUX2_X1 U2495 ( .A(\REGISTERS[8][21] ), .B(n3188), .S(n50), .Z(n1897) );
  MUX2_X1 U2496 ( .A(\REGISTERS[8][20] ), .B(n3189), .S(n50), .Z(n1896) );
  MUX2_X1 U2497 ( .A(\REGISTERS[8][19] ), .B(n3190), .S(n50), .Z(n1895) );
  MUX2_X1 U2498 ( .A(\REGISTERS[8][18] ), .B(n3191), .S(n50), .Z(n1894) );
  MUX2_X1 U2499 ( .A(\REGISTERS[8][17] ), .B(n3192), .S(n50), .Z(n1893) );
  MUX2_X1 U2500 ( .A(\REGISTERS[8][16] ), .B(n3193), .S(n50), .Z(n1892) );
  MUX2_X1 U2501 ( .A(\REGISTERS[8][15] ), .B(n3194), .S(n50), .Z(n1891) );
  MUX2_X1 U2502 ( .A(\REGISTERS[8][14] ), .B(n3195), .S(n50), .Z(n1890) );
  MUX2_X1 U2503 ( .A(\REGISTERS[8][13] ), .B(n3196), .S(n50), .Z(n1889) );
  MUX2_X1 U2504 ( .A(\REGISTERS[8][12] ), .B(n3197), .S(n50), .Z(n1888) );
  MUX2_X1 U2505 ( .A(\REGISTERS[8][11] ), .B(n3198), .S(n50), .Z(n1887) );
  MUX2_X1 U2506 ( .A(\REGISTERS[8][10] ), .B(n3199), .S(n50), .Z(n1886) );
  MUX2_X1 U2507 ( .A(\REGISTERS[8][9] ), .B(n3200), .S(n50), .Z(n1885) );
  MUX2_X1 U2508 ( .A(\REGISTERS[8][8] ), .B(n3201), .S(n50), .Z(n1884) );
  MUX2_X1 U2509 ( .A(\REGISTERS[8][7] ), .B(n3202), .S(n50), .Z(n1883) );
  MUX2_X1 U2510 ( .A(\REGISTERS[8][6] ), .B(n3203), .S(n50), .Z(n1882) );
  MUX2_X1 U2511 ( .A(\REGISTERS[8][5] ), .B(n3204), .S(n50), .Z(n1881) );
  MUX2_X1 U2512 ( .A(\REGISTERS[8][4] ), .B(n3205), .S(n50), .Z(n1880) );
  MUX2_X1 U2513 ( .A(\REGISTERS[8][3] ), .B(n3206), .S(n50), .Z(n1879) );
  MUX2_X1 U2514 ( .A(\REGISTERS[8][2] ), .B(n3207), .S(n50), .Z(n1878) );
  MUX2_X1 U2515 ( .A(\REGISTERS[8][1] ), .B(n3208), .S(n50), .Z(n1877) );
  MUX2_X1 U2516 ( .A(\REGISTERS[8][0] ), .B(n3209), .S(n50), .Z(n1876) );
  OAI21_X1 U2517 ( .B1(n3211), .B2(n3231), .A(n3212), .ZN(n3230) );
  MUX2_X1 U2518 ( .A(\REGISTERS[9][31] ), .B(n3177), .S(n44), .Z(n1875) );
  MUX2_X1 U2519 ( .A(\REGISTERS[9][30] ), .B(n3179), .S(n44), .Z(n1874) );
  MUX2_X1 U2520 ( .A(\REGISTERS[9][29] ), .B(n3180), .S(n44), .Z(n1873) );
  MUX2_X1 U2521 ( .A(\REGISTERS[9][28] ), .B(n3181), .S(n44), .Z(n1872) );
  MUX2_X1 U2522 ( .A(\REGISTERS[9][27] ), .B(n3182), .S(n44), .Z(n1871) );
  MUX2_X1 U2523 ( .A(\REGISTERS[9][26] ), .B(n3183), .S(n44), .Z(n1870) );
  MUX2_X1 U2524 ( .A(\REGISTERS[9][25] ), .B(n3184), .S(n44), .Z(n1869) );
  MUX2_X1 U2525 ( .A(\REGISTERS[9][24] ), .B(n3185), .S(n44), .Z(n1868) );
  MUX2_X1 U2526 ( .A(\REGISTERS[9][23] ), .B(n3186), .S(n44), .Z(n1867) );
  MUX2_X1 U2527 ( .A(\REGISTERS[9][22] ), .B(n3187), .S(n44), .Z(n1866) );
  MUX2_X1 U2528 ( .A(\REGISTERS[9][21] ), .B(n3188), .S(n44), .Z(n1865) );
  MUX2_X1 U2529 ( .A(\REGISTERS[9][20] ), .B(n3189), .S(n44), .Z(n1864) );
  MUX2_X1 U2530 ( .A(\REGISTERS[9][19] ), .B(n3190), .S(n44), .Z(n1863) );
  MUX2_X1 U2531 ( .A(\REGISTERS[9][18] ), .B(n3191), .S(n44), .Z(n1862) );
  MUX2_X1 U2532 ( .A(\REGISTERS[9][17] ), .B(n3192), .S(n44), .Z(n1861) );
  MUX2_X1 U2533 ( .A(\REGISTERS[9][16] ), .B(n3193), .S(n44), .Z(n1860) );
  MUX2_X1 U2534 ( .A(\REGISTERS[9][15] ), .B(n3194), .S(n44), .Z(n1859) );
  MUX2_X1 U2535 ( .A(\REGISTERS[9][14] ), .B(n3195), .S(n44), .Z(n1858) );
  MUX2_X1 U2536 ( .A(\REGISTERS[9][13] ), .B(n3196), .S(n44), .Z(n1857) );
  MUX2_X1 U2537 ( .A(\REGISTERS[9][12] ), .B(n3197), .S(n44), .Z(n1856) );
  MUX2_X1 U2538 ( .A(\REGISTERS[9][11] ), .B(n3198), .S(n44), .Z(n1855) );
  MUX2_X1 U2539 ( .A(\REGISTERS[9][10] ), .B(n3199), .S(n44), .Z(n1854) );
  MUX2_X1 U2540 ( .A(\REGISTERS[9][9] ), .B(n3200), .S(n44), .Z(n1853) );
  MUX2_X1 U2541 ( .A(\REGISTERS[9][8] ), .B(n3201), .S(n44), .Z(n1852) );
  MUX2_X1 U2542 ( .A(\REGISTERS[9][7] ), .B(n3202), .S(n44), .Z(n1851) );
  MUX2_X1 U2543 ( .A(\REGISTERS[9][6] ), .B(n3203), .S(n44), .Z(n1850) );
  MUX2_X1 U2544 ( .A(\REGISTERS[9][5] ), .B(n3204), .S(n44), .Z(n1849) );
  MUX2_X1 U2545 ( .A(\REGISTERS[9][4] ), .B(n3205), .S(n44), .Z(n1848) );
  MUX2_X1 U2546 ( .A(\REGISTERS[9][3] ), .B(n3206), .S(n44), .Z(n1847) );
  MUX2_X1 U2547 ( .A(\REGISTERS[9][2] ), .B(n3207), .S(n44), .Z(n1846) );
  MUX2_X1 U2548 ( .A(\REGISTERS[9][1] ), .B(n3208), .S(n44), .Z(n1845) );
  MUX2_X1 U2549 ( .A(\REGISTERS[9][0] ), .B(n3209), .S(n44), .Z(n1844) );
  OAI21_X1 U2550 ( .B1(n3214), .B2(n3231), .A(n3212), .ZN(n3232) );
  MUX2_X1 U2551 ( .A(\REGISTERS[10][31] ), .B(n3177), .S(n46), .Z(n1843) );
  MUX2_X1 U2552 ( .A(\REGISTERS[10][30] ), .B(n3179), .S(n46), .Z(n1842) );
  MUX2_X1 U2553 ( .A(\REGISTERS[10][29] ), .B(n3180), .S(n46), .Z(n1841) );
  MUX2_X1 U2554 ( .A(\REGISTERS[10][28] ), .B(n3181), .S(n46), .Z(n1840) );
  MUX2_X1 U2555 ( .A(\REGISTERS[10][27] ), .B(n3182), .S(n46), .Z(n1839) );
  MUX2_X1 U2556 ( .A(\REGISTERS[10][26] ), .B(n3183), .S(n46), .Z(n1838) );
  MUX2_X1 U2557 ( .A(\REGISTERS[10][25] ), .B(n3184), .S(n46), .Z(n1837) );
  MUX2_X1 U2558 ( .A(\REGISTERS[10][24] ), .B(n3185), .S(n46), .Z(n1836) );
  MUX2_X1 U2559 ( .A(\REGISTERS[10][23] ), .B(n3186), .S(n46), .Z(n1835) );
  MUX2_X1 U2560 ( .A(\REGISTERS[10][22] ), .B(n3187), .S(n46), .Z(n1834) );
  MUX2_X1 U2561 ( .A(\REGISTERS[10][21] ), .B(n3188), .S(n46), .Z(n1833) );
  MUX2_X1 U2562 ( .A(\REGISTERS[10][20] ), .B(n3189), .S(n46), .Z(n1832) );
  MUX2_X1 U2563 ( .A(\REGISTERS[10][19] ), .B(n3190), .S(n46), .Z(n1831) );
  MUX2_X1 U2564 ( .A(\REGISTERS[10][18] ), .B(n3191), .S(n46), .Z(n1830) );
  MUX2_X1 U2565 ( .A(\REGISTERS[10][17] ), .B(n3192), .S(n46), .Z(n1829) );
  MUX2_X1 U2566 ( .A(\REGISTERS[10][16] ), .B(n3193), .S(n46), .Z(n1828) );
  MUX2_X1 U2567 ( .A(\REGISTERS[10][15] ), .B(n3194), .S(n46), .Z(n1827) );
  MUX2_X1 U2568 ( .A(\REGISTERS[10][14] ), .B(n3195), .S(n46), .Z(n1826) );
  MUX2_X1 U2569 ( .A(\REGISTERS[10][13] ), .B(n3196), .S(n46), .Z(n1825) );
  MUX2_X1 U2570 ( .A(\REGISTERS[10][12] ), .B(n3197), .S(n46), .Z(n1824) );
  MUX2_X1 U2571 ( .A(\REGISTERS[10][11] ), .B(n3198), .S(n46), .Z(n1823) );
  MUX2_X1 U2572 ( .A(\REGISTERS[10][10] ), .B(n3199), .S(n46), .Z(n1822) );
  MUX2_X1 U2573 ( .A(\REGISTERS[10][9] ), .B(n3200), .S(n46), .Z(n1821) );
  MUX2_X1 U2574 ( .A(\REGISTERS[10][8] ), .B(n3201), .S(n46), .Z(n1820) );
  MUX2_X1 U2575 ( .A(\REGISTERS[10][7] ), .B(n3202), .S(n46), .Z(n1819) );
  MUX2_X1 U2576 ( .A(\REGISTERS[10][6] ), .B(n3203), .S(n46), .Z(n1818) );
  MUX2_X1 U2577 ( .A(\REGISTERS[10][5] ), .B(n3204), .S(n46), .Z(n1817) );
  MUX2_X1 U2578 ( .A(\REGISTERS[10][4] ), .B(n3205), .S(n46), .Z(n1816) );
  MUX2_X1 U2579 ( .A(\REGISTERS[10][3] ), .B(n3206), .S(n46), .Z(n1815) );
  MUX2_X1 U2580 ( .A(\REGISTERS[10][2] ), .B(n3207), .S(n46), .Z(n1814) );
  MUX2_X1 U2581 ( .A(\REGISTERS[10][1] ), .B(n3208), .S(n46), .Z(n1813) );
  MUX2_X1 U2582 ( .A(\REGISTERS[10][0] ), .B(n3209), .S(n46), .Z(n1812) );
  OAI21_X1 U2583 ( .B1(n3216), .B2(n3231), .A(n3212), .ZN(n3233) );
  MUX2_X1 U2584 ( .A(\REGISTERS[11][31] ), .B(n3177), .S(n40), .Z(n1811) );
  MUX2_X1 U2585 ( .A(\REGISTERS[11][30] ), .B(n3179), .S(n40), .Z(n1810) );
  MUX2_X1 U2586 ( .A(\REGISTERS[11][29] ), .B(n3180), .S(n40), .Z(n1809) );
  MUX2_X1 U2587 ( .A(\REGISTERS[11][28] ), .B(n3181), .S(n40), .Z(n1808) );
  MUX2_X1 U2588 ( .A(\REGISTERS[11][27] ), .B(n3182), .S(n40), .Z(n1807) );
  MUX2_X1 U2589 ( .A(\REGISTERS[11][26] ), .B(n3183), .S(n40), .Z(n1806) );
  MUX2_X1 U2590 ( .A(\REGISTERS[11][25] ), .B(n3184), .S(n40), .Z(n1805) );
  MUX2_X1 U2591 ( .A(\REGISTERS[11][24] ), .B(n3185), .S(n40), .Z(n1804) );
  MUX2_X1 U2592 ( .A(\REGISTERS[11][23] ), .B(n3186), .S(n40), .Z(n1803) );
  MUX2_X1 U2593 ( .A(\REGISTERS[11][22] ), .B(n3187), .S(n40), .Z(n1802) );
  MUX2_X1 U2594 ( .A(\REGISTERS[11][21] ), .B(n3188), .S(n40), .Z(n1801) );
  MUX2_X1 U2595 ( .A(\REGISTERS[11][20] ), .B(n3189), .S(n40), .Z(n1800) );
  MUX2_X1 U2596 ( .A(\REGISTERS[11][19] ), .B(n3190), .S(n40), .Z(n1799) );
  MUX2_X1 U2597 ( .A(\REGISTERS[11][18] ), .B(n3191), .S(n40), .Z(n1798) );
  MUX2_X1 U2598 ( .A(\REGISTERS[11][17] ), .B(n3192), .S(n40), .Z(n1797) );
  MUX2_X1 U2599 ( .A(\REGISTERS[11][16] ), .B(n3193), .S(n40), .Z(n1796) );
  MUX2_X1 U2600 ( .A(\REGISTERS[11][15] ), .B(n3194), .S(n40), .Z(n1795) );
  MUX2_X1 U2601 ( .A(\REGISTERS[11][14] ), .B(n3195), .S(n40), .Z(n1794) );
  MUX2_X1 U2602 ( .A(\REGISTERS[11][13] ), .B(n3196), .S(n40), .Z(n1793) );
  MUX2_X1 U2603 ( .A(\REGISTERS[11][12] ), .B(n3197), .S(n40), .Z(n1792) );
  MUX2_X1 U2604 ( .A(\REGISTERS[11][11] ), .B(n3198), .S(n40), .Z(n1791) );
  MUX2_X1 U2605 ( .A(\REGISTERS[11][10] ), .B(n3199), .S(n40), .Z(n1790) );
  MUX2_X1 U2606 ( .A(\REGISTERS[11][9] ), .B(n3200), .S(n40), .Z(n1789) );
  MUX2_X1 U2607 ( .A(\REGISTERS[11][8] ), .B(n3201), .S(n40), .Z(n1788) );
  MUX2_X1 U2608 ( .A(\REGISTERS[11][7] ), .B(n3202), .S(n40), .Z(n1787) );
  MUX2_X1 U2609 ( .A(\REGISTERS[11][6] ), .B(n3203), .S(n40), .Z(n1786) );
  MUX2_X1 U2610 ( .A(\REGISTERS[11][5] ), .B(n3204), .S(n40), .Z(n1785) );
  MUX2_X1 U2611 ( .A(\REGISTERS[11][4] ), .B(n3205), .S(n40), .Z(n1784) );
  MUX2_X1 U2612 ( .A(\REGISTERS[11][3] ), .B(n3206), .S(n40), .Z(n1783) );
  MUX2_X1 U2613 ( .A(\REGISTERS[11][2] ), .B(n3207), .S(n40), .Z(n1782) );
  MUX2_X1 U2614 ( .A(\REGISTERS[11][1] ), .B(n3208), .S(n40), .Z(n1781) );
  MUX2_X1 U2615 ( .A(\REGISTERS[11][0] ), .B(n3209), .S(n40), .Z(n1780) );
  OAI21_X1 U2616 ( .B1(n3218), .B2(n3231), .A(n3212), .ZN(n3234) );
  MUX2_X1 U2617 ( .A(\REGISTERS[12][31] ), .B(n3177), .S(n42), .Z(n1779) );
  MUX2_X1 U2618 ( .A(\REGISTERS[12][30] ), .B(n3179), .S(n42), .Z(n1778) );
  MUX2_X1 U2619 ( .A(\REGISTERS[12][29] ), .B(n3180), .S(n42), .Z(n1777) );
  MUX2_X1 U2620 ( .A(\REGISTERS[12][28] ), .B(n3181), .S(n42), .Z(n1776) );
  MUX2_X1 U2621 ( .A(\REGISTERS[12][27] ), .B(n3182), .S(n42), .Z(n1775) );
  MUX2_X1 U2622 ( .A(\REGISTERS[12][26] ), .B(n3183), .S(n42), .Z(n1774) );
  MUX2_X1 U2623 ( .A(\REGISTERS[12][25] ), .B(n3184), .S(n42), .Z(n1773) );
  MUX2_X1 U2624 ( .A(\REGISTERS[12][24] ), .B(n3185), .S(n42), .Z(n1772) );
  MUX2_X1 U2625 ( .A(\REGISTERS[12][23] ), .B(n3186), .S(n42), .Z(n1771) );
  MUX2_X1 U2626 ( .A(\REGISTERS[12][22] ), .B(n3187), .S(n42), .Z(n1770) );
  MUX2_X1 U2627 ( .A(\REGISTERS[12][21] ), .B(n3188), .S(n42), .Z(n1769) );
  MUX2_X1 U2628 ( .A(\REGISTERS[12][20] ), .B(n3189), .S(n42), .Z(n1768) );
  MUX2_X1 U2629 ( .A(\REGISTERS[12][19] ), .B(n3190), .S(n42), .Z(n1767) );
  MUX2_X1 U2630 ( .A(\REGISTERS[12][18] ), .B(n3191), .S(n42), .Z(n1766) );
  MUX2_X1 U2631 ( .A(\REGISTERS[12][17] ), .B(n3192), .S(n42), .Z(n1765) );
  MUX2_X1 U2632 ( .A(\REGISTERS[12][16] ), .B(n3193), .S(n42), .Z(n1764) );
  MUX2_X1 U2633 ( .A(\REGISTERS[12][15] ), .B(n3194), .S(n42), .Z(n1763) );
  MUX2_X1 U2634 ( .A(\REGISTERS[12][14] ), .B(n3195), .S(n42), .Z(n1762) );
  MUX2_X1 U2635 ( .A(\REGISTERS[12][13] ), .B(n3196), .S(n42), .Z(n1761) );
  MUX2_X1 U2636 ( .A(\REGISTERS[12][12] ), .B(n3197), .S(n42), .Z(n1760) );
  MUX2_X1 U2637 ( .A(\REGISTERS[12][11] ), .B(n3198), .S(n42), .Z(n1759) );
  MUX2_X1 U2638 ( .A(\REGISTERS[12][10] ), .B(n3199), .S(n42), .Z(n1758) );
  MUX2_X1 U2639 ( .A(\REGISTERS[12][9] ), .B(n3200), .S(n42), .Z(n1757) );
  MUX2_X1 U2640 ( .A(\REGISTERS[12][8] ), .B(n3201), .S(n42), .Z(n1756) );
  MUX2_X1 U2641 ( .A(\REGISTERS[12][7] ), .B(n3202), .S(n42), .Z(n1755) );
  MUX2_X1 U2642 ( .A(\REGISTERS[12][6] ), .B(n3203), .S(n42), .Z(n1754) );
  MUX2_X1 U2643 ( .A(\REGISTERS[12][5] ), .B(n3204), .S(n42), .Z(n1753) );
  MUX2_X1 U2644 ( .A(\REGISTERS[12][4] ), .B(n3205), .S(n42), .Z(n1752) );
  MUX2_X1 U2645 ( .A(\REGISTERS[12][3] ), .B(n3206), .S(n42), .Z(n1751) );
  MUX2_X1 U2646 ( .A(\REGISTERS[12][2] ), .B(n3207), .S(n42), .Z(n1750) );
  MUX2_X1 U2647 ( .A(\REGISTERS[12][1] ), .B(n3208), .S(n42), .Z(n1749) );
  MUX2_X1 U2648 ( .A(\REGISTERS[12][0] ), .B(n3209), .S(n42), .Z(n1748) );
  OAI21_X1 U2649 ( .B1(n3220), .B2(n3231), .A(n3212), .ZN(n3235) );
  MUX2_X1 U2650 ( .A(\REGISTERS[13][31] ), .B(n3177), .S(n36), .Z(n1747) );
  MUX2_X1 U2651 ( .A(\REGISTERS[13][30] ), .B(n3179), .S(n36), .Z(n1746) );
  MUX2_X1 U2652 ( .A(\REGISTERS[13][29] ), .B(n3180), .S(n36), .Z(n1745) );
  MUX2_X1 U2653 ( .A(\REGISTERS[13][28] ), .B(n3181), .S(n36), .Z(n1744) );
  MUX2_X1 U2654 ( .A(\REGISTERS[13][27] ), .B(n3182), .S(n36), .Z(n1743) );
  MUX2_X1 U2655 ( .A(\REGISTERS[13][26] ), .B(n3183), .S(n36), .Z(n1742) );
  MUX2_X1 U2656 ( .A(\REGISTERS[13][25] ), .B(n3184), .S(n36), .Z(n1741) );
  MUX2_X1 U2657 ( .A(\REGISTERS[13][24] ), .B(n3185), .S(n36), .Z(n1740) );
  MUX2_X1 U2658 ( .A(\REGISTERS[13][23] ), .B(n3186), .S(n36), .Z(n1739) );
  MUX2_X1 U2659 ( .A(\REGISTERS[13][22] ), .B(n3187), .S(n36), .Z(n1738) );
  MUX2_X1 U2660 ( .A(\REGISTERS[13][21] ), .B(n3188), .S(n36), .Z(n1737) );
  MUX2_X1 U2661 ( .A(\REGISTERS[13][20] ), .B(n3189), .S(n36), .Z(n1736) );
  MUX2_X1 U2662 ( .A(\REGISTERS[13][19] ), .B(n3190), .S(n36), .Z(n1735) );
  MUX2_X1 U2663 ( .A(\REGISTERS[13][18] ), .B(n3191), .S(n36), .Z(n1734) );
  MUX2_X1 U2664 ( .A(\REGISTERS[13][17] ), .B(n3192), .S(n36), .Z(n1733) );
  MUX2_X1 U2665 ( .A(\REGISTERS[13][16] ), .B(n3193), .S(n36), .Z(n1732) );
  MUX2_X1 U2666 ( .A(\REGISTERS[13][15] ), .B(n3194), .S(n36), .Z(n1731) );
  MUX2_X1 U2667 ( .A(\REGISTERS[13][14] ), .B(n3195), .S(n36), .Z(n1730) );
  MUX2_X1 U2668 ( .A(\REGISTERS[13][13] ), .B(n3196), .S(n36), .Z(n1729) );
  MUX2_X1 U2669 ( .A(\REGISTERS[13][12] ), .B(n3197), .S(n36), .Z(n1728) );
  MUX2_X1 U2670 ( .A(\REGISTERS[13][11] ), .B(n3198), .S(n36), .Z(n1727) );
  MUX2_X1 U2671 ( .A(\REGISTERS[13][10] ), .B(n3199), .S(n36), .Z(n1726) );
  MUX2_X1 U2672 ( .A(\REGISTERS[13][9] ), .B(n3200), .S(n36), .Z(n1725) );
  MUX2_X1 U2673 ( .A(\REGISTERS[13][8] ), .B(n3201), .S(n36), .Z(n1724) );
  MUX2_X1 U2674 ( .A(\REGISTERS[13][7] ), .B(n3202), .S(n36), .Z(n1723) );
  MUX2_X1 U2675 ( .A(\REGISTERS[13][6] ), .B(n3203), .S(n36), .Z(n1722) );
  MUX2_X1 U2676 ( .A(\REGISTERS[13][5] ), .B(n3204), .S(n36), .Z(n1721) );
  MUX2_X1 U2677 ( .A(\REGISTERS[13][4] ), .B(n3205), .S(n36), .Z(n1720) );
  MUX2_X1 U2678 ( .A(\REGISTERS[13][3] ), .B(n3206), .S(n36), .Z(n1719) );
  MUX2_X1 U2679 ( .A(\REGISTERS[13][2] ), .B(n3207), .S(n36), .Z(n1718) );
  MUX2_X1 U2680 ( .A(\REGISTERS[13][1] ), .B(n3208), .S(n36), .Z(n1717) );
  MUX2_X1 U2681 ( .A(\REGISTERS[13][0] ), .B(n3209), .S(n36), .Z(n1716) );
  OAI21_X1 U2682 ( .B1(n3222), .B2(n3231), .A(n3212), .ZN(n3236) );
  MUX2_X1 U2683 ( .A(\REGISTERS[14][31] ), .B(n3177), .S(n38), .Z(n1715) );
  MUX2_X1 U2684 ( .A(\REGISTERS[14][30] ), .B(n3179), .S(n38), .Z(n1714) );
  MUX2_X1 U2685 ( .A(\REGISTERS[14][29] ), .B(n3180), .S(n38), .Z(n1713) );
  MUX2_X1 U2686 ( .A(\REGISTERS[14][28] ), .B(n3181), .S(n38), .Z(n1712) );
  MUX2_X1 U2687 ( .A(\REGISTERS[14][27] ), .B(n3182), .S(n38), .Z(n1711) );
  MUX2_X1 U2688 ( .A(\REGISTERS[14][26] ), .B(n3183), .S(n38), .Z(n1710) );
  MUX2_X1 U2689 ( .A(\REGISTERS[14][25] ), .B(n3184), .S(n38), .Z(n1709) );
  MUX2_X1 U2690 ( .A(\REGISTERS[14][24] ), .B(n3185), .S(n38), .Z(n1708) );
  MUX2_X1 U2691 ( .A(\REGISTERS[14][23] ), .B(n3186), .S(n38), .Z(n1707) );
  MUX2_X1 U2692 ( .A(\REGISTERS[14][22] ), .B(n3187), .S(n38), .Z(n1706) );
  MUX2_X1 U2693 ( .A(\REGISTERS[14][21] ), .B(n3188), .S(n38), .Z(n1705) );
  MUX2_X1 U2694 ( .A(\REGISTERS[14][20] ), .B(n3189), .S(n38), .Z(n1704) );
  MUX2_X1 U2695 ( .A(\REGISTERS[14][19] ), .B(n3190), .S(n38), .Z(n1703) );
  MUX2_X1 U2696 ( .A(\REGISTERS[14][18] ), .B(n3191), .S(n38), .Z(n1702) );
  MUX2_X1 U2697 ( .A(\REGISTERS[14][17] ), .B(n3192), .S(n38), .Z(n1701) );
  MUX2_X1 U2698 ( .A(\REGISTERS[14][16] ), .B(n3193), .S(n38), .Z(n1700) );
  MUX2_X1 U2699 ( .A(\REGISTERS[14][15] ), .B(n3194), .S(n38), .Z(n1699) );
  MUX2_X1 U2700 ( .A(\REGISTERS[14][14] ), .B(n3195), .S(n38), .Z(n1698) );
  MUX2_X1 U2701 ( .A(\REGISTERS[14][13] ), .B(n3196), .S(n38), .Z(n1697) );
  MUX2_X1 U2702 ( .A(\REGISTERS[14][12] ), .B(n3197), .S(n38), .Z(n1696) );
  MUX2_X1 U2703 ( .A(\REGISTERS[14][11] ), .B(n3198), .S(n38), .Z(n1695) );
  MUX2_X1 U2704 ( .A(\REGISTERS[14][10] ), .B(n3199), .S(n38), .Z(n1694) );
  MUX2_X1 U2705 ( .A(\REGISTERS[14][9] ), .B(n3200), .S(n38), .Z(n1693) );
  MUX2_X1 U2706 ( .A(\REGISTERS[14][8] ), .B(n3201), .S(n38), .Z(n1692) );
  MUX2_X1 U2707 ( .A(\REGISTERS[14][7] ), .B(n3202), .S(n38), .Z(n1691) );
  MUX2_X1 U2708 ( .A(\REGISTERS[14][6] ), .B(n3203), .S(n38), .Z(n1690) );
  MUX2_X1 U2709 ( .A(\REGISTERS[14][5] ), .B(n3204), .S(n38), .Z(n1689) );
  MUX2_X1 U2710 ( .A(\REGISTERS[14][4] ), .B(n3205), .S(n38), .Z(n1688) );
  MUX2_X1 U2711 ( .A(\REGISTERS[14][3] ), .B(n3206), .S(n38), .Z(n1687) );
  MUX2_X1 U2712 ( .A(\REGISTERS[14][2] ), .B(n3207), .S(n38), .Z(n1686) );
  MUX2_X1 U2713 ( .A(\REGISTERS[14][1] ), .B(n3208), .S(n38), .Z(n1685) );
  MUX2_X1 U2714 ( .A(\REGISTERS[14][0] ), .B(n3209), .S(n38), .Z(n1684) );
  OAI21_X1 U2715 ( .B1(n3224), .B2(n3231), .A(n3212), .ZN(n3237) );
  MUX2_X1 U2716 ( .A(\REGISTERS[15][31] ), .B(n3177), .S(n32), .Z(n1683) );
  MUX2_X1 U2717 ( .A(\REGISTERS[15][30] ), .B(n3179), .S(n32), .Z(n1682) );
  MUX2_X1 U2718 ( .A(\REGISTERS[15][29] ), .B(n3180), .S(n32), .Z(n1681) );
  MUX2_X1 U2719 ( .A(\REGISTERS[15][28] ), .B(n3181), .S(n32), .Z(n1680) );
  MUX2_X1 U2720 ( .A(\REGISTERS[15][27] ), .B(n3182), .S(n32), .Z(n1679) );
  MUX2_X1 U2721 ( .A(\REGISTERS[15][26] ), .B(n3183), .S(n32), .Z(n1678) );
  MUX2_X1 U2722 ( .A(\REGISTERS[15][25] ), .B(n3184), .S(n32), .Z(n1677) );
  MUX2_X1 U2723 ( .A(\REGISTERS[15][24] ), .B(n3185), .S(n32), .Z(n1676) );
  MUX2_X1 U2724 ( .A(\REGISTERS[15][23] ), .B(n3186), .S(n32), .Z(n1675) );
  MUX2_X1 U2725 ( .A(\REGISTERS[15][22] ), .B(n3187), .S(n32), .Z(n1674) );
  MUX2_X1 U2726 ( .A(\REGISTERS[15][21] ), .B(n3188), .S(n32), .Z(n1673) );
  MUX2_X1 U2727 ( .A(\REGISTERS[15][20] ), .B(n3189), .S(n32), .Z(n1672) );
  MUX2_X1 U2728 ( .A(\REGISTERS[15][19] ), .B(n3190), .S(n32), .Z(n1671) );
  MUX2_X1 U2729 ( .A(\REGISTERS[15][18] ), .B(n3191), .S(n32), .Z(n1670) );
  MUX2_X1 U2730 ( .A(\REGISTERS[15][17] ), .B(n3192), .S(n32), .Z(n1669) );
  MUX2_X1 U2731 ( .A(\REGISTERS[15][16] ), .B(n3193), .S(n32), .Z(n1668) );
  MUX2_X1 U2732 ( .A(\REGISTERS[15][15] ), .B(n3194), .S(n32), .Z(n1667) );
  MUX2_X1 U2733 ( .A(\REGISTERS[15][14] ), .B(n3195), .S(n32), .Z(n1666) );
  MUX2_X1 U2734 ( .A(\REGISTERS[15][13] ), .B(n3196), .S(n32), .Z(n1665) );
  MUX2_X1 U2735 ( .A(\REGISTERS[15][12] ), .B(n3197), .S(n32), .Z(n1664) );
  MUX2_X1 U2736 ( .A(\REGISTERS[15][11] ), .B(n3198), .S(n32), .Z(n1663) );
  MUX2_X1 U2737 ( .A(\REGISTERS[15][10] ), .B(n3199), .S(n32), .Z(n1662) );
  MUX2_X1 U2738 ( .A(\REGISTERS[15][9] ), .B(n3200), .S(n32), .Z(n1661) );
  MUX2_X1 U2739 ( .A(\REGISTERS[15][8] ), .B(n3201), .S(n32), .Z(n1660) );
  MUX2_X1 U2740 ( .A(\REGISTERS[15][7] ), .B(n3202), .S(n32), .Z(n1659) );
  MUX2_X1 U2741 ( .A(\REGISTERS[15][6] ), .B(n3203), .S(n32), .Z(n1658) );
  MUX2_X1 U2742 ( .A(\REGISTERS[15][5] ), .B(n3204), .S(n32), .Z(n1657) );
  MUX2_X1 U2743 ( .A(\REGISTERS[15][4] ), .B(n3205), .S(n32), .Z(n1656) );
  MUX2_X1 U2744 ( .A(\REGISTERS[15][3] ), .B(n3206), .S(n32), .Z(n1655) );
  MUX2_X1 U2745 ( .A(\REGISTERS[15][2] ), .B(n3207), .S(n32), .Z(n1654) );
  MUX2_X1 U2746 ( .A(\REGISTERS[15][1] ), .B(n3208), .S(n32), .Z(n1653) );
  MUX2_X1 U2747 ( .A(\REGISTERS[15][0] ), .B(n3209), .S(n32), .Z(n1652) );
  OAI21_X1 U2748 ( .B1(n3226), .B2(n3231), .A(n3212), .ZN(n3238) );
  NAND3_X1 U2749 ( .A1(n3229), .A2(n3228), .A3(ADD_WR[3]), .ZN(n3231) );
  INV_X1 U2750 ( .A(ADD_WR[4]), .ZN(n3228) );
  MUX2_X1 U2751 ( .A(\REGISTERS[16][31] ), .B(n3177), .S(n34), .Z(n1651) );
  MUX2_X1 U2752 ( .A(\REGISTERS[16][30] ), .B(n3179), .S(n34), .Z(n1650) );
  MUX2_X1 U2753 ( .A(\REGISTERS[16][29] ), .B(n3180), .S(n34), .Z(n1649) );
  MUX2_X1 U2754 ( .A(\REGISTERS[16][28] ), .B(n3181), .S(n34), .Z(n1648) );
  MUX2_X1 U2755 ( .A(\REGISTERS[16][27] ), .B(n3182), .S(n34), .Z(n1647) );
  MUX2_X1 U2756 ( .A(\REGISTERS[16][26] ), .B(n3183), .S(n34), .Z(n1646) );
  MUX2_X1 U2757 ( .A(\REGISTERS[16][25] ), .B(n3184), .S(n34), .Z(n1645) );
  MUX2_X1 U2758 ( .A(\REGISTERS[16][24] ), .B(n3185), .S(n34), .Z(n1644) );
  MUX2_X1 U2759 ( .A(\REGISTERS[16][23] ), .B(n3186), .S(n34), .Z(n1643) );
  MUX2_X1 U2760 ( .A(\REGISTERS[16][22] ), .B(n3187), .S(n34), .Z(n1642) );
  MUX2_X1 U2761 ( .A(\REGISTERS[16][21] ), .B(n3188), .S(n34), .Z(n1641) );
  MUX2_X1 U2762 ( .A(\REGISTERS[16][20] ), .B(n3189), .S(n34), .Z(n1640) );
  MUX2_X1 U2763 ( .A(\REGISTERS[16][19] ), .B(n3190), .S(n34), .Z(n1639) );
  MUX2_X1 U2764 ( .A(\REGISTERS[16][18] ), .B(n3191), .S(n34), .Z(n1638) );
  MUX2_X1 U2765 ( .A(\REGISTERS[16][17] ), .B(n3192), .S(n34), .Z(n1637) );
  MUX2_X1 U2766 ( .A(\REGISTERS[16][16] ), .B(n3193), .S(n34), .Z(n1636) );
  MUX2_X1 U2767 ( .A(\REGISTERS[16][15] ), .B(n3194), .S(n34), .Z(n1635) );
  MUX2_X1 U2768 ( .A(\REGISTERS[16][14] ), .B(n3195), .S(n34), .Z(n1634) );
  MUX2_X1 U2769 ( .A(\REGISTERS[16][13] ), .B(n3196), .S(n34), .Z(n1633) );
  MUX2_X1 U2770 ( .A(\REGISTERS[16][12] ), .B(n3197), .S(n34), .Z(n1632) );
  MUX2_X1 U2771 ( .A(\REGISTERS[16][11] ), .B(n3198), .S(n34), .Z(n1631) );
  MUX2_X1 U2772 ( .A(\REGISTERS[16][10] ), .B(n3199), .S(n34), .Z(n1630) );
  MUX2_X1 U2773 ( .A(\REGISTERS[16][9] ), .B(n3200), .S(n34), .Z(n1629) );
  MUX2_X1 U2774 ( .A(\REGISTERS[16][8] ), .B(n3201), .S(n34), .Z(n1628) );
  MUX2_X1 U2775 ( .A(\REGISTERS[16][7] ), .B(n3202), .S(n34), .Z(n1627) );
  MUX2_X1 U2776 ( .A(\REGISTERS[16][6] ), .B(n3203), .S(n34), .Z(n1626) );
  MUX2_X1 U2777 ( .A(\REGISTERS[16][5] ), .B(n3204), .S(n34), .Z(n1625) );
  MUX2_X1 U2778 ( .A(\REGISTERS[16][4] ), .B(n3205), .S(n34), .Z(n1624) );
  MUX2_X1 U2779 ( .A(\REGISTERS[16][3] ), .B(n3206), .S(n34), .Z(n1623) );
  MUX2_X1 U2780 ( .A(\REGISTERS[16][2] ), .B(n3207), .S(n34), .Z(n1622) );
  MUX2_X1 U2781 ( .A(\REGISTERS[16][1] ), .B(n3208), .S(n34), .Z(n1621) );
  MUX2_X1 U2782 ( .A(\REGISTERS[16][0] ), .B(n3209), .S(n34), .Z(n1620) );
  OAI21_X1 U2783 ( .B1(n3211), .B2(n3240), .A(n3212), .ZN(n3239) );
  MUX2_X1 U2784 ( .A(\REGISTERS[17][31] ), .B(n3177), .S(n28), .Z(n1619) );
  MUX2_X1 U2785 ( .A(\REGISTERS[17][30] ), .B(n3179), .S(n28), .Z(n1618) );
  MUX2_X1 U2786 ( .A(\REGISTERS[17][29] ), .B(n3180), .S(n28), .Z(n1617) );
  MUX2_X1 U2787 ( .A(\REGISTERS[17][28] ), .B(n3181), .S(n28), .Z(n1616) );
  MUX2_X1 U2788 ( .A(\REGISTERS[17][27] ), .B(n3182), .S(n28), .Z(n1615) );
  MUX2_X1 U2789 ( .A(\REGISTERS[17][26] ), .B(n3183), .S(n28), .Z(n1614) );
  MUX2_X1 U2790 ( .A(\REGISTERS[17][25] ), .B(n3184), .S(n28), .Z(n1613) );
  MUX2_X1 U2791 ( .A(\REGISTERS[17][24] ), .B(n3185), .S(n28), .Z(n1612) );
  MUX2_X1 U2792 ( .A(\REGISTERS[17][23] ), .B(n3186), .S(n28), .Z(n1611) );
  MUX2_X1 U2793 ( .A(\REGISTERS[17][22] ), .B(n3187), .S(n28), .Z(n1610) );
  MUX2_X1 U2794 ( .A(\REGISTERS[17][21] ), .B(n3188), .S(n28), .Z(n1609) );
  MUX2_X1 U2795 ( .A(\REGISTERS[17][20] ), .B(n3189), .S(n28), .Z(n1608) );
  MUX2_X1 U2796 ( .A(\REGISTERS[17][19] ), .B(n3190), .S(n28), .Z(n1607) );
  MUX2_X1 U2797 ( .A(\REGISTERS[17][18] ), .B(n3191), .S(n28), .Z(n1606) );
  MUX2_X1 U2798 ( .A(\REGISTERS[17][17] ), .B(n3192), .S(n28), .Z(n1605) );
  MUX2_X1 U2799 ( .A(\REGISTERS[17][16] ), .B(n3193), .S(n28), .Z(n1604) );
  MUX2_X1 U2800 ( .A(\REGISTERS[17][15] ), .B(n3194), .S(n28), .Z(n1603) );
  MUX2_X1 U2801 ( .A(\REGISTERS[17][14] ), .B(n3195), .S(n28), .Z(n1602) );
  MUX2_X1 U2802 ( .A(\REGISTERS[17][13] ), .B(n3196), .S(n28), .Z(n1601) );
  MUX2_X1 U2803 ( .A(\REGISTERS[17][12] ), .B(n3197), .S(n28), .Z(n1600) );
  MUX2_X1 U2804 ( .A(\REGISTERS[17][11] ), .B(n3198), .S(n28), .Z(n1599) );
  MUX2_X1 U2805 ( .A(\REGISTERS[17][10] ), .B(n3199), .S(n28), .Z(n1598) );
  MUX2_X1 U2806 ( .A(\REGISTERS[17][9] ), .B(n3200), .S(n28), .Z(n1597) );
  MUX2_X1 U2807 ( .A(\REGISTERS[17][8] ), .B(n3201), .S(n28), .Z(n1596) );
  MUX2_X1 U2808 ( .A(\REGISTERS[17][7] ), .B(n3202), .S(n28), .Z(n1595) );
  MUX2_X1 U2809 ( .A(\REGISTERS[17][6] ), .B(n3203), .S(n28), .Z(n1594) );
  MUX2_X1 U2810 ( .A(\REGISTERS[17][5] ), .B(n3204), .S(n28), .Z(n1593) );
  MUX2_X1 U2811 ( .A(\REGISTERS[17][4] ), .B(n3205), .S(n28), .Z(n1592) );
  MUX2_X1 U2812 ( .A(\REGISTERS[17][3] ), .B(n3206), .S(n28), .Z(n1591) );
  MUX2_X1 U2813 ( .A(\REGISTERS[17][2] ), .B(n3207), .S(n28), .Z(n1590) );
  MUX2_X1 U2814 ( .A(\REGISTERS[17][1] ), .B(n3208), .S(n28), .Z(n1589) );
  MUX2_X1 U2815 ( .A(\REGISTERS[17][0] ), .B(n3209), .S(n28), .Z(n1588) );
  OAI21_X1 U2816 ( .B1(n3214), .B2(n3240), .A(n3212), .ZN(n3241) );
  MUX2_X1 U2817 ( .A(\REGISTERS[18][31] ), .B(n3177), .S(n30), .Z(n1587) );
  MUX2_X1 U2818 ( .A(\REGISTERS[18][30] ), .B(n3179), .S(n30), .Z(n1586) );
  MUX2_X1 U2819 ( .A(\REGISTERS[18][29] ), .B(n3180), .S(n30), .Z(n1585) );
  MUX2_X1 U2820 ( .A(\REGISTERS[18][28] ), .B(n3181), .S(n30), .Z(n1584) );
  MUX2_X1 U2821 ( .A(\REGISTERS[18][27] ), .B(n3182), .S(n30), .Z(n1583) );
  MUX2_X1 U2822 ( .A(\REGISTERS[18][26] ), .B(n3183), .S(n30), .Z(n1582) );
  MUX2_X1 U2823 ( .A(\REGISTERS[18][25] ), .B(n3184), .S(n30), .Z(n1581) );
  MUX2_X1 U2824 ( .A(\REGISTERS[18][24] ), .B(n3185), .S(n30), .Z(n1580) );
  MUX2_X1 U2825 ( .A(\REGISTERS[18][23] ), .B(n3186), .S(n30), .Z(n1579) );
  MUX2_X1 U2826 ( .A(\REGISTERS[18][22] ), .B(n3187), .S(n30), .Z(n1578) );
  MUX2_X1 U2827 ( .A(\REGISTERS[18][21] ), .B(n3188), .S(n30), .Z(n1577) );
  MUX2_X1 U2828 ( .A(\REGISTERS[18][20] ), .B(n3189), .S(n30), .Z(n1576) );
  MUX2_X1 U2829 ( .A(\REGISTERS[18][19] ), .B(n3190), .S(n30), .Z(n1575) );
  MUX2_X1 U2830 ( .A(\REGISTERS[18][18] ), .B(n3191), .S(n30), .Z(n1574) );
  MUX2_X1 U2831 ( .A(\REGISTERS[18][17] ), .B(n3192), .S(n30), .Z(n1573) );
  MUX2_X1 U2832 ( .A(\REGISTERS[18][16] ), .B(n3193), .S(n30), .Z(n1572) );
  MUX2_X1 U2833 ( .A(\REGISTERS[18][15] ), .B(n3194), .S(n30), .Z(n1571) );
  MUX2_X1 U2834 ( .A(\REGISTERS[18][14] ), .B(n3195), .S(n30), .Z(n1570) );
  MUX2_X1 U2835 ( .A(\REGISTERS[18][13] ), .B(n3196), .S(n30), .Z(n1569) );
  MUX2_X1 U2836 ( .A(\REGISTERS[18][12] ), .B(n3197), .S(n30), .Z(n1568) );
  MUX2_X1 U2837 ( .A(\REGISTERS[18][11] ), .B(n3198), .S(n30), .Z(n1567) );
  MUX2_X1 U2838 ( .A(\REGISTERS[18][10] ), .B(n3199), .S(n30), .Z(n1566) );
  MUX2_X1 U2839 ( .A(\REGISTERS[18][9] ), .B(n3200), .S(n30), .Z(n1565) );
  MUX2_X1 U2840 ( .A(\REGISTERS[18][8] ), .B(n3201), .S(n30), .Z(n1564) );
  MUX2_X1 U2841 ( .A(\REGISTERS[18][7] ), .B(n3202), .S(n30), .Z(n1563) );
  MUX2_X1 U2842 ( .A(\REGISTERS[18][6] ), .B(n3203), .S(n30), .Z(n1562) );
  MUX2_X1 U2843 ( .A(\REGISTERS[18][5] ), .B(n3204), .S(n30), .Z(n1561) );
  MUX2_X1 U2844 ( .A(\REGISTERS[18][4] ), .B(n3205), .S(n30), .Z(n1560) );
  MUX2_X1 U2845 ( .A(\REGISTERS[18][3] ), .B(n3206), .S(n30), .Z(n1559) );
  MUX2_X1 U2846 ( .A(\REGISTERS[18][2] ), .B(n3207), .S(n30), .Z(n1558) );
  MUX2_X1 U2847 ( .A(\REGISTERS[18][1] ), .B(n3208), .S(n30), .Z(n1557) );
  MUX2_X1 U2848 ( .A(\REGISTERS[18][0] ), .B(n3209), .S(n30), .Z(n1556) );
  OAI21_X1 U2849 ( .B1(n3216), .B2(n3240), .A(n3212), .ZN(n3242) );
  MUX2_X1 U2850 ( .A(\REGISTERS[19][31] ), .B(n3177), .S(n2), .Z(n1555) );
  MUX2_X1 U2851 ( .A(\REGISTERS[19][30] ), .B(n3179), .S(n2), .Z(n1554) );
  MUX2_X1 U2852 ( .A(\REGISTERS[19][29] ), .B(n3180), .S(n2), .Z(n1553) );
  MUX2_X1 U2853 ( .A(\REGISTERS[19][28] ), .B(n3181), .S(n2), .Z(n1552) );
  MUX2_X1 U2854 ( .A(\REGISTERS[19][27] ), .B(n3182), .S(n2), .Z(n1551) );
  MUX2_X1 U2855 ( .A(\REGISTERS[19][26] ), .B(n3183), .S(n2), .Z(n1550) );
  MUX2_X1 U2856 ( .A(\REGISTERS[19][25] ), .B(n3184), .S(n2), .Z(n1549) );
  MUX2_X1 U2857 ( .A(\REGISTERS[19][24] ), .B(n3185), .S(n2), .Z(n1548) );
  MUX2_X1 U2858 ( .A(\REGISTERS[19][23] ), .B(n3186), .S(n2), .Z(n1547) );
  MUX2_X1 U2859 ( .A(\REGISTERS[19][22] ), .B(n3187), .S(n2), .Z(n1546) );
  MUX2_X1 U2860 ( .A(\REGISTERS[19][21] ), .B(n3188), .S(n2), .Z(n1545) );
  MUX2_X1 U2861 ( .A(\REGISTERS[19][20] ), .B(n3189), .S(n2), .Z(n1544) );
  MUX2_X1 U2862 ( .A(\REGISTERS[19][19] ), .B(n3190), .S(n2), .Z(n1543) );
  MUX2_X1 U2863 ( .A(\REGISTERS[19][18] ), .B(n3191), .S(n2), .Z(n1542) );
  MUX2_X1 U2864 ( .A(\REGISTERS[19][17] ), .B(n3192), .S(n2), .Z(n1541) );
  MUX2_X1 U2865 ( .A(\REGISTERS[19][16] ), .B(n3193), .S(n2), .Z(n1540) );
  MUX2_X1 U2866 ( .A(\REGISTERS[19][15] ), .B(n3194), .S(n2), .Z(n1539) );
  MUX2_X1 U2867 ( .A(\REGISTERS[19][14] ), .B(n3195), .S(n2), .Z(n1538) );
  MUX2_X1 U2868 ( .A(\REGISTERS[19][13] ), .B(n3196), .S(n2), .Z(n1537) );
  MUX2_X1 U2869 ( .A(\REGISTERS[19][12] ), .B(n3197), .S(n2), .Z(n1536) );
  MUX2_X1 U2870 ( .A(\REGISTERS[19][11] ), .B(n3198), .S(n2), .Z(n1535) );
  MUX2_X1 U2871 ( .A(\REGISTERS[19][10] ), .B(n3199), .S(n2), .Z(n1534) );
  MUX2_X1 U2872 ( .A(\REGISTERS[19][9] ), .B(n3200), .S(n2), .Z(n1533) );
  MUX2_X1 U2873 ( .A(\REGISTERS[19][8] ), .B(n3201), .S(n2), .Z(n1532) );
  MUX2_X1 U2874 ( .A(\REGISTERS[19][7] ), .B(n3202), .S(n2), .Z(n1531) );
  MUX2_X1 U2875 ( .A(\REGISTERS[19][6] ), .B(n3203), .S(n2), .Z(n1530) );
  MUX2_X1 U2876 ( .A(\REGISTERS[19][5] ), .B(n3204), .S(n2), .Z(n1529) );
  MUX2_X1 U2877 ( .A(\REGISTERS[19][4] ), .B(n3205), .S(n2), .Z(n1528) );
  MUX2_X1 U2878 ( .A(\REGISTERS[19][3] ), .B(n3206), .S(n2), .Z(n1527) );
  MUX2_X1 U2879 ( .A(\REGISTERS[19][2] ), .B(n3207), .S(n2), .Z(n1526) );
  MUX2_X1 U2880 ( .A(\REGISTERS[19][1] ), .B(n3208), .S(n2), .Z(n1525) );
  MUX2_X1 U2881 ( .A(\REGISTERS[19][0] ), .B(n3209), .S(n2), .Z(n1524) );
  OAI21_X1 U2882 ( .B1(n3218), .B2(n3240), .A(n3212), .ZN(n3243) );
  MUX2_X1 U2883 ( .A(\REGISTERS[20][31] ), .B(n3177), .S(n4), .Z(n1523) );
  MUX2_X1 U2884 ( .A(\REGISTERS[20][30] ), .B(n3179), .S(n4), .Z(n1522) );
  MUX2_X1 U2885 ( .A(\REGISTERS[20][29] ), .B(n3180), .S(n4), .Z(n1521) );
  MUX2_X1 U2886 ( .A(\REGISTERS[20][28] ), .B(n3181), .S(n4), .Z(n1520) );
  MUX2_X1 U2887 ( .A(\REGISTERS[20][27] ), .B(n3182), .S(n4), .Z(n1519) );
  MUX2_X1 U2888 ( .A(\REGISTERS[20][26] ), .B(n3183), .S(n4), .Z(n1518) );
  MUX2_X1 U2889 ( .A(\REGISTERS[20][25] ), .B(n3184), .S(n4), .Z(n1517) );
  MUX2_X1 U2890 ( .A(\REGISTERS[20][24] ), .B(n3185), .S(n4), .Z(n1516) );
  MUX2_X1 U2891 ( .A(\REGISTERS[20][23] ), .B(n3186), .S(n4), .Z(n1515) );
  MUX2_X1 U2892 ( .A(\REGISTERS[20][22] ), .B(n3187), .S(n4), .Z(n1514) );
  MUX2_X1 U2893 ( .A(\REGISTERS[20][21] ), .B(n3188), .S(n4), .Z(n1513) );
  MUX2_X1 U2894 ( .A(\REGISTERS[20][20] ), .B(n3189), .S(n4), .Z(n1512) );
  MUX2_X1 U2895 ( .A(\REGISTERS[20][19] ), .B(n3190), .S(n4), .Z(n1511) );
  MUX2_X1 U2896 ( .A(\REGISTERS[20][18] ), .B(n3191), .S(n4), .Z(n1510) );
  MUX2_X1 U2897 ( .A(\REGISTERS[20][17] ), .B(n3192), .S(n4), .Z(n1509) );
  MUX2_X1 U2898 ( .A(\REGISTERS[20][16] ), .B(n3193), .S(n4), .Z(n1508) );
  MUX2_X1 U2899 ( .A(\REGISTERS[20][15] ), .B(n3194), .S(n4), .Z(n1507) );
  MUX2_X1 U2900 ( .A(\REGISTERS[20][14] ), .B(n3195), .S(n4), .Z(n1506) );
  MUX2_X1 U2901 ( .A(\REGISTERS[20][13] ), .B(n3196), .S(n4), .Z(n1505) );
  MUX2_X1 U2902 ( .A(\REGISTERS[20][12] ), .B(n3197), .S(n4), .Z(n1504) );
  MUX2_X1 U2903 ( .A(\REGISTERS[20][11] ), .B(n3198), .S(n4), .Z(n1503) );
  MUX2_X1 U2904 ( .A(\REGISTERS[20][10] ), .B(n3199), .S(n4), .Z(n1502) );
  MUX2_X1 U2905 ( .A(\REGISTERS[20][9] ), .B(n3200), .S(n4), .Z(n1501) );
  MUX2_X1 U2906 ( .A(\REGISTERS[20][8] ), .B(n3201), .S(n4), .Z(n1500) );
  MUX2_X1 U2907 ( .A(\REGISTERS[20][7] ), .B(n3202), .S(n4), .Z(n1499) );
  MUX2_X1 U2908 ( .A(\REGISTERS[20][6] ), .B(n3203), .S(n4), .Z(n1498) );
  MUX2_X1 U2909 ( .A(\REGISTERS[20][5] ), .B(n3204), .S(n4), .Z(n1497) );
  MUX2_X1 U2910 ( .A(\REGISTERS[20][4] ), .B(n3205), .S(n4), .Z(n1496) );
  MUX2_X1 U2911 ( .A(\REGISTERS[20][3] ), .B(n3206), .S(n4), .Z(n1495) );
  MUX2_X1 U2912 ( .A(\REGISTERS[20][2] ), .B(n3207), .S(n4), .Z(n1494) );
  MUX2_X1 U2913 ( .A(\REGISTERS[20][1] ), .B(n3208), .S(n4), .Z(n1493) );
  MUX2_X1 U2914 ( .A(\REGISTERS[20][0] ), .B(n3209), .S(n4), .Z(n1492) );
  OAI21_X1 U2915 ( .B1(n3220), .B2(n3240), .A(n3212), .ZN(n3244) );
  MUX2_X1 U2916 ( .A(\REGISTERS[21][31] ), .B(n3177), .S(n6), .Z(n1491) );
  MUX2_X1 U2917 ( .A(\REGISTERS[21][30] ), .B(n3179), .S(n6), .Z(n1490) );
  MUX2_X1 U2918 ( .A(\REGISTERS[21][29] ), .B(n3180), .S(n6), .Z(n1489) );
  MUX2_X1 U2919 ( .A(\REGISTERS[21][28] ), .B(n3181), .S(n6), .Z(n1488) );
  MUX2_X1 U2920 ( .A(\REGISTERS[21][27] ), .B(n3182), .S(n6), .Z(n1487) );
  MUX2_X1 U2921 ( .A(\REGISTERS[21][26] ), .B(n3183), .S(n6), .Z(n1486) );
  MUX2_X1 U2922 ( .A(\REGISTERS[21][25] ), .B(n3184), .S(n6), .Z(n1485) );
  MUX2_X1 U2923 ( .A(\REGISTERS[21][24] ), .B(n3185), .S(n6), .Z(n1484) );
  MUX2_X1 U2924 ( .A(\REGISTERS[21][23] ), .B(n3186), .S(n6), .Z(n1483) );
  MUX2_X1 U2925 ( .A(\REGISTERS[21][22] ), .B(n3187), .S(n6), .Z(n1482) );
  MUX2_X1 U2926 ( .A(\REGISTERS[21][21] ), .B(n3188), .S(n6), .Z(n1481) );
  MUX2_X1 U2927 ( .A(\REGISTERS[21][20] ), .B(n3189), .S(n6), .Z(n1480) );
  MUX2_X1 U2928 ( .A(\REGISTERS[21][19] ), .B(n3190), .S(n6), .Z(n1479) );
  MUX2_X1 U2929 ( .A(\REGISTERS[21][18] ), .B(n3191), .S(n6), .Z(n1478) );
  MUX2_X1 U2930 ( .A(\REGISTERS[21][17] ), .B(n3192), .S(n6), .Z(n1477) );
  MUX2_X1 U2931 ( .A(\REGISTERS[21][16] ), .B(n3193), .S(n6), .Z(n1476) );
  MUX2_X1 U2932 ( .A(\REGISTERS[21][15] ), .B(n3194), .S(n6), .Z(n1475) );
  MUX2_X1 U2933 ( .A(\REGISTERS[21][14] ), .B(n3195), .S(n6), .Z(n1474) );
  MUX2_X1 U2934 ( .A(\REGISTERS[21][13] ), .B(n3196), .S(n6), .Z(n1473) );
  MUX2_X1 U2935 ( .A(\REGISTERS[21][12] ), .B(n3197), .S(n6), .Z(n1472) );
  MUX2_X1 U2936 ( .A(\REGISTERS[21][11] ), .B(n3198), .S(n6), .Z(n1471) );
  MUX2_X1 U2937 ( .A(\REGISTERS[21][10] ), .B(n3199), .S(n6), .Z(n1470) );
  MUX2_X1 U2938 ( .A(\REGISTERS[21][9] ), .B(n3200), .S(n6), .Z(n1469) );
  MUX2_X1 U2939 ( .A(\REGISTERS[21][8] ), .B(n3201), .S(n6), .Z(n1468) );
  MUX2_X1 U2940 ( .A(\REGISTERS[21][7] ), .B(n3202), .S(n6), .Z(n1467) );
  MUX2_X1 U2941 ( .A(\REGISTERS[21][6] ), .B(n3203), .S(n6), .Z(n1466) );
  MUX2_X1 U2942 ( .A(\REGISTERS[21][5] ), .B(n3204), .S(n6), .Z(n1465) );
  MUX2_X1 U2943 ( .A(\REGISTERS[21][4] ), .B(n3205), .S(n6), .Z(n1464) );
  MUX2_X1 U2944 ( .A(\REGISTERS[21][3] ), .B(n3206), .S(n6), .Z(n1463) );
  MUX2_X1 U2945 ( .A(\REGISTERS[21][2] ), .B(n3207), .S(n6), .Z(n1462) );
  MUX2_X1 U2946 ( .A(\REGISTERS[21][1] ), .B(n3208), .S(n6), .Z(n1461) );
  MUX2_X1 U2947 ( .A(\REGISTERS[21][0] ), .B(n3209), .S(n6), .Z(n1460) );
  OAI21_X1 U2948 ( .B1(n3222), .B2(n3240), .A(n3212), .ZN(n3245) );
  MUX2_X1 U2949 ( .A(\REGISTERS[22][31] ), .B(n3177), .S(n8), .Z(n1459) );
  MUX2_X1 U2950 ( .A(\REGISTERS[22][30] ), .B(n3179), .S(n8), .Z(n1458) );
  MUX2_X1 U2951 ( .A(\REGISTERS[22][29] ), .B(n3180), .S(n8), .Z(n1457) );
  MUX2_X1 U2952 ( .A(\REGISTERS[22][28] ), .B(n3181), .S(n8), .Z(n1456) );
  MUX2_X1 U2953 ( .A(\REGISTERS[22][27] ), .B(n3182), .S(n8), .Z(n1455) );
  MUX2_X1 U2954 ( .A(\REGISTERS[22][26] ), .B(n3183), .S(n8), .Z(n1454) );
  MUX2_X1 U2955 ( .A(\REGISTERS[22][25] ), .B(n3184), .S(n8), .Z(n1453) );
  MUX2_X1 U2956 ( .A(\REGISTERS[22][24] ), .B(n3185), .S(n8), .Z(n1452) );
  MUX2_X1 U2957 ( .A(\REGISTERS[22][23] ), .B(n3186), .S(n8), .Z(n1451) );
  MUX2_X1 U2958 ( .A(\REGISTERS[22][22] ), .B(n3187), .S(n8), .Z(n1450) );
  MUX2_X1 U2959 ( .A(\REGISTERS[22][21] ), .B(n3188), .S(n8), .Z(n1449) );
  MUX2_X1 U2960 ( .A(\REGISTERS[22][20] ), .B(n3189), .S(n8), .Z(n1448) );
  MUX2_X1 U2961 ( .A(\REGISTERS[22][19] ), .B(n3190), .S(n8), .Z(n1447) );
  MUX2_X1 U2962 ( .A(\REGISTERS[22][18] ), .B(n3191), .S(n8), .Z(n1446) );
  MUX2_X1 U2963 ( .A(\REGISTERS[22][17] ), .B(n3192), .S(n8), .Z(n1445) );
  MUX2_X1 U2964 ( .A(\REGISTERS[22][16] ), .B(n3193), .S(n8), .Z(n1444) );
  MUX2_X1 U2965 ( .A(\REGISTERS[22][15] ), .B(n3194), .S(n8), .Z(n1443) );
  MUX2_X1 U2966 ( .A(\REGISTERS[22][14] ), .B(n3195), .S(n8), .Z(n1442) );
  MUX2_X1 U2967 ( .A(\REGISTERS[22][13] ), .B(n3196), .S(n8), .Z(n1441) );
  MUX2_X1 U2968 ( .A(\REGISTERS[22][12] ), .B(n3197), .S(n8), .Z(n1440) );
  MUX2_X1 U2969 ( .A(\REGISTERS[22][11] ), .B(n3198), .S(n8), .Z(n1439) );
  MUX2_X1 U2970 ( .A(\REGISTERS[22][10] ), .B(n3199), .S(n8), .Z(n1438) );
  MUX2_X1 U2971 ( .A(\REGISTERS[22][9] ), .B(n3200), .S(n8), .Z(n1437) );
  MUX2_X1 U2972 ( .A(\REGISTERS[22][8] ), .B(n3201), .S(n8), .Z(n1436) );
  MUX2_X1 U2973 ( .A(\REGISTERS[22][7] ), .B(n3202), .S(n8), .Z(n1435) );
  MUX2_X1 U2974 ( .A(\REGISTERS[22][6] ), .B(n3203), .S(n8), .Z(n1434) );
  MUX2_X1 U2975 ( .A(\REGISTERS[22][5] ), .B(n3204), .S(n8), .Z(n1433) );
  MUX2_X1 U2976 ( .A(\REGISTERS[22][4] ), .B(n3205), .S(n8), .Z(n1432) );
  MUX2_X1 U2977 ( .A(\REGISTERS[22][3] ), .B(n3206), .S(n8), .Z(n1431) );
  MUX2_X1 U2978 ( .A(\REGISTERS[22][2] ), .B(n3207), .S(n8), .Z(n1430) );
  MUX2_X1 U2979 ( .A(\REGISTERS[22][1] ), .B(n3208), .S(n8), .Z(n1429) );
  MUX2_X1 U2980 ( .A(\REGISTERS[22][0] ), .B(n3209), .S(n8), .Z(n1428) );
  OAI21_X1 U2981 ( .B1(n3224), .B2(n3240), .A(n3212), .ZN(n3246) );
  MUX2_X1 U2982 ( .A(\REGISTERS[23][31] ), .B(n3177), .S(n10), .Z(n1427) );
  MUX2_X1 U2983 ( .A(\REGISTERS[23][30] ), .B(n3179), .S(n10), .Z(n1426) );
  MUX2_X1 U2984 ( .A(\REGISTERS[23][29] ), .B(n3180), .S(n10), .Z(n1425) );
  MUX2_X1 U2985 ( .A(\REGISTERS[23][28] ), .B(n3181), .S(n10), .Z(n1424) );
  MUX2_X1 U2986 ( .A(\REGISTERS[23][27] ), .B(n3182), .S(n10), .Z(n1423) );
  MUX2_X1 U2987 ( .A(\REGISTERS[23][26] ), .B(n3183), .S(n10), .Z(n1422) );
  MUX2_X1 U2988 ( .A(\REGISTERS[23][25] ), .B(n3184), .S(n10), .Z(n1421) );
  MUX2_X1 U2989 ( .A(\REGISTERS[23][24] ), .B(n3185), .S(n10), .Z(n1420) );
  MUX2_X1 U2990 ( .A(\REGISTERS[23][23] ), .B(n3186), .S(n10), .Z(n1419) );
  MUX2_X1 U2991 ( .A(\REGISTERS[23][22] ), .B(n3187), .S(n10), .Z(n1418) );
  MUX2_X1 U2992 ( .A(\REGISTERS[23][21] ), .B(n3188), .S(n10), .Z(n1417) );
  MUX2_X1 U2993 ( .A(\REGISTERS[23][20] ), .B(n3189), .S(n10), .Z(n1416) );
  MUX2_X1 U2994 ( .A(\REGISTERS[23][19] ), .B(n3190), .S(n10), .Z(n1415) );
  MUX2_X1 U2995 ( .A(\REGISTERS[23][18] ), .B(n3191), .S(n10), .Z(n1414) );
  MUX2_X1 U2996 ( .A(\REGISTERS[23][17] ), .B(n3192), .S(n10), .Z(n1413) );
  MUX2_X1 U2997 ( .A(\REGISTERS[23][16] ), .B(n3193), .S(n10), .Z(n1412) );
  MUX2_X1 U2998 ( .A(\REGISTERS[23][15] ), .B(n3194), .S(n10), .Z(n1411) );
  MUX2_X1 U2999 ( .A(\REGISTERS[23][14] ), .B(n3195), .S(n10), .Z(n1410) );
  MUX2_X1 U3000 ( .A(\REGISTERS[23][13] ), .B(n3196), .S(n10), .Z(n1409) );
  MUX2_X1 U3001 ( .A(\REGISTERS[23][12] ), .B(n3197), .S(n10), .Z(n1408) );
  MUX2_X1 U3002 ( .A(\REGISTERS[23][11] ), .B(n3198), .S(n10), .Z(n1407) );
  MUX2_X1 U3003 ( .A(\REGISTERS[23][10] ), .B(n3199), .S(n10), .Z(n1406) );
  MUX2_X1 U3004 ( .A(\REGISTERS[23][9] ), .B(n3200), .S(n10), .Z(n1405) );
  MUX2_X1 U3005 ( .A(\REGISTERS[23][8] ), .B(n3201), .S(n10), .Z(n1404) );
  MUX2_X1 U3006 ( .A(\REGISTERS[23][7] ), .B(n3202), .S(n10), .Z(n1403) );
  MUX2_X1 U3007 ( .A(\REGISTERS[23][6] ), .B(n3203), .S(n10), .Z(n1402) );
  MUX2_X1 U3008 ( .A(\REGISTERS[23][5] ), .B(n3204), .S(n10), .Z(n1401) );
  MUX2_X1 U3009 ( .A(\REGISTERS[23][4] ), .B(n3205), .S(n10), .Z(n1400) );
  MUX2_X1 U3010 ( .A(\REGISTERS[23][3] ), .B(n3206), .S(n10), .Z(n1399) );
  MUX2_X1 U3011 ( .A(\REGISTERS[23][2] ), .B(n3207), .S(n10), .Z(n1398) );
  MUX2_X1 U3012 ( .A(\REGISTERS[23][1] ), .B(n3208), .S(n10), .Z(n1397) );
  MUX2_X1 U3013 ( .A(\REGISTERS[23][0] ), .B(n3209), .S(n10), .Z(n1396) );
  OAI21_X1 U3014 ( .B1(n3226), .B2(n3240), .A(n3212), .ZN(n3247) );
  NAND3_X1 U3015 ( .A1(n3229), .A2(n3227), .A3(ADD_WR[4]), .ZN(n3240) );
  INV_X1 U3016 ( .A(ADD_WR[3]), .ZN(n3227) );
  MUX2_X1 U3017 ( .A(\REGISTERS[24][31] ), .B(n3177), .S(n12), .Z(n1395) );
  MUX2_X1 U3018 ( .A(\REGISTERS[24][30] ), .B(n3179), .S(n12), .Z(n1394) );
  MUX2_X1 U3019 ( .A(\REGISTERS[24][29] ), .B(n3180), .S(n12), .Z(n1393) );
  MUX2_X1 U3020 ( .A(\REGISTERS[24][28] ), .B(n3181), .S(n12), .Z(n1392) );
  MUX2_X1 U3021 ( .A(\REGISTERS[24][27] ), .B(n3182), .S(n12), .Z(n1391) );
  MUX2_X1 U3022 ( .A(\REGISTERS[24][26] ), .B(n3183), .S(n12), .Z(n1390) );
  MUX2_X1 U3023 ( .A(\REGISTERS[24][25] ), .B(n3184), .S(n12), .Z(n1389) );
  MUX2_X1 U3024 ( .A(\REGISTERS[24][24] ), .B(n3185), .S(n12), .Z(n1388) );
  MUX2_X1 U3025 ( .A(\REGISTERS[24][23] ), .B(n3186), .S(n12), .Z(n1387) );
  MUX2_X1 U3026 ( .A(\REGISTERS[24][22] ), .B(n3187), .S(n12), .Z(n1386) );
  MUX2_X1 U3027 ( .A(\REGISTERS[24][21] ), .B(n3188), .S(n12), .Z(n1385) );
  MUX2_X1 U3028 ( .A(\REGISTERS[24][20] ), .B(n3189), .S(n12), .Z(n1384) );
  MUX2_X1 U3029 ( .A(\REGISTERS[24][19] ), .B(n3190), .S(n12), .Z(n1383) );
  MUX2_X1 U3030 ( .A(\REGISTERS[24][18] ), .B(n3191), .S(n12), .Z(n1382) );
  MUX2_X1 U3031 ( .A(\REGISTERS[24][17] ), .B(n3192), .S(n12), .Z(n1381) );
  MUX2_X1 U3032 ( .A(\REGISTERS[24][16] ), .B(n3193), .S(n12), .Z(n1380) );
  MUX2_X1 U3033 ( .A(\REGISTERS[24][15] ), .B(n3194), .S(n12), .Z(n1379) );
  MUX2_X1 U3034 ( .A(\REGISTERS[24][14] ), .B(n3195), .S(n12), .Z(n1378) );
  MUX2_X1 U3035 ( .A(\REGISTERS[24][13] ), .B(n3196), .S(n12), .Z(n1377) );
  MUX2_X1 U3036 ( .A(\REGISTERS[24][12] ), .B(n3197), .S(n12), .Z(n1376) );
  MUX2_X1 U3037 ( .A(\REGISTERS[24][11] ), .B(n3198), .S(n12), .Z(n1375) );
  MUX2_X1 U3038 ( .A(\REGISTERS[24][10] ), .B(n3199), .S(n12), .Z(n1374) );
  MUX2_X1 U3039 ( .A(\REGISTERS[24][9] ), .B(n3200), .S(n12), .Z(n1373) );
  MUX2_X1 U3040 ( .A(\REGISTERS[24][8] ), .B(n3201), .S(n12), .Z(n1372) );
  MUX2_X1 U3041 ( .A(\REGISTERS[24][7] ), .B(n3202), .S(n12), .Z(n1371) );
  MUX2_X1 U3042 ( .A(\REGISTERS[24][6] ), .B(n3203), .S(n12), .Z(n1370) );
  MUX2_X1 U3043 ( .A(\REGISTERS[24][5] ), .B(n3204), .S(n12), .Z(n1369) );
  MUX2_X1 U3044 ( .A(\REGISTERS[24][4] ), .B(n3205), .S(n12), .Z(n1368) );
  MUX2_X1 U3045 ( .A(\REGISTERS[24][3] ), .B(n3206), .S(n12), .Z(n1367) );
  MUX2_X1 U3046 ( .A(\REGISTERS[24][2] ), .B(n3207), .S(n12), .Z(n1366) );
  MUX2_X1 U3047 ( .A(\REGISTERS[24][1] ), .B(n3208), .S(n12), .Z(n1365) );
  MUX2_X1 U3048 ( .A(\REGISTERS[24][0] ), .B(n3209), .S(n12), .Z(n1364) );
  OAI21_X1 U3049 ( .B1(n3211), .B2(n3249), .A(n3212), .ZN(n3248) );
  NAND3_X1 U3050 ( .A1(n3250), .A2(n3251), .A3(n3252), .ZN(n3211) );
  MUX2_X1 U3051 ( .A(\REGISTERS[25][31] ), .B(n3177), .S(n14), .Z(n1363) );
  MUX2_X1 U3052 ( .A(\REGISTERS[25][30] ), .B(n3179), .S(n14), .Z(n1362) );
  MUX2_X1 U3053 ( .A(\REGISTERS[25][29] ), .B(n3180), .S(n14), .Z(n1361) );
  MUX2_X1 U3054 ( .A(\REGISTERS[25][28] ), .B(n3181), .S(n14), .Z(n1360) );
  MUX2_X1 U3055 ( .A(\REGISTERS[25][27] ), .B(n3182), .S(n14), .Z(n1359) );
  MUX2_X1 U3056 ( .A(\REGISTERS[25][26] ), .B(n3183), .S(n14), .Z(n1358) );
  MUX2_X1 U3057 ( .A(\REGISTERS[25][25] ), .B(n3184), .S(n14), .Z(n1357) );
  MUX2_X1 U3058 ( .A(\REGISTERS[25][24] ), .B(n3185), .S(n14), .Z(n1356) );
  MUX2_X1 U3059 ( .A(\REGISTERS[25][23] ), .B(n3186), .S(n14), .Z(n1355) );
  MUX2_X1 U3060 ( .A(\REGISTERS[25][22] ), .B(n3187), .S(n14), .Z(n1354) );
  MUX2_X1 U3061 ( .A(\REGISTERS[25][21] ), .B(n3188), .S(n14), .Z(n1353) );
  MUX2_X1 U3062 ( .A(\REGISTERS[25][20] ), .B(n3189), .S(n14), .Z(n1352) );
  MUX2_X1 U3063 ( .A(\REGISTERS[25][19] ), .B(n3190), .S(n14), .Z(n1351) );
  MUX2_X1 U3064 ( .A(\REGISTERS[25][18] ), .B(n3191), .S(n14), .Z(n1350) );
  MUX2_X1 U3065 ( .A(\REGISTERS[25][17] ), .B(n3192), .S(n14), .Z(n1349) );
  MUX2_X1 U3066 ( .A(\REGISTERS[25][16] ), .B(n3193), .S(n14), .Z(n1348) );
  MUX2_X1 U3067 ( .A(\REGISTERS[25][15] ), .B(n3194), .S(n14), .Z(n1347) );
  MUX2_X1 U3068 ( .A(\REGISTERS[25][14] ), .B(n3195), .S(n14), .Z(n1346) );
  MUX2_X1 U3069 ( .A(\REGISTERS[25][13] ), .B(n3196), .S(n14), .Z(n1345) );
  MUX2_X1 U3070 ( .A(\REGISTERS[25][12] ), .B(n3197), .S(n14), .Z(n1344) );
  MUX2_X1 U3071 ( .A(\REGISTERS[25][11] ), .B(n3198), .S(n14), .Z(n1343) );
  MUX2_X1 U3072 ( .A(\REGISTERS[25][10] ), .B(n3199), .S(n14), .Z(n1342) );
  MUX2_X1 U3073 ( .A(\REGISTERS[25][9] ), .B(n3200), .S(n14), .Z(n1341) );
  MUX2_X1 U3074 ( .A(\REGISTERS[25][8] ), .B(n3201), .S(n14), .Z(n1340) );
  MUX2_X1 U3075 ( .A(\REGISTERS[25][7] ), .B(n3202), .S(n14), .Z(n1339) );
  MUX2_X1 U3076 ( .A(\REGISTERS[25][6] ), .B(n3203), .S(n14), .Z(n1338) );
  MUX2_X1 U3077 ( .A(\REGISTERS[25][5] ), .B(n3204), .S(n14), .Z(n1337) );
  MUX2_X1 U3078 ( .A(\REGISTERS[25][4] ), .B(n3205), .S(n14), .Z(n1336) );
  MUX2_X1 U3079 ( .A(\REGISTERS[25][3] ), .B(n3206), .S(n14), .Z(n1335) );
  MUX2_X1 U3080 ( .A(\REGISTERS[25][2] ), .B(n3207), .S(n14), .Z(n1334) );
  MUX2_X1 U3081 ( .A(\REGISTERS[25][1] ), .B(n3208), .S(n14), .Z(n1333) );
  MUX2_X1 U3082 ( .A(\REGISTERS[25][0] ), .B(n3209), .S(n14), .Z(n1332) );
  OAI21_X1 U3083 ( .B1(n3214), .B2(n3249), .A(n3212), .ZN(n3253) );
  NAND3_X1 U3084 ( .A1(n3250), .A2(n3251), .A3(ADD_WR[0]), .ZN(n3214) );
  MUX2_X1 U3085 ( .A(\REGISTERS[26][31] ), .B(n3177), .S(n16), .Z(n1331) );
  MUX2_X1 U3086 ( .A(\REGISTERS[26][30] ), .B(n3179), .S(n16), .Z(n1330) );
  MUX2_X1 U3087 ( .A(\REGISTERS[26][29] ), .B(n3180), .S(n16), .Z(n1329) );
  MUX2_X1 U3088 ( .A(\REGISTERS[26][28] ), .B(n3181), .S(n16), .Z(n1328) );
  MUX2_X1 U3089 ( .A(\REGISTERS[26][27] ), .B(n3182), .S(n16), .Z(n1327) );
  MUX2_X1 U3090 ( .A(\REGISTERS[26][26] ), .B(n3183), .S(n16), .Z(n1326) );
  MUX2_X1 U3091 ( .A(\REGISTERS[26][25] ), .B(n3184), .S(n16), .Z(n1325) );
  MUX2_X1 U3092 ( .A(\REGISTERS[26][24] ), .B(n3185), .S(n16), .Z(n1324) );
  MUX2_X1 U3093 ( .A(\REGISTERS[26][23] ), .B(n3186), .S(n16), .Z(n1323) );
  MUX2_X1 U3094 ( .A(\REGISTERS[26][22] ), .B(n3187), .S(n16), .Z(n1322) );
  MUX2_X1 U3095 ( .A(\REGISTERS[26][21] ), .B(n3188), .S(n16), .Z(n1321) );
  MUX2_X1 U3096 ( .A(\REGISTERS[26][20] ), .B(n3189), .S(n16), .Z(n1320) );
  MUX2_X1 U3097 ( .A(\REGISTERS[26][19] ), .B(n3190), .S(n16), .Z(n1319) );
  MUX2_X1 U3098 ( .A(\REGISTERS[26][18] ), .B(n3191), .S(n16), .Z(n1318) );
  MUX2_X1 U3099 ( .A(\REGISTERS[26][17] ), .B(n3192), .S(n16), .Z(n1317) );
  MUX2_X1 U3100 ( .A(\REGISTERS[26][16] ), .B(n3193), .S(n16), .Z(n1316) );
  MUX2_X1 U3101 ( .A(\REGISTERS[26][15] ), .B(n3194), .S(n16), .Z(n1315) );
  MUX2_X1 U3102 ( .A(\REGISTERS[26][14] ), .B(n3195), .S(n16), .Z(n1314) );
  MUX2_X1 U3103 ( .A(\REGISTERS[26][13] ), .B(n3196), .S(n16), .Z(n1313) );
  MUX2_X1 U3104 ( .A(\REGISTERS[26][12] ), .B(n3197), .S(n16), .Z(n1312) );
  MUX2_X1 U3105 ( .A(\REGISTERS[26][11] ), .B(n3198), .S(n16), .Z(n1311) );
  MUX2_X1 U3106 ( .A(\REGISTERS[26][10] ), .B(n3199), .S(n16), .Z(n1310) );
  MUX2_X1 U3107 ( .A(\REGISTERS[26][9] ), .B(n3200), .S(n16), .Z(n1309) );
  MUX2_X1 U3108 ( .A(\REGISTERS[26][8] ), .B(n3201), .S(n16), .Z(n1308) );
  MUX2_X1 U3109 ( .A(\REGISTERS[26][7] ), .B(n3202), .S(n16), .Z(n1307) );
  MUX2_X1 U3110 ( .A(\REGISTERS[26][6] ), .B(n3203), .S(n16), .Z(n1306) );
  MUX2_X1 U3111 ( .A(\REGISTERS[26][5] ), .B(n3204), .S(n16), .Z(n1305) );
  MUX2_X1 U3112 ( .A(\REGISTERS[26][4] ), .B(n3205), .S(n16), .Z(n1304) );
  MUX2_X1 U3113 ( .A(\REGISTERS[26][3] ), .B(n3206), .S(n16), .Z(n1303) );
  MUX2_X1 U3114 ( .A(\REGISTERS[26][2] ), .B(n3207), .S(n16), .Z(n1302) );
  MUX2_X1 U3115 ( .A(\REGISTERS[26][1] ), .B(n3208), .S(n16), .Z(n1301) );
  MUX2_X1 U3116 ( .A(\REGISTERS[26][0] ), .B(n3209), .S(n16), .Z(n1300) );
  OAI21_X1 U3117 ( .B1(n3216), .B2(n3249), .A(n3212), .ZN(n3254) );
  NAND3_X1 U3118 ( .A1(n3252), .A2(n3251), .A3(ADD_WR[1]), .ZN(n3216) );
  MUX2_X1 U3119 ( .A(\REGISTERS[27][31] ), .B(n3177), .S(n18), .Z(n1299) );
  MUX2_X1 U3120 ( .A(\REGISTERS[27][30] ), .B(n3179), .S(n18), .Z(n1298) );
  MUX2_X1 U3121 ( .A(\REGISTERS[27][29] ), .B(n3180), .S(n18), .Z(n1297) );
  MUX2_X1 U3122 ( .A(\REGISTERS[27][28] ), .B(n3181), .S(n18), .Z(n1296) );
  MUX2_X1 U3123 ( .A(\REGISTERS[27][27] ), .B(n3182), .S(n18), .Z(n1295) );
  MUX2_X1 U3124 ( .A(\REGISTERS[27][26] ), .B(n3183), .S(n18), .Z(n1294) );
  MUX2_X1 U3125 ( .A(\REGISTERS[27][25] ), .B(n3184), .S(n18), .Z(n1293) );
  MUX2_X1 U3126 ( .A(\REGISTERS[27][24] ), .B(n3185), .S(n18), .Z(n1292) );
  MUX2_X1 U3127 ( .A(\REGISTERS[27][23] ), .B(n3186), .S(n18), .Z(n1291) );
  MUX2_X1 U3128 ( .A(\REGISTERS[27][22] ), .B(n3187), .S(n18), .Z(n1290) );
  MUX2_X1 U3129 ( .A(\REGISTERS[27][21] ), .B(n3188), .S(n18), .Z(n1289) );
  MUX2_X1 U3130 ( .A(\REGISTERS[27][20] ), .B(n3189), .S(n18), .Z(n1288) );
  MUX2_X1 U3131 ( .A(\REGISTERS[27][19] ), .B(n3190), .S(n18), .Z(n1287) );
  MUX2_X1 U3132 ( .A(\REGISTERS[27][18] ), .B(n3191), .S(n18), .Z(n1286) );
  MUX2_X1 U3133 ( .A(\REGISTERS[27][17] ), .B(n3192), .S(n18), .Z(n1285) );
  MUX2_X1 U3134 ( .A(\REGISTERS[27][16] ), .B(n3193), .S(n18), .Z(n1284) );
  MUX2_X1 U3135 ( .A(\REGISTERS[27][15] ), .B(n3194), .S(n18), .Z(n1283) );
  MUX2_X1 U3136 ( .A(\REGISTERS[27][14] ), .B(n3195), .S(n18), .Z(n1282) );
  MUX2_X1 U3137 ( .A(\REGISTERS[27][13] ), .B(n3196), .S(n18), .Z(n1281) );
  MUX2_X1 U3138 ( .A(\REGISTERS[27][12] ), .B(n3197), .S(n18), .Z(n1280) );
  MUX2_X1 U3139 ( .A(\REGISTERS[27][11] ), .B(n3198), .S(n18), .Z(n1279) );
  MUX2_X1 U3140 ( .A(\REGISTERS[27][10] ), .B(n3199), .S(n18), .Z(n1278) );
  MUX2_X1 U3141 ( .A(\REGISTERS[27][9] ), .B(n3200), .S(n18), .Z(n1277) );
  MUX2_X1 U3142 ( .A(\REGISTERS[27][8] ), .B(n3201), .S(n18), .Z(n1276) );
  MUX2_X1 U3143 ( .A(\REGISTERS[27][7] ), .B(n3202), .S(n18), .Z(n1275) );
  MUX2_X1 U3144 ( .A(\REGISTERS[27][6] ), .B(n3203), .S(n18), .Z(n1274) );
  MUX2_X1 U3145 ( .A(\REGISTERS[27][5] ), .B(n3204), .S(n18), .Z(n1273) );
  MUX2_X1 U3146 ( .A(\REGISTERS[27][4] ), .B(n3205), .S(n18), .Z(n1272) );
  MUX2_X1 U3147 ( .A(\REGISTERS[27][3] ), .B(n3206), .S(n18), .Z(n1271) );
  MUX2_X1 U3148 ( .A(\REGISTERS[27][2] ), .B(n3207), .S(n18), .Z(n1270) );
  MUX2_X1 U3149 ( .A(\REGISTERS[27][1] ), .B(n3208), .S(n18), .Z(n1269) );
  MUX2_X1 U3150 ( .A(\REGISTERS[27][0] ), .B(n3209), .S(n18), .Z(n1268) );
  OAI21_X1 U3151 ( .B1(n3218), .B2(n3249), .A(n3212), .ZN(n3255) );
  NAND3_X1 U3152 ( .A1(ADD_WR[0]), .A2(n3251), .A3(ADD_WR[1]), .ZN(n3218) );
  INV_X1 U3153 ( .A(ADD_WR[2]), .ZN(n3251) );
  MUX2_X1 U3154 ( .A(\REGISTERS[28][31] ), .B(n3177), .S(n20), .Z(n1267) );
  MUX2_X1 U3155 ( .A(\REGISTERS[28][30] ), .B(n3179), .S(n20), .Z(n1266) );
  MUX2_X1 U3156 ( .A(\REGISTERS[28][29] ), .B(n3180), .S(n20), .Z(n1265) );
  MUX2_X1 U3157 ( .A(\REGISTERS[28][28] ), .B(n3181), .S(n20), .Z(n1264) );
  MUX2_X1 U3158 ( .A(\REGISTERS[28][27] ), .B(n3182), .S(n20), .Z(n1263) );
  MUX2_X1 U3159 ( .A(\REGISTERS[28][26] ), .B(n3183), .S(n20), .Z(n1262) );
  MUX2_X1 U3160 ( .A(\REGISTERS[28][25] ), .B(n3184), .S(n20), .Z(n1261) );
  MUX2_X1 U3161 ( .A(\REGISTERS[28][24] ), .B(n3185), .S(n20), .Z(n1260) );
  MUX2_X1 U3162 ( .A(\REGISTERS[28][23] ), .B(n3186), .S(n20), .Z(n1259) );
  MUX2_X1 U3163 ( .A(\REGISTERS[28][22] ), .B(n3187), .S(n20), .Z(n1258) );
  MUX2_X1 U3164 ( .A(\REGISTERS[28][21] ), .B(n3188), .S(n20), .Z(n1257) );
  MUX2_X1 U3165 ( .A(\REGISTERS[28][20] ), .B(n3189), .S(n20), .Z(n1256) );
  MUX2_X1 U3166 ( .A(\REGISTERS[28][19] ), .B(n3190), .S(n20), .Z(n1255) );
  MUX2_X1 U3167 ( .A(\REGISTERS[28][18] ), .B(n3191), .S(n20), .Z(n1254) );
  MUX2_X1 U3168 ( .A(\REGISTERS[28][17] ), .B(n3192), .S(n20), .Z(n1253) );
  MUX2_X1 U3169 ( .A(\REGISTERS[28][16] ), .B(n3193), .S(n20), .Z(n1252) );
  MUX2_X1 U3170 ( .A(\REGISTERS[28][15] ), .B(n3194), .S(n20), .Z(n1251) );
  MUX2_X1 U3171 ( .A(\REGISTERS[28][14] ), .B(n3195), .S(n20), .Z(n1250) );
  MUX2_X1 U3172 ( .A(\REGISTERS[28][13] ), .B(n3196), .S(n20), .Z(n1249) );
  MUX2_X1 U3173 ( .A(\REGISTERS[28][12] ), .B(n3197), .S(n20), .Z(n1248) );
  MUX2_X1 U3174 ( .A(\REGISTERS[28][11] ), .B(n3198), .S(n20), .Z(n1247) );
  MUX2_X1 U3175 ( .A(\REGISTERS[28][10] ), .B(n3199), .S(n20), .Z(n1246) );
  MUX2_X1 U3176 ( .A(\REGISTERS[28][9] ), .B(n3200), .S(n20), .Z(n1245) );
  MUX2_X1 U3177 ( .A(\REGISTERS[28][8] ), .B(n3201), .S(n20), .Z(n1244) );
  MUX2_X1 U3178 ( .A(\REGISTERS[28][7] ), .B(n3202), .S(n20), .Z(n1243) );
  MUX2_X1 U3179 ( .A(\REGISTERS[28][6] ), .B(n3203), .S(n20), .Z(n1242) );
  MUX2_X1 U3180 ( .A(\REGISTERS[28][5] ), .B(n3204), .S(n20), .Z(n1241) );
  MUX2_X1 U3181 ( .A(\REGISTERS[28][4] ), .B(n3205), .S(n20), .Z(n1240) );
  MUX2_X1 U3182 ( .A(\REGISTERS[28][3] ), .B(n3206), .S(n20), .Z(n1239) );
  MUX2_X1 U3183 ( .A(\REGISTERS[28][2] ), .B(n3207), .S(n20), .Z(n1238) );
  MUX2_X1 U3184 ( .A(\REGISTERS[28][1] ), .B(n3208), .S(n20), .Z(n1237) );
  MUX2_X1 U3185 ( .A(\REGISTERS[28][0] ), .B(n3209), .S(n20), .Z(n1236) );
  OAI21_X1 U3186 ( .B1(n3220), .B2(n3249), .A(n3212), .ZN(n3256) );
  NAND3_X1 U3187 ( .A1(n3252), .A2(n3250), .A3(ADD_WR[2]), .ZN(n3220) );
  MUX2_X1 U3188 ( .A(\REGISTERS[29][31] ), .B(n3177), .S(n22), .Z(n1235) );
  MUX2_X1 U3189 ( .A(\REGISTERS[29][30] ), .B(n3179), .S(n22), .Z(n1234) );
  MUX2_X1 U3190 ( .A(\REGISTERS[29][29] ), .B(n3180), .S(n22), .Z(n1233) );
  MUX2_X1 U3191 ( .A(\REGISTERS[29][28] ), .B(n3181), .S(n22), .Z(n1232) );
  MUX2_X1 U3192 ( .A(\REGISTERS[29][27] ), .B(n3182), .S(n22), .Z(n1231) );
  MUX2_X1 U3193 ( .A(\REGISTERS[29][26] ), .B(n3183), .S(n22), .Z(n1230) );
  MUX2_X1 U3194 ( .A(\REGISTERS[29][25] ), .B(n3184), .S(n22), .Z(n1229) );
  MUX2_X1 U3195 ( .A(\REGISTERS[29][24] ), .B(n3185), .S(n22), .Z(n1228) );
  MUX2_X1 U3196 ( .A(\REGISTERS[29][23] ), .B(n3186), .S(n22), .Z(n1227) );
  MUX2_X1 U3197 ( .A(\REGISTERS[29][22] ), .B(n3187), .S(n22), .Z(n1226) );
  MUX2_X1 U3198 ( .A(\REGISTERS[29][21] ), .B(n3188), .S(n22), .Z(n1225) );
  MUX2_X1 U3199 ( .A(\REGISTERS[29][20] ), .B(n3189), .S(n22), .Z(n1224) );
  MUX2_X1 U3200 ( .A(\REGISTERS[29][19] ), .B(n3190), .S(n22), .Z(n1223) );
  MUX2_X1 U3201 ( .A(\REGISTERS[29][18] ), .B(n3191), .S(n22), .Z(n1222) );
  MUX2_X1 U3202 ( .A(\REGISTERS[29][17] ), .B(n3192), .S(n22), .Z(n1221) );
  MUX2_X1 U3203 ( .A(\REGISTERS[29][16] ), .B(n3193), .S(n22), .Z(n1220) );
  MUX2_X1 U3204 ( .A(\REGISTERS[29][15] ), .B(n3194), .S(n22), .Z(n1219) );
  MUX2_X1 U3205 ( .A(\REGISTERS[29][14] ), .B(n3195), .S(n22), .Z(n1218) );
  MUX2_X1 U3206 ( .A(\REGISTERS[29][13] ), .B(n3196), .S(n22), .Z(n1217) );
  MUX2_X1 U3207 ( .A(\REGISTERS[29][12] ), .B(n3197), .S(n22), .Z(n1216) );
  MUX2_X1 U3208 ( .A(\REGISTERS[29][11] ), .B(n3198), .S(n22), .Z(n1215) );
  MUX2_X1 U3209 ( .A(\REGISTERS[29][10] ), .B(n3199), .S(n22), .Z(n1214) );
  MUX2_X1 U3210 ( .A(\REGISTERS[29][9] ), .B(n3200), .S(n22), .Z(n1213) );
  MUX2_X1 U3211 ( .A(\REGISTERS[29][8] ), .B(n3201), .S(n22), .Z(n1212) );
  MUX2_X1 U3212 ( .A(\REGISTERS[29][7] ), .B(n3202), .S(n22), .Z(n1211) );
  MUX2_X1 U3213 ( .A(\REGISTERS[29][6] ), .B(n3203), .S(n22), .Z(n1210) );
  MUX2_X1 U3214 ( .A(\REGISTERS[29][5] ), .B(n3204), .S(n22), .Z(n1209) );
  MUX2_X1 U3215 ( .A(\REGISTERS[29][4] ), .B(n3205), .S(n22), .Z(n1208) );
  MUX2_X1 U3216 ( .A(\REGISTERS[29][3] ), .B(n3206), .S(n22), .Z(n1207) );
  MUX2_X1 U3217 ( .A(\REGISTERS[29][2] ), .B(n3207), .S(n22), .Z(n1206) );
  MUX2_X1 U3218 ( .A(\REGISTERS[29][1] ), .B(n3208), .S(n22), .Z(n1205) );
  MUX2_X1 U3219 ( .A(\REGISTERS[29][0] ), .B(n3209), .S(n22), .Z(n1204) );
  OAI21_X1 U3220 ( .B1(n3222), .B2(n3249), .A(n3212), .ZN(n3257) );
  NAND3_X1 U3221 ( .A1(ADD_WR[0]), .A2(n3250), .A3(ADD_WR[2]), .ZN(n3222) );
  INV_X1 U3222 ( .A(ADD_WR[1]), .ZN(n3250) );
  MUX2_X1 U3223 ( .A(\REGISTERS[30][31] ), .B(n3177), .S(n24), .Z(n1203) );
  MUX2_X1 U3224 ( .A(\REGISTERS[30][30] ), .B(n3179), .S(n24), .Z(n1202) );
  MUX2_X1 U3225 ( .A(\REGISTERS[30][29] ), .B(n3180), .S(n24), .Z(n1201) );
  MUX2_X1 U3226 ( .A(\REGISTERS[30][28] ), .B(n3181), .S(n24), .Z(n1200) );
  MUX2_X1 U3227 ( .A(\REGISTERS[30][27] ), .B(n3182), .S(n24), .Z(n1199) );
  MUX2_X1 U3228 ( .A(\REGISTERS[30][26] ), .B(n3183), .S(n24), .Z(n1198) );
  MUX2_X1 U3229 ( .A(\REGISTERS[30][25] ), .B(n3184), .S(n24), .Z(n1197) );
  MUX2_X1 U3230 ( .A(\REGISTERS[30][24] ), .B(n3185), .S(n24), .Z(n1196) );
  MUX2_X1 U3231 ( .A(\REGISTERS[30][23] ), .B(n3186), .S(n24), .Z(n1195) );
  MUX2_X1 U3232 ( .A(\REGISTERS[30][22] ), .B(n3187), .S(n24), .Z(n1194) );
  MUX2_X1 U3233 ( .A(\REGISTERS[30][21] ), .B(n3188), .S(n24), .Z(n1193) );
  MUX2_X1 U3234 ( .A(\REGISTERS[30][20] ), .B(n3189), .S(n24), .Z(n1192) );
  MUX2_X1 U3235 ( .A(\REGISTERS[30][19] ), .B(n3190), .S(n24), .Z(n1191) );
  MUX2_X1 U3236 ( .A(\REGISTERS[30][18] ), .B(n3191), .S(n24), .Z(n1190) );
  MUX2_X1 U3237 ( .A(\REGISTERS[30][17] ), .B(n3192), .S(n24), .Z(n1189) );
  MUX2_X1 U3238 ( .A(\REGISTERS[30][16] ), .B(n3193), .S(n24), .Z(n1188) );
  MUX2_X1 U3239 ( .A(\REGISTERS[30][15] ), .B(n3194), .S(n24), .Z(n1187) );
  MUX2_X1 U3240 ( .A(\REGISTERS[30][14] ), .B(n3195), .S(n24), .Z(n1186) );
  MUX2_X1 U3241 ( .A(\REGISTERS[30][13] ), .B(n3196), .S(n24), .Z(n1185) );
  MUX2_X1 U3242 ( .A(\REGISTERS[30][12] ), .B(n3197), .S(n24), .Z(n1184) );
  MUX2_X1 U3243 ( .A(\REGISTERS[30][11] ), .B(n3198), .S(n24), .Z(n1183) );
  MUX2_X1 U3244 ( .A(\REGISTERS[30][10] ), .B(n3199), .S(n24), .Z(n1182) );
  MUX2_X1 U3245 ( .A(\REGISTERS[30][9] ), .B(n3200), .S(n24), .Z(n1181) );
  MUX2_X1 U3246 ( .A(\REGISTERS[30][8] ), .B(n3201), .S(n24), .Z(n1180) );
  MUX2_X1 U3247 ( .A(\REGISTERS[30][7] ), .B(n3202), .S(n24), .Z(n1179) );
  MUX2_X1 U3248 ( .A(\REGISTERS[30][6] ), .B(n3203), .S(n24), .Z(n1178) );
  MUX2_X1 U3249 ( .A(\REGISTERS[30][5] ), .B(n3204), .S(n24), .Z(n1177) );
  MUX2_X1 U3250 ( .A(\REGISTERS[30][4] ), .B(n3205), .S(n24), .Z(n1176) );
  MUX2_X1 U3251 ( .A(\REGISTERS[30][3] ), .B(n3206), .S(n24), .Z(n1175) );
  MUX2_X1 U3252 ( .A(\REGISTERS[30][2] ), .B(n3207), .S(n24), .Z(n1174) );
  MUX2_X1 U3253 ( .A(\REGISTERS[30][1] ), .B(n3208), .S(n24), .Z(n1173) );
  MUX2_X1 U3254 ( .A(\REGISTERS[30][0] ), .B(n3209), .S(n24), .Z(n1172) );
  OAI21_X1 U3255 ( .B1(n3224), .B2(n3249), .A(n3212), .ZN(n3258) );
  NAND3_X1 U3256 ( .A1(ADD_WR[1]), .A2(n3252), .A3(ADD_WR[2]), .ZN(n3224) );
  INV_X1 U3257 ( .A(ADD_WR[0]), .ZN(n3252) );
  MUX2_X1 U3258 ( .A(\REGISTERS[31][31] ), .B(n3177), .S(n26), .Z(n1171) );
  AND2_X1 U3259 ( .A1(DATAIN[31]), .A2(n3212), .ZN(n3177) );
  MUX2_X1 U3260 ( .A(\REGISTERS[31][30] ), .B(n3179), .S(n26), .Z(n1170) );
  AND2_X1 U3261 ( .A1(DATAIN[30]), .A2(n3212), .ZN(n3179) );
  MUX2_X1 U3262 ( .A(\REGISTERS[31][29] ), .B(n3180), .S(n26), .Z(n1169) );
  AND2_X1 U3263 ( .A1(DATAIN[29]), .A2(n3212), .ZN(n3180) );
  MUX2_X1 U3264 ( .A(\REGISTERS[31][28] ), .B(n3181), .S(n26), .Z(n1168) );
  AND2_X1 U3265 ( .A1(DATAIN[28]), .A2(n3212), .ZN(n3181) );
  MUX2_X1 U3266 ( .A(\REGISTERS[31][27] ), .B(n3182), .S(n26), .Z(n1167) );
  AND2_X1 U3267 ( .A1(DATAIN[27]), .A2(n3212), .ZN(n3182) );
  MUX2_X1 U3268 ( .A(\REGISTERS[31][26] ), .B(n3183), .S(n26), .Z(n1166) );
  AND2_X1 U3269 ( .A1(DATAIN[26]), .A2(n3212), .ZN(n3183) );
  MUX2_X1 U3270 ( .A(\REGISTERS[31][25] ), .B(n3184), .S(n26), .Z(n1165) );
  AND2_X1 U3271 ( .A1(DATAIN[25]), .A2(n3212), .ZN(n3184) );
  MUX2_X1 U3272 ( .A(\REGISTERS[31][24] ), .B(n3185), .S(n26), .Z(n1164) );
  AND2_X1 U3273 ( .A1(DATAIN[24]), .A2(n3212), .ZN(n3185) );
  MUX2_X1 U3274 ( .A(\REGISTERS[31][23] ), .B(n3186), .S(n26), .Z(n1163) );
  AND2_X1 U3275 ( .A1(DATAIN[23]), .A2(n3212), .ZN(n3186) );
  MUX2_X1 U3276 ( .A(\REGISTERS[31][22] ), .B(n3187), .S(n26), .Z(n1162) );
  AND2_X1 U3277 ( .A1(DATAIN[22]), .A2(n3212), .ZN(n3187) );
  MUX2_X1 U3278 ( .A(\REGISTERS[31][21] ), .B(n3188), .S(n26), .Z(n1161) );
  AND2_X1 U3279 ( .A1(DATAIN[21]), .A2(n3212), .ZN(n3188) );
  MUX2_X1 U3280 ( .A(\REGISTERS[31][20] ), .B(n3189), .S(n26), .Z(n1160) );
  AND2_X1 U3281 ( .A1(DATAIN[20]), .A2(n3212), .ZN(n3189) );
  MUX2_X1 U3282 ( .A(\REGISTERS[31][19] ), .B(n3190), .S(n26), .Z(n1159) );
  AND2_X1 U3283 ( .A1(DATAIN[19]), .A2(n3212), .ZN(n3190) );
  MUX2_X1 U3284 ( .A(\REGISTERS[31][18] ), .B(n3191), .S(n26), .Z(n1158) );
  AND2_X1 U3285 ( .A1(DATAIN[18]), .A2(n3212), .ZN(n3191) );
  MUX2_X1 U3286 ( .A(\REGISTERS[31][17] ), .B(n3192), .S(n26), .Z(n1157) );
  AND2_X1 U3287 ( .A1(DATAIN[17]), .A2(n3212), .ZN(n3192) );
  MUX2_X1 U3288 ( .A(\REGISTERS[31][16] ), .B(n3193), .S(n26), .Z(n1156) );
  AND2_X1 U3289 ( .A1(DATAIN[16]), .A2(n3212), .ZN(n3193) );
  MUX2_X1 U3290 ( .A(\REGISTERS[31][15] ), .B(n3194), .S(n26), .Z(n1155) );
  AND2_X1 U3291 ( .A1(DATAIN[15]), .A2(n3212), .ZN(n3194) );
  MUX2_X1 U3292 ( .A(\REGISTERS[31][14] ), .B(n3195), .S(n26), .Z(n1154) );
  AND2_X1 U3293 ( .A1(DATAIN[14]), .A2(n3212), .ZN(n3195) );
  MUX2_X1 U3294 ( .A(\REGISTERS[31][13] ), .B(n3196), .S(n26), .Z(n1153) );
  AND2_X1 U3295 ( .A1(DATAIN[13]), .A2(n3212), .ZN(n3196) );
  MUX2_X1 U3296 ( .A(\REGISTERS[31][12] ), .B(n3197), .S(n26), .Z(n1152) );
  AND2_X1 U3297 ( .A1(DATAIN[12]), .A2(n3212), .ZN(n3197) );
  MUX2_X1 U3298 ( .A(\REGISTERS[31][11] ), .B(n3198), .S(n26), .Z(n1151) );
  AND2_X1 U3299 ( .A1(DATAIN[11]), .A2(n3212), .ZN(n3198) );
  MUX2_X1 U3300 ( .A(\REGISTERS[31][10] ), .B(n3199), .S(n26), .Z(n1150) );
  AND2_X1 U3301 ( .A1(DATAIN[10]), .A2(n3212), .ZN(n3199) );
  MUX2_X1 U3302 ( .A(\REGISTERS[31][9] ), .B(n3200), .S(n26), .Z(n1149) );
  AND2_X1 U3303 ( .A1(DATAIN[9]), .A2(n3212), .ZN(n3200) );
  MUX2_X1 U3304 ( .A(\REGISTERS[31][8] ), .B(n3201), .S(n26), .Z(n1148) );
  AND2_X1 U3305 ( .A1(DATAIN[8]), .A2(n3212), .ZN(n3201) );
  MUX2_X1 U3306 ( .A(\REGISTERS[31][7] ), .B(n3202), .S(n26), .Z(n1147) );
  AND2_X1 U3307 ( .A1(DATAIN[7]), .A2(n3212), .ZN(n3202) );
  MUX2_X1 U3308 ( .A(\REGISTERS[31][6] ), .B(n3203), .S(n26), .Z(n1146) );
  AND2_X1 U3309 ( .A1(DATAIN[6]), .A2(n3212), .ZN(n3203) );
  MUX2_X1 U3310 ( .A(\REGISTERS[31][5] ), .B(n3204), .S(n26), .Z(n1145) );
  AND2_X1 U3311 ( .A1(DATAIN[5]), .A2(n3212), .ZN(n3204) );
  MUX2_X1 U3312 ( .A(\REGISTERS[31][4] ), .B(n3205), .S(n26), .Z(n1144) );
  AND2_X1 U3313 ( .A1(DATAIN[4]), .A2(n3212), .ZN(n3205) );
  MUX2_X1 U3314 ( .A(\REGISTERS[31][3] ), .B(n3206), .S(n26), .Z(n1143) );
  AND2_X1 U3315 ( .A1(DATAIN[3]), .A2(n3212), .ZN(n3206) );
  MUX2_X1 U3316 ( .A(\REGISTERS[31][2] ), .B(n3207), .S(n26), .Z(n1142) );
  AND2_X1 U3317 ( .A1(DATAIN[2]), .A2(n3212), .ZN(n3207) );
  MUX2_X1 U3318 ( .A(\REGISTERS[31][1] ), .B(n3208), .S(n26), .Z(n1141) );
  AND2_X1 U3319 ( .A1(DATAIN[1]), .A2(n3212), .ZN(n3208) );
  MUX2_X1 U3320 ( .A(\REGISTERS[31][0] ), .B(n3209), .S(n26), .Z(n1140) );
  OAI21_X1 U3321 ( .B1(n3226), .B2(n3249), .A(n3212), .ZN(n3259) );
  NAND3_X1 U3322 ( .A1(ADD_WR[3]), .A2(n3229), .A3(ADD_WR[4]), .ZN(n3249) );
  AND2_X1 U3323 ( .A1(WR), .A2(ENABLE), .ZN(n3229) );
  NAND3_X1 U3324 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n3226)
         );
  AND2_X1 U3325 ( .A1(DATAIN[0]), .A2(n3212), .ZN(n3209) );
  AND2_X1 U3326 ( .A1(RD2), .A2(ENABLE), .ZN(N445) );
  AND2_X1 U3327 ( .A1(RD1), .A2(ENABLE), .ZN(N444) );
endmodule


module ffd_234 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_233 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_232 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_231 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_230 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_229 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_228 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_227 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_226 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_225 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_224 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_223 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_222 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_221 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_220 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_219 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_218 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_217 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_216 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_215 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_214 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_213 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_212 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_211 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_210 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_209 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_208 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_207 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_206 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_205 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_204 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_203 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_7 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;
  wire   n1, n2, n3;

  ffd_234 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[31]) );
  ffd_233 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[30]) );
  ffd_232 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[29]) );
  ffd_231 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[28]) );
  ffd_230 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[27]) );
  ffd_229 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[26]) );
  ffd_228 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[25]) );
  ffd_227 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[24]) );
  ffd_226 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[23]) );
  ffd_225 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[22]) );
  ffd_224 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[21]) );
  ffd_223 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[20]) );
  ffd_222 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[19]) );
  ffd_221 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[18]) );
  ffd_220 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[17]) );
  ffd_219 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[16]) );
  ffd_218 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[15]) );
  ffd_217 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[14]) );
  ffd_216 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[13]) );
  ffd_215 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[12]) );
  ffd_214 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[11]) );
  ffd_213 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[10]) );
  ffd_212 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[9]) );
  ffd_211 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[8]) );
  ffd_210 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[7]) );
  ffd_209 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[6]) );
  ffd_208 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[5]) );
  ffd_207 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[4]) );
  ffd_206 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[3]) );
  ffd_205 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[2]) );
  ffd_204 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[1]) );
  ffd_203 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[0]) );
  BUF_X1 U1 ( .A(Enable), .Z(n1) );
  BUF_X1 U2 ( .A(Enable), .Z(n2) );
  BUF_X1 U3 ( .A(Enable), .Z(n3) );
endmodule


module ffd_202 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_201 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_200 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_199 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_198 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_197 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_196 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_195 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_194 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_193 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_192 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_191 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_190 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_189 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_188 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_187 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_186 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_185 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_184 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_183 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_182 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_181 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_180 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_179 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_178 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_177 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_176 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_175 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_174 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_173 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_172 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_171 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_6 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;
  wire   n1, n2, n3;

  ffd_202 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[31]) );
  ffd_201 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[30]) );
  ffd_200 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[29]) );
  ffd_199 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[28]) );
  ffd_198 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[27]) );
  ffd_197 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[26]) );
  ffd_196 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[25]) );
  ffd_195 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[24]) );
  ffd_194 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[23]) );
  ffd_193 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[22]) );
  ffd_192 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[21]) );
  ffd_191 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[20]) );
  ffd_190 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[19]) );
  ffd_189 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[18]) );
  ffd_188 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[17]) );
  ffd_187 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[16]) );
  ffd_186 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[15]) );
  ffd_185 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[14]) );
  ffd_184 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[13]) );
  ffd_183 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[12]) );
  ffd_182 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[11]) );
  ffd_181 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[10]) );
  ffd_180 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[9]) );
  ffd_179 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[8]) );
  ffd_178 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[7]) );
  ffd_177 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[6]) );
  ffd_176 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[5]) );
  ffd_175 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[4]) );
  ffd_174 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[3]) );
  ffd_173 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[2]) );
  ffd_172 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[1]) );
  ffd_171 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[0]) );
  BUF_X1 U1 ( .A(Enable), .Z(n1) );
  BUF_X1 U2 ( .A(Enable), .Z(n2) );
  BUF_X1 U3 ( .A(Enable), .Z(n3) );
endmodule


module ffd_170 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_169 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_168 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_167 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_166 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_165 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_164 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_163 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_162 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_161 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_160 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_159 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_158 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_157 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_156 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_155 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_154 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_153 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_152 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_151 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_150 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_149 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_148 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_147 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_146 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_145 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_144 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_143 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_142 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_141 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_140 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_139 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_5 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;
  wire   n1, n2, n3;

  ffd_170 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[31]) );
  ffd_169 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[30]) );
  ffd_168 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[29]) );
  ffd_167 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[28]) );
  ffd_166 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[27]) );
  ffd_165 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[26]) );
  ffd_164 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[25]) );
  ffd_163 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[24]) );
  ffd_162 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[23]) );
  ffd_161 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[22]) );
  ffd_160 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[21]) );
  ffd_159 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[20]) );
  ffd_158 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[19]) );
  ffd_157 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[18]) );
  ffd_156 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[17]) );
  ffd_155 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[16]) );
  ffd_154 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[15]) );
  ffd_153 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[14]) );
  ffd_152 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[13]) );
  ffd_151 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[12]) );
  ffd_150 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[11]) );
  ffd_149 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[10]) );
  ffd_148 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[9]) );
  ffd_147 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[8]) );
  ffd_146 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[7]) );
  ffd_145 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[6]) );
  ffd_144 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[5]) );
  ffd_143 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[4]) );
  ffd_142 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[3]) );
  ffd_141 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[2]) );
  ffd_140 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[1]) );
  ffd_139 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[0]) );
  BUF_X1 U1 ( .A(Enable), .Z(n1) );
  BUF_X1 U2 ( .A(Enable), .Z(n2) );
  BUF_X1 U3 ( .A(Enable), .Z(n3) );
endmodule


module ffd_138 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_137 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_136 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_135 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_134 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_133 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_132 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_131 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_130 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_129 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_128 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_127 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_126 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_125 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_124 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_123 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_122 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_121 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_120 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_119 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_118 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_117 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_116 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_115 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_114 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_113 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_112 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_111 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_110 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_109 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_108 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_107 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_4 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;
  wire   n1, n2, n3;

  ffd_138 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[31]) );
  ffd_137 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[30]) );
  ffd_136 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[29]) );
  ffd_135 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[28]) );
  ffd_134 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[27]) );
  ffd_133 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[26]) );
  ffd_132 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[25]) );
  ffd_131 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[24]) );
  ffd_130 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[23]) );
  ffd_129 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[22]) );
  ffd_128 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[21]) );
  ffd_127 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(n1), .Q(
        regOut[20]) );
  ffd_126 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[19]) );
  ffd_125 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[18]) );
  ffd_124 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[17]) );
  ffd_123 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[16]) );
  ffd_122 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[15]) );
  ffd_121 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[14]) );
  ffd_120 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[13]) );
  ffd_119 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[12]) );
  ffd_118 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[11]) );
  ffd_117 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(n2), .Q(
        regOut[10]) );
  ffd_116 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[9]) );
  ffd_115 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(n2), .Q(regOut[8]) );
  ffd_114 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[7]) );
  ffd_113 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[6]) );
  ffd_112 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[5]) );
  ffd_111 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[4]) );
  ffd_110 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[3]) );
  ffd_109 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[2]) );
  ffd_108 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[1]) );
  ffd_107 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(n3), .Q(regOut[0]) );
  BUF_X1 U1 ( .A(Enable), .Z(n1) );
  BUF_X1 U2 ( .A(Enable), .Z(n2) );
  BUF_X1 U3 ( .A(Enable), .Z(n3) );
endmodule


module ffd_106 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_105 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_104 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_103 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_102 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N5_0 ( regIn, Clk, Reset, Enable, regOut );
  input [4:0] regIn;
  output [4:0] regOut;
  input Clk, Reset, Enable;


  ffd_106 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_105 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_104 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_103 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_102 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module MUX41_GENERIC_N32_0 ( SHIFTER_OUT, ADD_OUT, CMP_OUT, LOGICALS_OUT, SEL, 
        Y );
  input [31:0] SHIFTER_OUT;
  input [31:0] ADD_OUT;
  input [31:0] CMP_OUT;
  input [31:0] LOGICALS_OUT;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;

  AND2_X2 U1 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n4) );
  AND2_X2 U2 ( .A1(SEL[1]), .A2(n69), .ZN(n3) );
  NOR2_X4 U3 ( .A1(n69), .A2(SEL[1]), .ZN(n6) );
  NOR2_X4 U4 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n1), .A2(n2), .ZN(Y[9]) );
  AOI22_X1 U6 ( .A1(CMP_OUT[9]), .A2(n3), .B1(LOGICALS_OUT[9]), .B2(n4), .ZN(
        n2) );
  AOI22_X1 U7 ( .A1(SHIFTER_OUT[9]), .A2(n5), .B1(ADD_OUT[9]), .B2(n6), .ZN(n1) );
  NAND2_X1 U8 ( .A1(n7), .A2(n8), .ZN(Y[8]) );
  AOI22_X1 U9 ( .A1(CMP_OUT[8]), .A2(n3), .B1(LOGICALS_OUT[8]), .B2(n4), .ZN(
        n8) );
  AOI22_X1 U10 ( .A1(SHIFTER_OUT[8]), .A2(n5), .B1(ADD_OUT[8]), .B2(n6), .ZN(
        n7) );
  NAND2_X1 U11 ( .A1(n9), .A2(n10), .ZN(Y[7]) );
  AOI22_X1 U12 ( .A1(CMP_OUT[7]), .A2(n3), .B1(LOGICALS_OUT[7]), .B2(n4), .ZN(
        n10) );
  AOI22_X1 U13 ( .A1(SHIFTER_OUT[7]), .A2(n5), .B1(ADD_OUT[7]), .B2(n6), .ZN(
        n9) );
  NAND2_X1 U14 ( .A1(n11), .A2(n12), .ZN(Y[6]) );
  AOI22_X1 U15 ( .A1(CMP_OUT[6]), .A2(n3), .B1(LOGICALS_OUT[6]), .B2(n4), .ZN(
        n12) );
  AOI22_X1 U16 ( .A1(SHIFTER_OUT[6]), .A2(n5), .B1(ADD_OUT[6]), .B2(n6), .ZN(
        n11) );
  NAND2_X1 U17 ( .A1(n13), .A2(n14), .ZN(Y[5]) );
  AOI22_X1 U18 ( .A1(CMP_OUT[5]), .A2(n3), .B1(LOGICALS_OUT[5]), .B2(n4), .ZN(
        n14) );
  AOI22_X1 U19 ( .A1(SHIFTER_OUT[5]), .A2(n5), .B1(ADD_OUT[5]), .B2(n6), .ZN(
        n13) );
  NAND2_X1 U20 ( .A1(n15), .A2(n16), .ZN(Y[4]) );
  AOI22_X1 U21 ( .A1(CMP_OUT[4]), .A2(n3), .B1(LOGICALS_OUT[4]), .B2(n4), .ZN(
        n16) );
  AOI22_X1 U22 ( .A1(SHIFTER_OUT[4]), .A2(n5), .B1(ADD_OUT[4]), .B2(n6), .ZN(
        n15) );
  NAND2_X1 U23 ( .A1(n17), .A2(n18), .ZN(Y[3]) );
  AOI22_X1 U24 ( .A1(CMP_OUT[3]), .A2(n3), .B1(LOGICALS_OUT[3]), .B2(n4), .ZN(
        n18) );
  AOI22_X1 U25 ( .A1(SHIFTER_OUT[3]), .A2(n5), .B1(ADD_OUT[3]), .B2(n6), .ZN(
        n17) );
  NAND2_X1 U26 ( .A1(n19), .A2(n20), .ZN(Y[31]) );
  AOI22_X1 U27 ( .A1(CMP_OUT[31]), .A2(n3), .B1(LOGICALS_OUT[31]), .B2(n4), 
        .ZN(n20) );
  AOI22_X1 U28 ( .A1(SHIFTER_OUT[31]), .A2(n5), .B1(ADD_OUT[31]), .B2(n6), 
        .ZN(n19) );
  NAND2_X1 U29 ( .A1(n21), .A2(n22), .ZN(Y[30]) );
  AOI22_X1 U30 ( .A1(CMP_OUT[30]), .A2(n3), .B1(LOGICALS_OUT[30]), .B2(n4), 
        .ZN(n22) );
  AOI22_X1 U31 ( .A1(SHIFTER_OUT[30]), .A2(n5), .B1(ADD_OUT[30]), .B2(n6), 
        .ZN(n21) );
  NAND2_X1 U32 ( .A1(n23), .A2(n24), .ZN(Y[2]) );
  AOI22_X1 U33 ( .A1(CMP_OUT[2]), .A2(n3), .B1(LOGICALS_OUT[2]), .B2(n4), .ZN(
        n24) );
  AOI22_X1 U34 ( .A1(SHIFTER_OUT[2]), .A2(n5), .B1(ADD_OUT[2]), .B2(n6), .ZN(
        n23) );
  NAND2_X1 U35 ( .A1(n25), .A2(n26), .ZN(Y[29]) );
  AOI22_X1 U36 ( .A1(CMP_OUT[29]), .A2(n3), .B1(LOGICALS_OUT[29]), .B2(n4), 
        .ZN(n26) );
  AOI22_X1 U37 ( .A1(SHIFTER_OUT[29]), .A2(n5), .B1(ADD_OUT[29]), .B2(n6), 
        .ZN(n25) );
  NAND2_X1 U38 ( .A1(n27), .A2(n28), .ZN(Y[28]) );
  AOI22_X1 U39 ( .A1(CMP_OUT[28]), .A2(n3), .B1(LOGICALS_OUT[28]), .B2(n4), 
        .ZN(n28) );
  AOI22_X1 U40 ( .A1(SHIFTER_OUT[28]), .A2(n5), .B1(ADD_OUT[28]), .B2(n6), 
        .ZN(n27) );
  NAND2_X1 U41 ( .A1(n29), .A2(n30), .ZN(Y[27]) );
  AOI22_X1 U42 ( .A1(CMP_OUT[27]), .A2(n3), .B1(LOGICALS_OUT[27]), .B2(n4), 
        .ZN(n30) );
  AOI22_X1 U43 ( .A1(SHIFTER_OUT[27]), .A2(n5), .B1(ADD_OUT[27]), .B2(n6), 
        .ZN(n29) );
  NAND2_X1 U44 ( .A1(n31), .A2(n32), .ZN(Y[26]) );
  AOI22_X1 U45 ( .A1(CMP_OUT[26]), .A2(n3), .B1(LOGICALS_OUT[26]), .B2(n4), 
        .ZN(n32) );
  AOI22_X1 U46 ( .A1(SHIFTER_OUT[26]), .A2(n5), .B1(ADD_OUT[26]), .B2(n6), 
        .ZN(n31) );
  NAND2_X1 U47 ( .A1(n33), .A2(n34), .ZN(Y[25]) );
  AOI22_X1 U48 ( .A1(CMP_OUT[25]), .A2(n3), .B1(LOGICALS_OUT[25]), .B2(n4), 
        .ZN(n34) );
  AOI22_X1 U49 ( .A1(SHIFTER_OUT[25]), .A2(n5), .B1(ADD_OUT[25]), .B2(n6), 
        .ZN(n33) );
  NAND2_X1 U50 ( .A1(n35), .A2(n36), .ZN(Y[24]) );
  AOI22_X1 U51 ( .A1(CMP_OUT[24]), .A2(n3), .B1(LOGICALS_OUT[24]), .B2(n4), 
        .ZN(n36) );
  AOI22_X1 U52 ( .A1(SHIFTER_OUT[24]), .A2(n5), .B1(ADD_OUT[24]), .B2(n6), 
        .ZN(n35) );
  NAND2_X1 U53 ( .A1(n37), .A2(n38), .ZN(Y[23]) );
  AOI22_X1 U54 ( .A1(CMP_OUT[23]), .A2(n3), .B1(LOGICALS_OUT[23]), .B2(n4), 
        .ZN(n38) );
  AOI22_X1 U55 ( .A1(SHIFTER_OUT[23]), .A2(n5), .B1(ADD_OUT[23]), .B2(n6), 
        .ZN(n37) );
  NAND2_X1 U56 ( .A1(n39), .A2(n40), .ZN(Y[22]) );
  AOI22_X1 U57 ( .A1(CMP_OUT[22]), .A2(n3), .B1(LOGICALS_OUT[22]), .B2(n4), 
        .ZN(n40) );
  AOI22_X1 U58 ( .A1(SHIFTER_OUT[22]), .A2(n5), .B1(ADD_OUT[22]), .B2(n6), 
        .ZN(n39) );
  NAND2_X1 U59 ( .A1(n41), .A2(n42), .ZN(Y[21]) );
  AOI22_X1 U60 ( .A1(CMP_OUT[21]), .A2(n3), .B1(LOGICALS_OUT[21]), .B2(n4), 
        .ZN(n42) );
  AOI22_X1 U61 ( .A1(SHIFTER_OUT[21]), .A2(n5), .B1(ADD_OUT[21]), .B2(n6), 
        .ZN(n41) );
  NAND2_X1 U62 ( .A1(n43), .A2(n44), .ZN(Y[20]) );
  AOI22_X1 U63 ( .A1(CMP_OUT[20]), .A2(n3), .B1(LOGICALS_OUT[20]), .B2(n4), 
        .ZN(n44) );
  AOI22_X1 U64 ( .A1(SHIFTER_OUT[20]), .A2(n5), .B1(ADD_OUT[20]), .B2(n6), 
        .ZN(n43) );
  NAND2_X1 U65 ( .A1(n45), .A2(n46), .ZN(Y[1]) );
  AOI22_X1 U66 ( .A1(CMP_OUT[1]), .A2(n3), .B1(LOGICALS_OUT[1]), .B2(n4), .ZN(
        n46) );
  AOI22_X1 U67 ( .A1(SHIFTER_OUT[1]), .A2(n5), .B1(ADD_OUT[1]), .B2(n6), .ZN(
        n45) );
  NAND2_X1 U68 ( .A1(n47), .A2(n48), .ZN(Y[19]) );
  AOI22_X1 U69 ( .A1(CMP_OUT[19]), .A2(n3), .B1(LOGICALS_OUT[19]), .B2(n4), 
        .ZN(n48) );
  AOI22_X1 U70 ( .A1(SHIFTER_OUT[19]), .A2(n5), .B1(ADD_OUT[19]), .B2(n6), 
        .ZN(n47) );
  NAND2_X1 U71 ( .A1(n49), .A2(n50), .ZN(Y[18]) );
  AOI22_X1 U72 ( .A1(CMP_OUT[18]), .A2(n3), .B1(LOGICALS_OUT[18]), .B2(n4), 
        .ZN(n50) );
  AOI22_X1 U73 ( .A1(SHIFTER_OUT[18]), .A2(n5), .B1(ADD_OUT[18]), .B2(n6), 
        .ZN(n49) );
  NAND2_X1 U74 ( .A1(n51), .A2(n52), .ZN(Y[17]) );
  AOI22_X1 U75 ( .A1(CMP_OUT[17]), .A2(n3), .B1(LOGICALS_OUT[17]), .B2(n4), 
        .ZN(n52) );
  AOI22_X1 U76 ( .A1(SHIFTER_OUT[17]), .A2(n5), .B1(ADD_OUT[17]), .B2(n6), 
        .ZN(n51) );
  NAND2_X1 U77 ( .A1(n53), .A2(n54), .ZN(Y[16]) );
  AOI22_X1 U78 ( .A1(CMP_OUT[16]), .A2(n3), .B1(LOGICALS_OUT[16]), .B2(n4), 
        .ZN(n54) );
  AOI22_X1 U79 ( .A1(SHIFTER_OUT[16]), .A2(n5), .B1(ADD_OUT[16]), .B2(n6), 
        .ZN(n53) );
  NAND2_X1 U80 ( .A1(n55), .A2(n56), .ZN(Y[15]) );
  AOI22_X1 U81 ( .A1(CMP_OUT[15]), .A2(n3), .B1(LOGICALS_OUT[15]), .B2(n4), 
        .ZN(n56) );
  AOI22_X1 U82 ( .A1(SHIFTER_OUT[15]), .A2(n5), .B1(ADD_OUT[15]), .B2(n6), 
        .ZN(n55) );
  NAND2_X1 U83 ( .A1(n57), .A2(n58), .ZN(Y[14]) );
  AOI22_X1 U84 ( .A1(CMP_OUT[14]), .A2(n3), .B1(LOGICALS_OUT[14]), .B2(n4), 
        .ZN(n58) );
  AOI22_X1 U85 ( .A1(SHIFTER_OUT[14]), .A2(n5), .B1(ADD_OUT[14]), .B2(n6), 
        .ZN(n57) );
  NAND2_X1 U86 ( .A1(n59), .A2(n60), .ZN(Y[13]) );
  AOI22_X1 U87 ( .A1(CMP_OUT[13]), .A2(n3), .B1(LOGICALS_OUT[13]), .B2(n4), 
        .ZN(n60) );
  AOI22_X1 U88 ( .A1(SHIFTER_OUT[13]), .A2(n5), .B1(ADD_OUT[13]), .B2(n6), 
        .ZN(n59) );
  NAND2_X1 U89 ( .A1(n61), .A2(n62), .ZN(Y[12]) );
  AOI22_X1 U90 ( .A1(CMP_OUT[12]), .A2(n3), .B1(LOGICALS_OUT[12]), .B2(n4), 
        .ZN(n62) );
  AOI22_X1 U91 ( .A1(SHIFTER_OUT[12]), .A2(n5), .B1(ADD_OUT[12]), .B2(n6), 
        .ZN(n61) );
  NAND2_X1 U92 ( .A1(n63), .A2(n64), .ZN(Y[11]) );
  AOI22_X1 U93 ( .A1(CMP_OUT[11]), .A2(n3), .B1(LOGICALS_OUT[11]), .B2(n4), 
        .ZN(n64) );
  AOI22_X1 U94 ( .A1(SHIFTER_OUT[11]), .A2(n5), .B1(ADD_OUT[11]), .B2(n6), 
        .ZN(n63) );
  NAND2_X1 U95 ( .A1(n65), .A2(n66), .ZN(Y[10]) );
  AOI22_X1 U96 ( .A1(CMP_OUT[10]), .A2(n3), .B1(LOGICALS_OUT[10]), .B2(n4), 
        .ZN(n66) );
  AOI22_X1 U97 ( .A1(SHIFTER_OUT[10]), .A2(n5), .B1(ADD_OUT[10]), .B2(n6), 
        .ZN(n65) );
  NAND2_X1 U98 ( .A1(n67), .A2(n68), .ZN(Y[0]) );
  AOI22_X1 U99 ( .A1(CMP_OUT[0]), .A2(n3), .B1(LOGICALS_OUT[0]), .B2(n4), .ZN(
        n68) );
  AOI22_X1 U100 ( .A1(SHIFTER_OUT[0]), .A2(n5), .B1(ADD_OUT[0]), .B2(n6), .ZN(
        n67) );
  INV_X1 U101 ( .A(SEL[0]), .ZN(n69) );
endmodule


module IR_decoder_N32 ( IR_IN, RS1, RS2, RD, imm16, imm26 );
  input [31:0] IR_IN;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [15:0] imm16;
  output [25:0] imm26;
  wire   \IR_IN[25] , \IR_IN[24] , \IR_IN[23] , \IR_IN[22] , \IR_IN[21] ,
         \IR_IN[20] , \IR_IN[19] , \IR_IN[18] , \IR_IN[17] , \IR_IN[16] ,
         \IR_IN[15] , \IR_IN[14] , \IR_IN[13] , \IR_IN[12] , \IR_IN[11] ,
         \IR_IN[10] , \IR_IN[9] , \IR_IN[8] , \IR_IN[7] , \IR_IN[6] ,
         \IR_IN[5] , \IR_IN[4] , \IR_IN[3] , \IR_IN[2] , \IR_IN[1] ,
         \IR_IN[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9;
  assign imm26[25] = \IR_IN[25] ;
  assign RS1[4] = \IR_IN[25] ;
  assign \IR_IN[25]  = IR_IN[25];
  assign imm26[24] = \IR_IN[24] ;
  assign RS1[3] = \IR_IN[24] ;
  assign \IR_IN[24]  = IR_IN[24];
  assign imm26[23] = \IR_IN[23] ;
  assign RS1[2] = \IR_IN[23] ;
  assign \IR_IN[23]  = IR_IN[23];
  assign imm26[22] = \IR_IN[22] ;
  assign RS1[1] = \IR_IN[22] ;
  assign \IR_IN[22]  = IR_IN[22];
  assign imm26[21] = \IR_IN[21] ;
  assign RS1[0] = \IR_IN[21] ;
  assign \IR_IN[21]  = IR_IN[21];
  assign imm26[20] = \IR_IN[20] ;
  assign RS2[4] = \IR_IN[20] ;
  assign \IR_IN[20]  = IR_IN[20];
  assign imm26[19] = \IR_IN[19] ;
  assign RS2[3] = \IR_IN[19] ;
  assign \IR_IN[19]  = IR_IN[19];
  assign imm26[18] = \IR_IN[18] ;
  assign RS2[2] = \IR_IN[18] ;
  assign \IR_IN[18]  = IR_IN[18];
  assign imm26[17] = \IR_IN[17] ;
  assign RS2[1] = \IR_IN[17] ;
  assign \IR_IN[17]  = IR_IN[17];
  assign imm26[16] = \IR_IN[16] ;
  assign RS2[0] = \IR_IN[16] ;
  assign \IR_IN[16]  = IR_IN[16];
  assign imm26[15] = \IR_IN[15] ;
  assign imm16[15] = \IR_IN[15] ;
  assign \IR_IN[15]  = IR_IN[15];
  assign imm26[14] = \IR_IN[14] ;
  assign imm16[14] = \IR_IN[14] ;
  assign \IR_IN[14]  = IR_IN[14];
  assign imm26[13] = \IR_IN[13] ;
  assign imm16[13] = \IR_IN[13] ;
  assign \IR_IN[13]  = IR_IN[13];
  assign imm26[12] = \IR_IN[12] ;
  assign imm16[12] = \IR_IN[12] ;
  assign \IR_IN[12]  = IR_IN[12];
  assign imm26[11] = \IR_IN[11] ;
  assign imm16[11] = \IR_IN[11] ;
  assign \IR_IN[11]  = IR_IN[11];
  assign imm26[10] = \IR_IN[10] ;
  assign imm16[10] = \IR_IN[10] ;
  assign \IR_IN[10]  = IR_IN[10];
  assign imm26[9] = \IR_IN[9] ;
  assign imm16[9] = \IR_IN[9] ;
  assign \IR_IN[9]  = IR_IN[9];
  assign imm26[8] = \IR_IN[8] ;
  assign imm16[8] = \IR_IN[8] ;
  assign \IR_IN[8]  = IR_IN[8];
  assign imm26[7] = \IR_IN[7] ;
  assign imm16[7] = \IR_IN[7] ;
  assign \IR_IN[7]  = IR_IN[7];
  assign imm26[6] = \IR_IN[6] ;
  assign imm16[6] = \IR_IN[6] ;
  assign \IR_IN[6]  = IR_IN[6];
  assign imm26[5] = \IR_IN[5] ;
  assign imm16[5] = \IR_IN[5] ;
  assign \IR_IN[5]  = IR_IN[5];
  assign imm26[4] = \IR_IN[4] ;
  assign imm16[4] = \IR_IN[4] ;
  assign \IR_IN[4]  = IR_IN[4];
  assign imm26[3] = \IR_IN[3] ;
  assign imm16[3] = \IR_IN[3] ;
  assign \IR_IN[3]  = IR_IN[3];
  assign imm26[2] = \IR_IN[2] ;
  assign imm16[2] = \IR_IN[2] ;
  assign \IR_IN[2]  = IR_IN[2];
  assign imm26[1] = \IR_IN[1] ;
  assign imm16[1] = \IR_IN[1] ;
  assign \IR_IN[1]  = IR_IN[1];
  assign imm26[0] = \IR_IN[0] ;
  assign imm16[0] = \IR_IN[0] ;
  assign \IR_IN[0]  = IR_IN[0];

  NOR4_X2 U2 ( .A1(IR_IN[26]), .A2(n8), .A3(IR_IN[30]), .A4(IR_IN[27]), .ZN(n3) );
  OR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(RD[4]) );
  MUX2_X1 U4 ( .A(\IR_IN[20] ), .B(\IR_IN[15] ), .S(n3), .Z(n2) );
  OR2_X1 U5 ( .A1(n1), .A2(n4), .ZN(RD[3]) );
  MUX2_X1 U6 ( .A(\IR_IN[19] ), .B(\IR_IN[14] ), .S(n3), .Z(n4) );
  OR2_X1 U7 ( .A1(n1), .A2(n5), .ZN(RD[2]) );
  MUX2_X1 U8 ( .A(\IR_IN[18] ), .B(\IR_IN[13] ), .S(n3), .Z(n5) );
  OR2_X1 U9 ( .A1(n1), .A2(n6), .ZN(RD[1]) );
  MUX2_X1 U10 ( .A(\IR_IN[17] ), .B(\IR_IN[12] ), .S(n3), .Z(n6) );
  OR2_X1 U11 ( .A1(n1), .A2(n7), .ZN(RD[0]) );
  MUX2_X1 U12 ( .A(\IR_IN[16] ), .B(\IR_IN[11] ), .S(n3), .Z(n7) );
  INV_X1 U13 ( .A(n9), .ZN(n8) );
  AND3_X1 U14 ( .A1(IR_IN[26]), .A2(n9), .A3(IR_IN[27]), .ZN(n1) );
  NOR3_X1 U15 ( .A1(IR_IN[31]), .A2(IR_IN[29]), .A3(IR_IN[28]), .ZN(n9) );
endmodule


module DU_N32 ( IR_IN, NPC, WR_ADDR_RF, DATAIN, EN1, RF1, RF2, WF1, CLK, RST, 
        SEL_IMM, NPC1_OUT, regA_OUT, regB_OUT, IMM_OUT, RD1_IN, RD1_OUT );
  input [31:0] IR_IN;
  input [31:0] NPC;
  input [4:0] WR_ADDR_RF;
  input [31:0] DATAIN;
  input [1:0] SEL_IMM;
  output [31:0] NPC1_OUT;
  output [31:0] regA_OUT;
  output [31:0] regB_OUT;
  output [31:0] IMM_OUT;
  output [4:0] RD1_IN;
  output [4:0] RD1_OUT;
  input EN1, RF1, RF2, WF1, CLK, RST;
  wire   imm1632_31, imm2632_31;
  wire   [14:0] imm1632;
  wire   [24:0] imm2632;
  wire   [4:0] RS1s;
  wire   [4:0] RS2s;
  wire   [31:0] registerA;
  wire   [31:0] registerB;
  wire   [31:0] immediate32;

  register_file_WORD_SIZE32_ADDR_SIZE5 RegisterFile ( .CLK(CLK), .RESET(RST), 
        .ENABLE(EN1), .RD1(RF1), .RD2(RF2), .WR(WF1), .ADD_WR(WR_ADDR_RF), 
        .ADD_RD1(RS1s), .ADD_RD2(RS2s), .DATAIN(DATAIN), .OUT1(registerA), 
        .OUT2(registerB) );
  regN_N32_7 NPC1reg ( .regIn(NPC), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(NPC1_OUT) );
  regN_N32_6 Areg ( .regIn(registerA), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(regA_OUT) );
  regN_N32_5 Breg ( .regIn(registerB), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(regB_OUT) );
  regN_N32_4 IMMreg ( .regIn(immediate32), .Clk(CLK), .Reset(RST), .Enable(EN1), .regOut(IMM_OUT) );
  regN_N5_0 RD1reg ( .regIn(RD1_IN), .Clk(CLK), .Reset(RST), .Enable(EN1), 
        .regOut(RD1_OUT) );
  MUX41_GENERIC_N32_0 MUXimm ( .SHIFTER_OUT({imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, imm1632_31, 
        imm1632_31, imm1632_31, imm1632_31, imm1632}), .ADD_OUT({imm2632_31, 
        imm2632_31, imm2632_31, imm2632_31, imm2632_31, imm2632_31, imm2632_31, 
        imm2632}), .CMP_OUT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, imm1632_31, imm1632}), 
        .LOGICALS_OUT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, imm2632_31, imm2632}), .SEL(SEL_IMM), .Y(immediate32) );
  IR_decoder_N32 DEC ( .IR_IN(IR_IN), .RS1(RS1s), .RS2(RS2s), .RD(RD1_IN), 
        .imm16({imm1632_31, imm1632}), .imm26({imm2632_31, imm2632}) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_160 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_159 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_158 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_157 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_156 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_155 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_154 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_153 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_152 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_151 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_150 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_149 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_148 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_147 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_146 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_145 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_144 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_143 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_142 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_141 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_140 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_139 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_138 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_137 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_136 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_135 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_134 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_133 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_132 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_131 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_130 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_129 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_128 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_127 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_126 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_125 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_124 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_123 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_122 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_121 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_120 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_119 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_118 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_117 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_116 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_115 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_114 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_113 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_112 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_111 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_110 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_109 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_108 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_107 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_106 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_105 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_104 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_103 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_102 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_101 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_100 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_99 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_98 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_97 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module XNOR2_0 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_31 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_30 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_29 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_28 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_27 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_26 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_25 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_24 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_23 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_22 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_21 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_20 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_19 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_18 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_17 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_16 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_15 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_14 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_13 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_12 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_11 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_10 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_9 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_8 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_7 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_6 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_5 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_4 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_3 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_2 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR2_1 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module AND2_0 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_45 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_44 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_43 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_42 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_41 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_40 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_39 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_38 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_37 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_36 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_35 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_34 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_33 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_32 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_31 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_30 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_29 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_28 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_27 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_26 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_25 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_24 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_23 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_22 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_21 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_20 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_19 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_18 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_17 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_16 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ZERODET_N32 ( A, Y );
  input [31:0] A;
  output Y;
  wire   \M[4][1] , \M[4][0] , \M[3][3] , \M[3][2] , \M[3][1] , \M[3][0] ,
         \M[2][7] , \M[2][6] , \M[2][5] , \M[2][4] , \M[2][3] , \M[2][2] ,
         \M[2][1] , \M[2][0] , \M[1][15] , \M[1][14] , \M[1][13] , \M[1][12] ,
         \M[1][11] , \M[1][10] , \M[1][9] , \M[1][8] , \M[1][7] , \M[1][6] ,
         \M[1][5] , \M[1][4] , \M[1][3] , \M[1][2] , \M[1][1] , \M[1][0] ,
         \M[0][31] , \M[0][30] , \M[0][29] , \M[0][28] , \M[0][27] ,
         \M[0][26] , \M[0][25] , \M[0][24] , \M[0][23] , \M[0][22] ,
         \M[0][21] , \M[0][20] , \M[0][19] , \M[0][18] , \M[0][17] ,
         \M[0][16] , \M[0][15] , \M[0][14] , \M[0][13] , \M[0][12] ,
         \M[0][11] , \M[0][10] , \M[0][9] , \M[0][8] , \M[0][7] , \M[0][6] ,
         \M[0][5] , \M[0][4] , \M[0][3] , \M[0][2] , \M[0][1] , \M[0][0] ;

  XNOR2_0 XOR0i_0_0 ( .A(A[0]), .B(1'b0), .Y(\M[0][0] ) );
  XNOR2_31 XOR0i_0_1 ( .A(A[1]), .B(1'b0), .Y(\M[0][1] ) );
  XNOR2_30 XOR0i_0_2 ( .A(A[2]), .B(1'b0), .Y(\M[0][2] ) );
  XNOR2_29 XOR0i_0_3 ( .A(A[3]), .B(1'b0), .Y(\M[0][3] ) );
  XNOR2_28 XOR0i_0_4 ( .A(A[4]), .B(1'b0), .Y(\M[0][4] ) );
  XNOR2_27 XOR0i_0_5 ( .A(A[5]), .B(1'b0), .Y(\M[0][5] ) );
  XNOR2_26 XOR0i_0_6 ( .A(A[6]), .B(1'b0), .Y(\M[0][6] ) );
  XNOR2_25 XOR0i_0_7 ( .A(A[7]), .B(1'b0), .Y(\M[0][7] ) );
  XNOR2_24 XOR0i_0_8 ( .A(A[8]), .B(1'b0), .Y(\M[0][8] ) );
  XNOR2_23 XOR0i_0_9 ( .A(A[9]), .B(1'b0), .Y(\M[0][9] ) );
  XNOR2_22 XOR0i_0_10 ( .A(A[10]), .B(1'b0), .Y(\M[0][10] ) );
  XNOR2_21 XOR0i_0_11 ( .A(A[11]), .B(1'b0), .Y(\M[0][11] ) );
  XNOR2_20 XOR0i_0_12 ( .A(A[12]), .B(1'b0), .Y(\M[0][12] ) );
  XNOR2_19 XOR0i_0_13 ( .A(A[13]), .B(1'b0), .Y(\M[0][13] ) );
  XNOR2_18 XOR0i_0_14 ( .A(A[14]), .B(1'b0), .Y(\M[0][14] ) );
  XNOR2_17 XOR0i_0_15 ( .A(A[15]), .B(1'b0), .Y(\M[0][15] ) );
  XNOR2_16 XOR0i_0_16 ( .A(A[16]), .B(1'b0), .Y(\M[0][16] ) );
  XNOR2_15 XOR0i_0_17 ( .A(A[17]), .B(1'b0), .Y(\M[0][17] ) );
  XNOR2_14 XOR0i_0_18 ( .A(A[18]), .B(1'b0), .Y(\M[0][18] ) );
  XNOR2_13 XOR0i_0_19 ( .A(A[19]), .B(1'b0), .Y(\M[0][19] ) );
  XNOR2_12 XOR0i_0_20 ( .A(A[20]), .B(1'b0), .Y(\M[0][20] ) );
  XNOR2_11 XOR0i_0_21 ( .A(A[21]), .B(1'b0), .Y(\M[0][21] ) );
  XNOR2_10 XOR0i_0_22 ( .A(A[22]), .B(1'b0), .Y(\M[0][22] ) );
  XNOR2_9 XOR0i_0_23 ( .A(A[23]), .B(1'b0), .Y(\M[0][23] ) );
  XNOR2_8 XOR0i_0_24 ( .A(A[24]), .B(1'b0), .Y(\M[0][24] ) );
  XNOR2_7 XOR0i_0_25 ( .A(A[25]), .B(1'b0), .Y(\M[0][25] ) );
  XNOR2_6 XOR0i_0_26 ( .A(A[26]), .B(1'b0), .Y(\M[0][26] ) );
  XNOR2_5 XOR0i_0_27 ( .A(A[27]), .B(1'b0), .Y(\M[0][27] ) );
  XNOR2_4 XOR0i_0_28 ( .A(A[28]), .B(1'b0), .Y(\M[0][28] ) );
  XNOR2_3 XOR0i_0_29 ( .A(A[29]), .B(1'b0), .Y(\M[0][29] ) );
  XNOR2_2 XOR0i_0_30 ( .A(A[30]), .B(1'b0), .Y(\M[0][30] ) );
  XNOR2_1 XOR0i_0_31 ( .A(A[31]), .B(1'b0), .Y(\M[0][31] ) );
  AND2_0 ANDi_1_0 ( .A(\M[0][0] ), .B(\M[0][1] ), .Y(\M[1][0] ) );
  AND2_45 ANDi_1_1 ( .A(\M[0][2] ), .B(\M[0][3] ), .Y(\M[1][1] ) );
  AND2_44 ANDi_1_2 ( .A(\M[0][4] ), .B(\M[0][5] ), .Y(\M[1][2] ) );
  AND2_43 ANDi_1_3 ( .A(\M[0][6] ), .B(\M[0][7] ), .Y(\M[1][3] ) );
  AND2_42 ANDi_1_4 ( .A(\M[0][8] ), .B(\M[0][9] ), .Y(\M[1][4] ) );
  AND2_41 ANDi_1_5 ( .A(\M[0][10] ), .B(\M[0][11] ), .Y(\M[1][5] ) );
  AND2_40 ANDi_1_6 ( .A(\M[0][12] ), .B(\M[0][13] ), .Y(\M[1][6] ) );
  AND2_39 ANDi_1_7 ( .A(\M[0][14] ), .B(\M[0][15] ), .Y(\M[1][7] ) );
  AND2_38 ANDi_1_8 ( .A(\M[0][16] ), .B(\M[0][17] ), .Y(\M[1][8] ) );
  AND2_37 ANDi_1_9 ( .A(\M[0][18] ), .B(\M[0][19] ), .Y(\M[1][9] ) );
  AND2_36 ANDi_1_10 ( .A(\M[0][20] ), .B(\M[0][21] ), .Y(\M[1][10] ) );
  AND2_35 ANDi_1_11 ( .A(\M[0][22] ), .B(\M[0][23] ), .Y(\M[1][11] ) );
  AND2_34 ANDi_1_12 ( .A(\M[0][24] ), .B(\M[0][25] ), .Y(\M[1][12] ) );
  AND2_33 ANDi_1_13 ( .A(\M[0][26] ), .B(\M[0][27] ), .Y(\M[1][13] ) );
  AND2_32 ANDi_1_14 ( .A(\M[0][28] ), .B(\M[0][29] ), .Y(\M[1][14] ) );
  AND2_31 ANDi_1_15 ( .A(\M[0][30] ), .B(\M[0][31] ), .Y(\M[1][15] ) );
  AND2_30 ANDi_2_0 ( .A(\M[1][0] ), .B(\M[1][1] ), .Y(\M[2][0] ) );
  AND2_29 ANDi_2_1 ( .A(\M[1][2] ), .B(\M[1][3] ), .Y(\M[2][1] ) );
  AND2_28 ANDi_2_2 ( .A(\M[1][4] ), .B(\M[1][5] ), .Y(\M[2][2] ) );
  AND2_27 ANDi_2_3 ( .A(\M[1][6] ), .B(\M[1][7] ), .Y(\M[2][3] ) );
  AND2_26 ANDi_2_4 ( .A(\M[1][8] ), .B(\M[1][9] ), .Y(\M[2][4] ) );
  AND2_25 ANDi_2_5 ( .A(\M[1][10] ), .B(\M[1][11] ), .Y(\M[2][5] ) );
  AND2_24 ANDi_2_6 ( .A(\M[1][12] ), .B(\M[1][13] ), .Y(\M[2][6] ) );
  AND2_23 ANDi_2_7 ( .A(\M[1][14] ), .B(\M[1][15] ), .Y(\M[2][7] ) );
  AND2_22 ANDi_3_0 ( .A(\M[2][0] ), .B(\M[2][1] ), .Y(\M[3][0] ) );
  AND2_21 ANDi_3_1 ( .A(\M[2][2] ), .B(\M[2][3] ), .Y(\M[3][1] ) );
  AND2_20 ANDi_3_2 ( .A(\M[2][4] ), .B(\M[2][5] ), .Y(\M[3][2] ) );
  AND2_19 ANDi_3_3 ( .A(\M[2][6] ), .B(\M[2][7] ), .Y(\M[3][3] ) );
  AND2_18 ANDi_4_0 ( .A(\M[3][0] ), .B(\M[3][1] ), .Y(\M[4][0] ) );
  AND2_17 ANDi_4_1 ( .A(\M[3][2] ), .B(\M[3][3] ), .Y(\M[4][1] ) );
  AND2_16 ANDi_5_0 ( .A(\M[4][0] ), .B(\M[4][1] ), .Y(Y) );
endmodule


module MUX4_1 ( ZERO, ONE, INV_CMP, CMP, Sel, Y );
  input [1:0] Sel;
  input ZERO, ONE, INV_CMP, CMP;
  output Y;
  wire   n4, n2, n3;

  CLKBUF_X3 U1 ( .A(n4), .Z(Y) );
  MUX2_X1 U2 ( .A(n2), .B(n3), .S(Sel[1]), .Z(n4) );
  MUX2_X1 U3 ( .A(INV_CMP), .B(CMP), .S(Sel[0]), .Z(n3) );
  MUX2_X1 U4 ( .A(ZERO), .B(ONE), .S(Sel[0]), .Z(n2) );
endmodule


module ffd_101 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_100 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_99 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_98 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_97 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_96 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_95 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_94 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_93 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_92 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_91 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_90 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_89 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_88 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_87 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_86 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_85 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_84 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_83 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_82 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_81 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_80 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_79 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_78 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_77 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_76 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_75 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_74 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_73 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_72 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_71 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_70 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_3 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_101 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_100 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_99 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_98 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_97 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_96 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_95 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_94 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_93 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_92 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_91 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_90 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_89 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_88 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_87 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_86 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_85 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_84 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_83 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_82 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_81 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_80 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_79 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_78 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_77 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_76 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_75 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_74 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_73 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_72 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_71 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_70 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module xorGrid_N32 ( B, Cin, Bx );
  input [31:0] B;
  output [31:0] Bx;
  input Cin;


  XOR2_X1 U1 ( .A(Cin), .B(B[9]), .Z(Bx[9]) );
  XOR2_X1 U2 ( .A(Cin), .B(B[8]), .Z(Bx[8]) );
  XOR2_X1 U3 ( .A(Cin), .B(B[7]), .Z(Bx[7]) );
  XOR2_X1 U4 ( .A(Cin), .B(B[6]), .Z(Bx[6]) );
  XOR2_X1 U5 ( .A(Cin), .B(B[5]), .Z(Bx[5]) );
  XOR2_X1 U6 ( .A(Cin), .B(B[4]), .Z(Bx[4]) );
  XOR2_X1 U7 ( .A(Cin), .B(B[3]), .Z(Bx[3]) );
  XOR2_X1 U8 ( .A(Cin), .B(B[31]), .Z(Bx[31]) );
  XOR2_X1 U9 ( .A(Cin), .B(B[30]), .Z(Bx[30]) );
  XOR2_X1 U10 ( .A(Cin), .B(B[2]), .Z(Bx[2]) );
  XOR2_X1 U11 ( .A(Cin), .B(B[29]), .Z(Bx[29]) );
  XOR2_X1 U12 ( .A(Cin), .B(B[28]), .Z(Bx[28]) );
  XOR2_X1 U13 ( .A(Cin), .B(B[27]), .Z(Bx[27]) );
  XOR2_X1 U14 ( .A(Cin), .B(B[26]), .Z(Bx[26]) );
  XOR2_X1 U15 ( .A(Cin), .B(B[25]), .Z(Bx[25]) );
  XOR2_X1 U16 ( .A(Cin), .B(B[24]), .Z(Bx[24]) );
  XOR2_X1 U17 ( .A(Cin), .B(B[23]), .Z(Bx[23]) );
  XOR2_X1 U18 ( .A(Cin), .B(B[22]), .Z(Bx[22]) );
  XOR2_X1 U19 ( .A(Cin), .B(B[21]), .Z(Bx[21]) );
  XOR2_X1 U20 ( .A(Cin), .B(B[20]), .Z(Bx[20]) );
  XOR2_X1 U21 ( .A(Cin), .B(B[1]), .Z(Bx[1]) );
  XOR2_X1 U22 ( .A(Cin), .B(B[19]), .Z(Bx[19]) );
  XOR2_X1 U23 ( .A(Cin), .B(B[18]), .Z(Bx[18]) );
  XOR2_X1 U24 ( .A(Cin), .B(B[17]), .Z(Bx[17]) );
  XOR2_X1 U25 ( .A(Cin), .B(B[16]), .Z(Bx[16]) );
  XOR2_X1 U26 ( .A(Cin), .B(B[15]), .Z(Bx[15]) );
  XOR2_X1 U27 ( .A(Cin), .B(B[14]), .Z(Bx[14]) );
  XOR2_X1 U28 ( .A(Cin), .B(B[13]), .Z(Bx[13]) );
  XOR2_X1 U29 ( .A(Cin), .B(B[12]), .Z(Bx[12]) );
  XOR2_X1 U30 ( .A(Cin), .B(B[11]), .Z(Bx[11]) );
  XOR2_X1 U31 ( .A(Cin), .B(B[10]), .Z(Bx[10]) );
  XOR2_X1 U32 ( .A(Cin), .B(B[0]), .Z(Bx[0]) );
endmodule


module PG_NET_0 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_30 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_29 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_28 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_27 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_26 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_25 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_24 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_23 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_22 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_21 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_20 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_19 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_18 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_17 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_16 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_15 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_14 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_13 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_12 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_11 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_10 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_9 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_8 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_7 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_6 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_5 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_4 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_3 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_2 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_NET_1 ( A, B, P, G );
  input A, B;
  output P, G;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module G_BLOCK_0 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module PG_BLOCK_0 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_26 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_25 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_24 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_23 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_22 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_21 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_20 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_19 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_18 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_17 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_16 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_15 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_14 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_13 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module G_BLOCK_8 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module PG_BLOCK_12 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_11 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_10 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_9 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_8 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_7 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_6 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module G_BLOCK_7 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module PG_BLOCK_5 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_4 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_3 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module G_BLOCK_6 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module G_BLOCK_5 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module PG_BLOCK_2 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module PG_BLOCK_1 ( PIK, GIK, PK1J, GK1J, GIJ, PIJ );
  input PIK, GIK, PK1J, GK1J;
  output GIJ, PIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
  AND2_X1 U3 ( .A1(PK1J), .A2(PIK), .ZN(PIJ) );
endmodule


module G_BLOCK_4 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module G_BLOCK_3 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module G_BLOCK_2 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module G_BLOCK_1 ( PIK, GIK, GK1J, GIJ );
  input PIK, GIK, GK1J;
  output GIJ;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(GIJ) );
  AOI21_X1 U2 ( .B1(PIK), .B2(GK1J), .A(GIK), .ZN(n1) );
endmodule


module CARRY_GENERATOR_NBIT32_NBLOCK4 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Co;
  input Cin;
  wire   Cin, \PGNET_G[4][31] , \PGNET_G[4][27] , \PGNET_G[3][31] ,
         \PGNET_G[3][23] , \PGNET_G[3][15] , \PGNET_G[2][31] ,
         \PGNET_G[2][27] , \PGNET_G[2][23] , \PGNET_G[2][19] ,
         \PGNET_G[2][15] , \PGNET_G[2][11] , \PGNET_G[2][7] , \PGNET_G[1][31] ,
         \PGNET_G[1][29] , \PGNET_G[1][27] , \PGNET_G[1][25] ,
         \PGNET_G[1][23] , \PGNET_G[1][21] , \PGNET_G[1][19] ,
         \PGNET_G[1][17] , \PGNET_G[1][15] , \PGNET_G[1][13] ,
         \PGNET_G[1][11] , \PGNET_G[1][9] , \PGNET_G[1][7] , \PGNET_G[1][5] ,
         \PGNET_G[1][3] , \PGNET_G[1][1] , \PGNET_G[0][31] , \PGNET_G[0][30] ,
         \PGNET_G[0][29] , \PGNET_G[0][28] , \PGNET_G[0][27] ,
         \PGNET_G[0][26] , \PGNET_G[0][25] , \PGNET_G[0][24] ,
         \PGNET_G[0][23] , \PGNET_G[0][22] , \PGNET_G[0][21] ,
         \PGNET_G[0][20] , \PGNET_G[0][19] , \PGNET_G[0][18] ,
         \PGNET_G[0][17] , \PGNET_G[0][16] , \PGNET_G[0][15] ,
         \PGNET_G[0][14] , \PGNET_G[0][13] , \PGNET_G[0][12] ,
         \PGNET_G[0][11] , \PGNET_G[0][10] , \PGNET_G[0][9] , \PGNET_G[0][8] ,
         \PGNET_G[0][7] , \PGNET_G[0][6] , \PGNET_G[0][5] , \PGNET_G[0][4] ,
         \PGNET_G[0][3] , \PGNET_G[0][2] , \PGNET_G[0][1] , \PGNET_G[0][0] ,
         \PGNET_P[4][31] , \PGNET_P[4][27] , \PGNET_P[3][31] ,
         \PGNET_P[3][23] , \PGNET_P[3][15] , \PGNET_P[3][11] ,
         \PGNET_P[2][31] , \PGNET_P[2][27] , \PGNET_P[2][23] ,
         \PGNET_P[2][19] , \PGNET_P[2][15] , \PGNET_P[2][7] , \PGNET_P[1][31] ,
         \PGNET_P[1][29] , \PGNET_P[1][27] , \PGNET_P[1][25] ,
         \PGNET_P[1][23] , \PGNET_P[1][21] , \PGNET_P[1][19] ,
         \PGNET_P[1][17] , \PGNET_P[1][15] , \PGNET_P[1][13] ,
         \PGNET_P[1][11] , \PGNET_P[1][9] , \PGNET_P[1][7] , \PGNET_P[1][5] ,
         \PGNET_P[1][3] , \PGNET_P[0][31] , \PGNET_P[0][30] , \PGNET_P[0][29] ,
         \PGNET_P[0][28] , \PGNET_P[0][27] , \PGNET_P[0][26] ,
         \PGNET_P[0][25] , \PGNET_P[0][24] , \PGNET_P[0][23] ,
         \PGNET_P[0][22] , \PGNET_P[0][21] , \PGNET_P[0][20] ,
         \PGNET_P[0][19] , \PGNET_P[0][18] , \PGNET_P[0][17] ,
         \PGNET_P[0][16] , \PGNET_P[0][15] , \PGNET_P[0][14] ,
         \PGNET_P[0][13] , \PGNET_P[0][12] , \PGNET_P[0][11] ,
         \PGNET_P[0][10] , \PGNET_P[0][9] , \PGNET_P[0][8] , \PGNET_P[0][7] ,
         \PGNET_P[0][6] , \PGNET_P[0][5] , \PGNET_P[0][4] , \PGNET_P[0][3] ,
         \PGNET_P[0][2] , \PGNET_P[0][1] , n1, n2, n3;
  assign Co[0] = Cin;

  PG_NET_0 pgport_1 ( .A(A[1]), .B(B[1]), .P(\PGNET_P[0][1] ), .G(
        \PGNET_G[0][1] ) );
  PG_NET_30 pgport_2 ( .A(A[2]), .B(B[2]), .P(\PGNET_P[0][2] ), .G(
        \PGNET_G[0][2] ) );
  PG_NET_29 pgport_3 ( .A(A[3]), .B(B[3]), .P(\PGNET_P[0][3] ), .G(
        \PGNET_G[0][3] ) );
  PG_NET_28 pgport_4 ( .A(A[4]), .B(B[4]), .P(\PGNET_P[0][4] ), .G(
        \PGNET_G[0][4] ) );
  PG_NET_27 pgport_5 ( .A(A[5]), .B(B[5]), .P(\PGNET_P[0][5] ), .G(
        \PGNET_G[0][5] ) );
  PG_NET_26 pgport_6 ( .A(A[6]), .B(B[6]), .P(\PGNET_P[0][6] ), .G(
        \PGNET_G[0][6] ) );
  PG_NET_25 pgport_7 ( .A(A[7]), .B(B[7]), .P(\PGNET_P[0][7] ), .G(
        \PGNET_G[0][7] ) );
  PG_NET_24 pgport_8 ( .A(A[8]), .B(B[8]), .P(\PGNET_P[0][8] ), .G(
        \PGNET_G[0][8] ) );
  PG_NET_23 pgport_9 ( .A(A[9]), .B(B[9]), .P(\PGNET_P[0][9] ), .G(
        \PGNET_G[0][9] ) );
  PG_NET_22 pgport_10 ( .A(A[10]), .B(B[10]), .P(\PGNET_P[0][10] ), .G(
        \PGNET_G[0][10] ) );
  PG_NET_21 pgport_11 ( .A(A[11]), .B(B[11]), .P(\PGNET_P[0][11] ), .G(
        \PGNET_G[0][11] ) );
  PG_NET_20 pgport_12 ( .A(A[12]), .B(B[12]), .P(\PGNET_P[0][12] ), .G(
        \PGNET_G[0][12] ) );
  PG_NET_19 pgport_13 ( .A(A[13]), .B(B[13]), .P(\PGNET_P[0][13] ), .G(
        \PGNET_G[0][13] ) );
  PG_NET_18 pgport_14 ( .A(A[14]), .B(B[14]), .P(\PGNET_P[0][14] ), .G(
        \PGNET_G[0][14] ) );
  PG_NET_17 pgport_15 ( .A(A[15]), .B(B[15]), .P(\PGNET_P[0][15] ), .G(
        \PGNET_G[0][15] ) );
  PG_NET_16 pgport_16 ( .A(A[16]), .B(B[16]), .P(\PGNET_P[0][16] ), .G(
        \PGNET_G[0][16] ) );
  PG_NET_15 pgport_17 ( .A(A[17]), .B(B[17]), .P(\PGNET_P[0][17] ), .G(
        \PGNET_G[0][17] ) );
  PG_NET_14 pgport_18 ( .A(A[18]), .B(B[18]), .P(\PGNET_P[0][18] ), .G(
        \PGNET_G[0][18] ) );
  PG_NET_13 pgport_19 ( .A(A[19]), .B(B[19]), .P(\PGNET_P[0][19] ), .G(
        \PGNET_G[0][19] ) );
  PG_NET_12 pgport_20 ( .A(A[20]), .B(B[20]), .P(\PGNET_P[0][20] ), .G(
        \PGNET_G[0][20] ) );
  PG_NET_11 pgport_21 ( .A(A[21]), .B(B[21]), .P(\PGNET_P[0][21] ), .G(
        \PGNET_G[0][21] ) );
  PG_NET_10 pgport_22 ( .A(A[22]), .B(B[22]), .P(\PGNET_P[0][22] ), .G(
        \PGNET_G[0][22] ) );
  PG_NET_9 pgport_23 ( .A(A[23]), .B(B[23]), .P(\PGNET_P[0][23] ), .G(
        \PGNET_G[0][23] ) );
  PG_NET_8 pgport_24 ( .A(A[24]), .B(B[24]), .P(\PGNET_P[0][24] ), .G(
        \PGNET_G[0][24] ) );
  PG_NET_7 pgport_25 ( .A(A[25]), .B(B[25]), .P(\PGNET_P[0][25] ), .G(
        \PGNET_G[0][25] ) );
  PG_NET_6 pgport_26 ( .A(A[26]), .B(B[26]), .P(\PGNET_P[0][26] ), .G(
        \PGNET_G[0][26] ) );
  PG_NET_5 pgport_27 ( .A(A[27]), .B(B[27]), .P(\PGNET_P[0][27] ), .G(
        \PGNET_G[0][27] ) );
  PG_NET_4 pgport_28 ( .A(A[28]), .B(B[28]), .P(\PGNET_P[0][28] ), .G(
        \PGNET_G[0][28] ) );
  PG_NET_3 pgport_29 ( .A(A[29]), .B(B[29]), .P(\PGNET_P[0][29] ), .G(
        \PGNET_G[0][29] ) );
  PG_NET_2 pgport_30 ( .A(A[30]), .B(B[30]), .P(\PGNET_P[0][30] ), .G(
        \PGNET_G[0][30] ) );
  PG_NET_1 pgport_31 ( .A(A[31]), .B(B[31]), .P(\PGNET_P[0][31] ), .G(
        \PGNET_G[0][31] ) );
  G_BLOCK_0 gi_1_1 ( .PIK(\PGNET_P[0][1] ), .GIK(\PGNET_G[0][1] ), .GK1J(
        \PGNET_G[0][0] ), .GIJ(\PGNET_G[1][1] ) );
  PG_BLOCK_0 pgi_1_3 ( .PIK(\PGNET_P[0][3] ), .GIK(\PGNET_G[0][3] ), .PK1J(
        \PGNET_P[0][2] ), .GK1J(\PGNET_G[0][2] ), .GIJ(\PGNET_G[1][3] ), .PIJ(
        \PGNET_P[1][3] ) );
  PG_BLOCK_26 pgi_1_5 ( .PIK(\PGNET_P[0][5] ), .GIK(\PGNET_G[0][5] ), .PK1J(
        \PGNET_P[0][4] ), .GK1J(\PGNET_G[0][4] ), .GIJ(\PGNET_G[1][5] ), .PIJ(
        \PGNET_P[1][5] ) );
  PG_BLOCK_25 pgi_1_7 ( .PIK(\PGNET_P[0][7] ), .GIK(\PGNET_G[0][7] ), .PK1J(
        \PGNET_P[0][6] ), .GK1J(\PGNET_G[0][6] ), .GIJ(\PGNET_G[1][7] ), .PIJ(
        \PGNET_P[1][7] ) );
  PG_BLOCK_24 pgi_1_9 ( .PIK(\PGNET_P[0][9] ), .GIK(\PGNET_G[0][9] ), .PK1J(
        \PGNET_P[0][8] ), .GK1J(\PGNET_G[0][8] ), .GIJ(\PGNET_G[1][9] ), .PIJ(
        \PGNET_P[1][9] ) );
  PG_BLOCK_23 pgi_1_11 ( .PIK(\PGNET_P[0][11] ), .GIK(\PGNET_G[0][11] ), 
        .PK1J(\PGNET_P[0][10] ), .GK1J(\PGNET_G[0][10] ), .GIJ(
        \PGNET_G[1][11] ), .PIJ(\PGNET_P[1][11] ) );
  PG_BLOCK_22 pgi_1_13 ( .PIK(\PGNET_P[0][13] ), .GIK(\PGNET_G[0][13] ), 
        .PK1J(\PGNET_P[0][12] ), .GK1J(\PGNET_G[0][12] ), .GIJ(
        \PGNET_G[1][13] ), .PIJ(\PGNET_P[1][13] ) );
  PG_BLOCK_21 pgi_1_15 ( .PIK(\PGNET_P[0][15] ), .GIK(\PGNET_G[0][15] ), 
        .PK1J(\PGNET_P[0][14] ), .GK1J(\PGNET_G[0][14] ), .GIJ(
        \PGNET_G[1][15] ), .PIJ(\PGNET_P[1][15] ) );
  PG_BLOCK_20 pgi_1_17 ( .PIK(\PGNET_P[0][17] ), .GIK(\PGNET_G[0][17] ), 
        .PK1J(\PGNET_P[0][16] ), .GK1J(\PGNET_G[0][16] ), .GIJ(
        \PGNET_G[1][17] ), .PIJ(\PGNET_P[1][17] ) );
  PG_BLOCK_19 pgi_1_19 ( .PIK(\PGNET_P[0][19] ), .GIK(\PGNET_G[0][19] ), 
        .PK1J(\PGNET_P[0][18] ), .GK1J(\PGNET_G[0][18] ), .GIJ(
        \PGNET_G[1][19] ), .PIJ(\PGNET_P[1][19] ) );
  PG_BLOCK_18 pgi_1_21 ( .PIK(\PGNET_P[0][21] ), .GIK(\PGNET_G[0][21] ), 
        .PK1J(\PGNET_P[0][20] ), .GK1J(\PGNET_G[0][20] ), .GIJ(
        \PGNET_G[1][21] ), .PIJ(\PGNET_P[1][21] ) );
  PG_BLOCK_17 pgi_1_23 ( .PIK(\PGNET_P[0][23] ), .GIK(\PGNET_G[0][23] ), 
        .PK1J(\PGNET_P[0][22] ), .GK1J(\PGNET_G[0][22] ), .GIJ(
        \PGNET_G[1][23] ), .PIJ(\PGNET_P[1][23] ) );
  PG_BLOCK_16 pgi_1_25 ( .PIK(\PGNET_P[0][25] ), .GIK(\PGNET_G[0][25] ), 
        .PK1J(\PGNET_P[0][24] ), .GK1J(\PGNET_G[0][24] ), .GIJ(
        \PGNET_G[1][25] ), .PIJ(\PGNET_P[1][25] ) );
  PG_BLOCK_15 pgi_1_27 ( .PIK(\PGNET_P[0][27] ), .GIK(\PGNET_G[0][27] ), 
        .PK1J(\PGNET_P[0][26] ), .GK1J(\PGNET_G[0][26] ), .GIJ(
        \PGNET_G[1][27] ), .PIJ(\PGNET_P[1][27] ) );
  PG_BLOCK_14 pgi_1_29 ( .PIK(\PGNET_P[0][29] ), .GIK(\PGNET_G[0][29] ), 
        .PK1J(\PGNET_P[0][28] ), .GK1J(\PGNET_G[0][28] ), .GIJ(
        \PGNET_G[1][29] ), .PIJ(\PGNET_P[1][29] ) );
  PG_BLOCK_13 pgi_1_31 ( .PIK(\PGNET_P[0][31] ), .GIK(\PGNET_G[0][31] ), 
        .PK1J(\PGNET_P[0][30] ), .GK1J(\PGNET_G[0][30] ), .GIJ(
        \PGNET_G[1][31] ), .PIJ(\PGNET_P[1][31] ) );
  G_BLOCK_8 gi_2_3 ( .PIK(\PGNET_P[1][3] ), .GIK(\PGNET_G[1][3] ), .GK1J(
        \PGNET_G[1][1] ), .GIJ(Co[1]) );
  PG_BLOCK_12 pgi_2_7 ( .PIK(\PGNET_P[1][7] ), .GIK(\PGNET_G[1][7] ), .PK1J(
        \PGNET_P[1][5] ), .GK1J(\PGNET_G[1][5] ), .GIJ(\PGNET_G[2][7] ), .PIJ(
        \PGNET_P[2][7] ) );
  PG_BLOCK_11 pgi_2_11 ( .PIK(\PGNET_P[1][11] ), .GIK(\PGNET_G[1][11] ), 
        .PK1J(\PGNET_P[1][9] ), .GK1J(\PGNET_G[1][9] ), .GIJ(\PGNET_G[2][11] ), 
        .PIJ(\PGNET_P[3][11] ) );
  PG_BLOCK_10 pgi_2_15 ( .PIK(\PGNET_P[1][15] ), .GIK(\PGNET_G[1][15] ), 
        .PK1J(\PGNET_P[1][13] ), .GK1J(\PGNET_G[1][13] ), .GIJ(
        \PGNET_G[2][15] ), .PIJ(\PGNET_P[2][15] ) );
  PG_BLOCK_9 pgi_2_19 ( .PIK(\PGNET_P[1][19] ), .GIK(\PGNET_G[1][19] ), .PK1J(
        \PGNET_P[1][17] ), .GK1J(\PGNET_G[1][17] ), .GIJ(\PGNET_G[2][19] ), 
        .PIJ(\PGNET_P[2][19] ) );
  PG_BLOCK_8 pgi_2_23 ( .PIK(\PGNET_P[1][23] ), .GIK(\PGNET_G[1][23] ), .PK1J(
        \PGNET_P[1][21] ), .GK1J(\PGNET_G[1][21] ), .GIJ(\PGNET_G[2][23] ), 
        .PIJ(\PGNET_P[2][23] ) );
  PG_BLOCK_7 pgi_2_27 ( .PIK(\PGNET_P[1][27] ), .GIK(\PGNET_G[1][27] ), .PK1J(
        \PGNET_P[1][25] ), .GK1J(\PGNET_G[1][25] ), .GIJ(\PGNET_G[2][27] ), 
        .PIJ(\PGNET_P[2][27] ) );
  PG_BLOCK_6 pgi_2_31 ( .PIK(\PGNET_P[1][31] ), .GIK(\PGNET_G[1][31] ), .PK1J(
        \PGNET_P[1][29] ), .GK1J(\PGNET_G[1][29] ), .GIJ(\PGNET_G[2][31] ), 
        .PIJ(\PGNET_P[2][31] ) );
  G_BLOCK_7 gi_3_7 ( .PIK(\PGNET_P[2][7] ), .GIK(\PGNET_G[2][7] ), .GK1J(Co[1]), .GIJ(Co[2]) );
  PG_BLOCK_5 pgi_3_15 ( .PIK(\PGNET_P[2][15] ), .GIK(\PGNET_G[2][15] ), .PK1J(
        \PGNET_P[3][11] ), .GK1J(\PGNET_G[2][11] ), .GIJ(\PGNET_G[3][15] ), 
        .PIJ(\PGNET_P[3][15] ) );
  PG_BLOCK_4 pgi_3_23 ( .PIK(\PGNET_P[2][23] ), .GIK(\PGNET_G[2][23] ), .PK1J(
        \PGNET_P[2][19] ), .GK1J(\PGNET_G[2][19] ), .GIJ(\PGNET_G[3][23] ), 
        .PIJ(\PGNET_P[3][23] ) );
  PG_BLOCK_3 pgi_3_31 ( .PIK(\PGNET_P[2][31] ), .GIK(\PGNET_G[2][31] ), .PK1J(
        \PGNET_P[2][27] ), .GK1J(\PGNET_G[2][27] ), .GIJ(\PGNET_G[3][31] ), 
        .PIJ(\PGNET_P[3][31] ) );
  G_BLOCK_6 gi_4_11 ( .PIK(\PGNET_P[3][11] ), .GIK(\PGNET_G[2][11] ), .GK1J(
        Co[2]), .GIJ(Co[3]) );
  G_BLOCK_5 gi_4_15 ( .PIK(\PGNET_P[3][15] ), .GIK(\PGNET_G[3][15] ), .GK1J(
        Co[2]), .GIJ(Co[4]) );
  PG_BLOCK_2 pgi_4_27 ( .PIK(\PGNET_P[2][27] ), .GIK(\PGNET_G[2][27] ), .PK1J(
        \PGNET_P[3][23] ), .GK1J(\PGNET_G[3][23] ), .GIJ(\PGNET_G[4][27] ), 
        .PIJ(\PGNET_P[4][27] ) );
  PG_BLOCK_1 pgi_4_31 ( .PIK(\PGNET_P[3][31] ), .GIK(\PGNET_G[3][31] ), .PK1J(
        \PGNET_P[3][23] ), .GK1J(\PGNET_G[3][23] ), .GIJ(\PGNET_G[4][31] ), 
        .PIJ(\PGNET_P[4][31] ) );
  G_BLOCK_4 gi_5_19 ( .PIK(\PGNET_P[2][19] ), .GIK(\PGNET_G[2][19] ), .GK1J(
        Co[4]), .GIJ(Co[5]) );
  G_BLOCK_3 gi_5_23 ( .PIK(\PGNET_P[3][23] ), .GIK(\PGNET_G[3][23] ), .GK1J(
        Co[4]), .GIJ(Co[6]) );
  G_BLOCK_2 gi_5_27 ( .PIK(\PGNET_P[4][27] ), .GIK(\PGNET_G[4][27] ), .GK1J(
        Co[4]), .GIJ(Co[7]) );
  G_BLOCK_1 gi_5_31 ( .PIK(\PGNET_P[4][31] ), .GIK(\PGNET_G[4][31] ), .GK1J(
        Co[4]), .GIJ(Co[8]) );
  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(\PGNET_G[0][0] ) );
  OAI21_X1 U2 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n3) );
  INV_X1 U3 ( .A(B[0]), .ZN(n2) );
  INV_X1 U4 ( .A(A[0]), .ZN(n1) );
endmodule


module FA_0 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_63 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_62 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_61 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_0 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_0 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_63 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_62 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_61 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_60 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_59 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_58 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_57 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_15 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_60 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_59 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_58 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_57 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_32 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_0 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_0 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_15 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_0 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_56 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_55 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_54 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_53 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_14 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_56 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_55 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_54 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_53 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_52 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_51 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_50 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_49 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_13 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_52 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_51 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_50 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_49 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_7 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_14 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_13 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_7 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_48 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_47 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_46 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_45 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_12 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_48 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_47 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_46 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_45 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_44 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_43 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_42 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_41 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_11 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_44 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_43 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_42 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_41 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_6 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_12 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_11 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_6 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_40 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_39 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_38 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_37 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_10 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_40 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_39 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_38 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_37 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_36 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_35 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_34 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_33 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_9 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_36 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_35 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_34 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_33 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_5 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_10 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_9 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_5 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_32 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_31 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_30 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_29 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_8 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_32 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_31 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_30 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_29 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_28 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_27 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_26 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_25 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_7 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_28 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_27 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_26 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_25 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_4 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_8 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_7 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_4 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_24 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_23 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_22 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_21 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_6 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_24 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_23 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_22 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_21 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_20 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_19 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_18 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_17 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_5 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_20 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_19 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_18 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_17 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_3 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_6 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_5 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_3 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_16 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_15 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_14 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_13 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_4 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_16 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_15 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_14 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_13 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_12 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_11 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_10 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_9 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_3 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_12 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_11 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(
        sum[1]) );
  FA_10 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(
        sum[2]) );
  FA_9 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_2 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_4 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_3 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_2 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module FA_8 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_7 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_6 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_5 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_2 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_8 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_7 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(sum[1]) );
  FA_6 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(sum[2]) );
  FA_5 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module FA_4 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_3 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_2 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FA_1 ( a, b, c_in, c_out, s );
  input a, b, c_in;
  output c_out, s;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(c_in), .B(n1), .Z(s) );
  INV_X1 U2 ( .A(n2), .ZN(c_out) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(c_in), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module RCA_size4_1 ( a, b, c_in, c_out, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  FA_4 fa_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .c_out(temp[1]), .s(sum[0])
         );
  FA_3 fa_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .c_out(temp[2]), .s(sum[1]) );
  FA_2 fa_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .c_out(temp[3]), .s(sum[2]) );
  FA_1 fa_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .c_out(c_out), .s(sum[3])
         );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module SUM_BLOCK_K4_1 ( a, b, C_gen, sum );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input C_gen;

  wire   [3:0] SUM1;
  wire   [3:0] SUM2;

  RCA_size4_2 RCA_CIN0 ( .a(a), .b(b), .c_in(1'b0), .sum(SUM1) );
  RCA_size4_1 RCA_CIN1 ( .a(a), .b(b), .c_in(1'b1), .sum(SUM2) );
  MUX21_GENERIC_NBIT4_1 MPX ( .A(SUM2), .B(SUM1), .SEL(C_gen), .Y(sum) );
endmodule


module SUM_GENERATOR_N32_K4 ( carries, A, B, SUM );
  input [7:0] carries;
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;


  SUM_BLOCK_K4_0 SBi_0 ( .a(A[3:0]), .b(B[3:0]), .C_gen(carries[0]), .sum(
        SUM[3:0]) );
  SUM_BLOCK_K4_7 SBi_1 ( .a(A[7:4]), .b(B[7:4]), .C_gen(carries[1]), .sum(
        SUM[7:4]) );
  SUM_BLOCK_K4_6 SBi_2 ( .a(A[11:8]), .b(B[11:8]), .C_gen(carries[2]), .sum(
        SUM[11:8]) );
  SUM_BLOCK_K4_5 SBi_3 ( .a(A[15:12]), .b(B[15:12]), .C_gen(carries[3]), .sum(
        SUM[15:12]) );
  SUM_BLOCK_K4_4 SBi_4 ( .a(A[19:16]), .b(B[19:16]), .C_gen(carries[4]), .sum(
        SUM[19:16]) );
  SUM_BLOCK_K4_3 SBi_5 ( .a(A[23:20]), .b(B[23:20]), .C_gen(carries[5]), .sum(
        SUM[23:20]) );
  SUM_BLOCK_K4_2 SBi_6 ( .a(A[27:24]), .b(B[27:24]), .C_gen(carries[6]), .sum(
        SUM[27:24]) );
  SUM_BLOCK_K4_1 SBi_7 ( .a(A[31:28]), .b(B[31:28]), .C_gen(carries[7]), .sum(
        SUM[31:28]) );
endmodule


module P4Adder_N32_K4 ( A, B, CIN, Cout, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CIN;
  output Cout;

  wire   [31:0] Bx_s;
  wire   [7:0] carries_s;

  xorGrid_N32 CPL ( .B(B), .Cin(CIN), .Bx(Bx_s) );
  CARRY_GENERATOR_NBIT32_NBLOCK4 CG ( .A(A), .B(Bx_s), .Cin(CIN), .Co({Cout, 
        carries_s}) );
  SUM_GENERATOR_N32_K4 SG ( .carries(carries_s), .A(A), .B(Bx_s), .SUM(SUM) );
endmodule


module ShifterT2_N32 ( A, B, sel, \output  );
  input [31:0] A;
  input [4:0] B;
  input [1:0] sel;
  output [31:0] \output ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298;

  AOI221_X1 U2 ( .B1(n84), .B2(A[8]), .C1(n85), .C2(A[0]), .A(n96), .ZN(n158)
         );
  AOI221_X1 U3 ( .B1(n3), .B2(n250), .C1(n223), .C2(n15), .A(n269), .ZN(n268)
         );
  AOI221_X1 U4 ( .B1(n28), .B2(n14), .C1(n17), .C2(n15), .A(n29), .ZN(n23) );
  AOI221_X1 U5 ( .B1(n16), .B2(n4), .C1(n5), .C2(n25), .A(n34), .ZN(n33) );
  AOI221_X1 U6 ( .B1(n84), .B2(A[13]), .C1(n85), .C2(A[5]), .A(n96), .ZN(n114)
         );
  AOI221_X1 U7 ( .B1(n84), .B2(A[12]), .C1(n85), .C2(A[4]), .A(n96), .ZN(n125)
         );
  AOI221_X1 U8 ( .B1(n84), .B2(A[11]), .C1(n85), .C2(A[3]), .A(n96), .ZN(n134)
         );
  AOI221_X1 U9 ( .B1(n84), .B2(A[10]), .C1(n85), .C2(A[2]), .A(n96), .ZN(n142)
         );
  AOI221_X1 U10 ( .B1(n84), .B2(A[9]), .C1(n85), .C2(A[1]), .A(n96), .ZN(n150)
         );
  NOR4_X2 U11 ( .A1(n159), .A2(n160), .A3(sel[0]), .A4(sel[1]), .ZN(n85) );
  NOR3_X2 U12 ( .A1(n81), .A2(n103), .A3(n237), .ZN(n96) );
  INV_X2 U13 ( .A(n20), .ZN(n28) );
  INV_X2 U14 ( .A(n31), .ZN(n16) );
  NOR3_X4 U15 ( .A1(n286), .A2(B[0]), .A3(n288), .ZN(n116) );
  OAI21_X2 U16 ( .B1(n293), .B2(n294), .A(n295), .ZN(n6) );
  OAI21_X4 U17 ( .B1(n287), .B2(n290), .A(n291), .ZN(n39) );
  NOR2_X4 U18 ( .A1(n294), .A2(B[0]), .ZN(n3) );
  OAI21_X4 U19 ( .B1(n287), .B2(n293), .A(n298), .ZN(n15) );
  NAND2_X2 U20 ( .A1(n276), .A2(n160), .ZN(n82) );
  OAI21_X4 U21 ( .B1(n290), .B2(n294), .A(n297), .ZN(n25) );
  NAND2_X1 U22 ( .A1(n1), .A2(n2), .ZN(\output [9]) );
  AOI221_X1 U23 ( .B1(n3), .B2(n4), .C1(n5), .C2(n6), .A(n7), .ZN(n2) );
  OAI222_X1 U24 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C1(n12), .C2(n13), 
        .ZN(n7) );
  AOI221_X1 U25 ( .B1(n14), .B2(n15), .C1(n16), .C2(n17), .A(n18), .ZN(n1) );
  OAI22_X1 U26 ( .A1(n19), .A2(n20), .B1(n21), .B2(n22), .ZN(n18) );
  NAND2_X1 U27 ( .A1(n23), .A2(n24), .ZN(\output [8]) );
  AOI221_X1 U28 ( .B1(n4), .B2(n25), .C1(n3), .C2(n5), .A(n26), .ZN(n24) );
  OAI222_X1 U29 ( .A1(n9), .A2(n13), .B1(n8), .B2(n10), .C1(n27), .C2(n12), 
        .ZN(n26) );
  OAI22_X1 U30 ( .A1(n30), .A2(n11), .B1(n22), .B2(n31), .ZN(n29) );
  NAND2_X1 U31 ( .A1(n32), .A2(n33), .ZN(\output [7]) );
  OAI222_X1 U32 ( .A1(n27), .A2(n9), .B1(n10), .B2(n13), .C1(n12), .C2(n35), 
        .ZN(n34) );
  INV_X1 U33 ( .A(n36), .ZN(n12) );
  INV_X1 U34 ( .A(n37), .ZN(n9) );
  AOI221_X1 U35 ( .B1(n38), .B2(n39), .C1(n40), .C2(n41), .A(n42), .ZN(n32) );
  OAI22_X1 U36 ( .A1(n43), .A2(n22), .B1(n44), .B2(n20), .ZN(n42) );
  NAND3_X1 U37 ( .A1(n45), .A2(n46), .A3(n47), .ZN(\output [6]) );
  AOI221_X1 U38 ( .B1(n48), .B2(n41), .C1(n40), .C2(n39), .A(n49), .ZN(n47) );
  OAI22_X1 U39 ( .A1(n30), .A2(n13), .B1(n22), .B2(n20), .ZN(n49) );
  AOI222_X1 U40 ( .A1(n36), .A2(n25), .B1(n50), .B2(n6), .C1(n3), .C2(n37), 
        .ZN(n46) );
  AOI22_X1 U41 ( .A1(n4), .A2(n15), .B1(n16), .B2(n5), .ZN(n45) );
  NAND3_X1 U42 ( .A1(n51), .A2(n52), .A3(n53), .ZN(\output [5]) );
  AOI221_X1 U43 ( .B1(n38), .B2(n6), .C1(n54), .C2(n41), .A(n55), .ZN(n53) );
  OAI22_X1 U44 ( .A1(n13), .A2(n56), .B1(n8), .B2(n57), .ZN(n55) );
  AOI222_X1 U45 ( .A1(n16), .A2(n36), .B1(n3), .B2(n50), .C1(n37), .C2(n25), 
        .ZN(n52) );
  AOI22_X1 U46 ( .A1(n28), .A2(n4), .B1(n5), .B2(n15), .ZN(n51) );
  NAND3_X1 U47 ( .A1(n58), .A2(n59), .A3(n60), .ZN(\output [4]) );
  AOI221_X1 U48 ( .B1(n61), .B2(n41), .C1(n54), .C2(n39), .A(n62), .ZN(n60) );
  OAI22_X1 U49 ( .A1(n13), .A2(n57), .B1(n27), .B2(n56), .ZN(n62) );
  AOI222_X1 U50 ( .A1(n36), .A2(n15), .B1(n50), .B2(n25), .C1(n16), .C2(n37), 
        .ZN(n59) );
  AOI22_X1 U51 ( .A1(n28), .A2(n5), .B1(n3), .B2(n38), .ZN(n58) );
  NAND3_X1 U52 ( .A1(n63), .A2(n64), .A3(n65), .ZN(\output [3]) );
  AOI221_X1 U53 ( .B1(n61), .B2(n39), .C1(n48), .C2(n6), .A(n66), .ZN(n65) );
  OAI22_X1 U54 ( .A1(n35), .A2(n56), .B1(n13), .B2(n67), .ZN(n66) );
  AOI222_X1 U55 ( .A1(n37), .A2(n15), .B1(A[3]), .B2(n41), .C1(n16), .C2(n50), 
        .ZN(n64) );
  AOI22_X1 U56 ( .A1(n28), .A2(n36), .B1(n38), .B2(n25), .ZN(n63) );
  NAND3_X1 U57 ( .A1(n68), .A2(n69), .A3(n70), .ZN(\output [31]) );
  AOI221_X1 U58 ( .B1(n3), .B2(n71), .C1(n72), .C2(n6), .A(n73), .ZN(n70) );
  OAI22_X1 U59 ( .A1(n8), .A2(n74), .B1(n75), .B2(n13), .ZN(n73) );
  AOI22_X1 U60 ( .A1(n76), .A2(n77), .B1(n78), .B2(n15), .ZN(n69) );
  OAI221_X1 U61 ( .B1(n79), .B2(n80), .C1(n81), .C2(n82), .A(n83), .ZN(n77) );
  AOI222_X1 U62 ( .A1(n84), .A2(A[15]), .B1(n85), .B2(A[7]), .C1(sel[0]), .C2(
        n86), .ZN(n83) );
  AOI22_X1 U63 ( .A1(n16), .A2(n87), .B1(n88), .B2(n25), .ZN(n68) );
  NAND2_X1 U64 ( .A1(n89), .A2(n90), .ZN(\output [30]) );
  AOI221_X1 U65 ( .B1(n71), .B2(n25), .C1(n3), .C2(n72), .A(n91), .ZN(n90) );
  INV_X1 U66 ( .A(n92), .ZN(n91) );
  AOI222_X1 U67 ( .A1(n15), .A2(n87), .B1(n78), .B2(n28), .C1(n88), .C2(n16), 
        .ZN(n92) );
  OAI221_X1 U68 ( .B1(n79), .B2(n93), .C1(n82), .C2(n94), .A(n95), .ZN(n78) );
  AOI221_X1 U69 ( .B1(n84), .B2(A[14]), .C1(n85), .C2(A[6]), .A(n96), .ZN(n95)
         );
  INV_X1 U70 ( .A(A[30]), .ZN(n94) );
  AOI221_X1 U71 ( .B1(n86), .B2(n39), .C1(n41), .C2(n97), .A(n98), .ZN(n89) );
  OAI22_X1 U72 ( .A1(n74), .A2(n13), .B1(n27), .B2(n75), .ZN(n98) );
  NAND2_X1 U73 ( .A1(n99), .A2(n100), .ZN(\output [2]) );
  AOI221_X1 U74 ( .B1(n28), .B2(n37), .C1(n16), .C2(n38), .A(n101), .ZN(n100)
         );
  OAI22_X1 U75 ( .A1(n43), .A2(n10), .B1(n102), .B2(n103), .ZN(n101) );
  AOI22_X1 U76 ( .A1(A[2]), .A2(n41), .B1(A[3]), .B2(n39), .ZN(n102) );
  INV_X1 U77 ( .A(n50), .ZN(n10) );
  AOI221_X1 U78 ( .B1(n48), .B2(n3), .C1(n40), .C2(n25), .A(n104), .ZN(n99) );
  OAI22_X1 U79 ( .A1(n13), .A2(n105), .B1(n27), .B2(n67), .ZN(n104) );
  NAND3_X1 U80 ( .A1(n106), .A2(n107), .A3(n108), .ZN(\output [29]) );
  AOI221_X1 U81 ( .B1(n72), .B2(n25), .C1(n3), .C2(n109), .A(n110), .ZN(n108)
         );
  INV_X1 U82 ( .A(n111), .ZN(n110) );
  AOI222_X1 U83 ( .A1(n15), .A2(n88), .B1(n87), .B2(n28), .C1(n71), .C2(n16), 
        .ZN(n111) );
  OAI221_X1 U84 ( .B1(n79), .B2(n112), .C1(n82), .C2(n113), .A(n114), .ZN(n87)
         );
  INV_X1 U85 ( .A(A[29]), .ZN(n113) );
  AOI22_X1 U86 ( .A1(n115), .A2(n6), .B1(n116), .B2(n86), .ZN(n107) );
  AOI22_X1 U87 ( .A1(n97), .A2(n39), .B1(n41), .B2(n117), .ZN(n106) );
  NAND3_X1 U88 ( .A1(n118), .A2(n119), .A3(n120), .ZN(\output [28]) );
  INV_X1 U89 ( .A(n121), .ZN(n120) );
  OAI221_X1 U90 ( .B1(n75), .B2(n21), .C1(n35), .C2(n74), .A(n122), .ZN(n121)
         );
  AOI222_X1 U91 ( .A1(n15), .A2(n71), .B1(n88), .B2(n28), .C1(n72), .C2(n16), 
        .ZN(n122) );
  OAI221_X1 U92 ( .B1(n79), .B2(n123), .C1(n82), .C2(n124), .A(n125), .ZN(n88)
         );
  INV_X1 U93 ( .A(A[28]), .ZN(n124) );
  INV_X1 U94 ( .A(n115), .ZN(n74) );
  INV_X1 U95 ( .A(n109), .ZN(n75) );
  AOI22_X1 U96 ( .A1(n86), .A2(n6), .B1(n116), .B2(n97), .ZN(n119) );
  AOI22_X1 U97 ( .A1(n117), .A2(n39), .B1(n41), .B2(n126), .ZN(n118) );
  NAND3_X1 U98 ( .A1(n127), .A2(n128), .A3(n129), .ZN(\output [27]) );
  AOI221_X1 U99 ( .B1(n115), .B2(n25), .C1(n3), .C2(n86), .A(n130), .ZN(n129)
         );
  INV_X1 U100 ( .A(n131), .ZN(n130) );
  AOI222_X1 U101 ( .A1(n15), .A2(n72), .B1(n71), .B2(n28), .C1(n109), .C2(n16), 
        .ZN(n131) );
  OAI221_X1 U102 ( .B1(n79), .B2(n132), .C1(n82), .C2(n133), .A(n134), .ZN(n71) );
  INV_X1 U103 ( .A(A[27]), .ZN(n133) );
  AOI22_X1 U104 ( .A1(n97), .A2(n6), .B1(n116), .B2(n117), .ZN(n128) );
  AOI22_X1 U105 ( .A1(n126), .A2(n39), .B1(n41), .B2(n135), .ZN(n127) );
  NAND4_X1 U106 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(\output [26]) );
  AOI222_X1 U107 ( .A1(n16), .A2(n115), .B1(n28), .B2(n72), .C1(n109), .C2(n15), .ZN(n139) );
  OAI221_X1 U108 ( .B1(n79), .B2(n140), .C1(n82), .C2(n141), .A(n142), .ZN(n72) );
  INV_X1 U109 ( .A(A[26]), .ZN(n141) );
  AOI22_X1 U110 ( .A1(n86), .A2(n25), .B1(n3), .B2(n97), .ZN(n138) );
  AOI22_X1 U111 ( .A1(n117), .A2(n6), .B1(n116), .B2(n126), .ZN(n137) );
  AOI22_X1 U112 ( .A1(n135), .A2(n39), .B1(n41), .B2(n143), .ZN(n136) );
  NAND4_X1 U113 ( .A1(n144), .A2(n145), .A3(n146), .A4(n147), .ZN(\output [25]) );
  AOI222_X1 U114 ( .A1(n16), .A2(n86), .B1(n28), .B2(n109), .C1(n115), .C2(n15), .ZN(n147) );
  OAI221_X1 U115 ( .B1(n79), .B2(n148), .C1(n82), .C2(n149), .A(n150), .ZN(
        n109) );
  INV_X1 U116 ( .A(A[25]), .ZN(n149) );
  AOI22_X1 U117 ( .A1(n97), .A2(n25), .B1(n3), .B2(n117), .ZN(n146) );
  AOI22_X1 U118 ( .A1(n126), .A2(n6), .B1(n116), .B2(n135), .ZN(n145) );
  AOI22_X1 U119 ( .A1(n143), .A2(n39), .B1(n41), .B2(n151), .ZN(n144) );
  NAND4_X1 U120 ( .A1(n152), .A2(n153), .A3(n154), .A4(n155), .ZN(\output [24]) );
  AOI222_X1 U121 ( .A1(n16), .A2(n97), .B1(n28), .B2(n115), .C1(n86), .C2(n15), 
        .ZN(n155) );
  OAI221_X1 U122 ( .B1(n79), .B2(n156), .C1(n82), .C2(n157), .A(n158), .ZN(
        n115) );
  INV_X1 U123 ( .A(A[24]), .ZN(n157) );
  AOI22_X1 U124 ( .A1(n117), .A2(n25), .B1(n3), .B2(n126), .ZN(n154) );
  AOI22_X1 U125 ( .A1(n135), .A2(n6), .B1(n116), .B2(n143), .ZN(n153) );
  AOI22_X1 U126 ( .A1(n151), .A2(n39), .B1(n41), .B2(n161), .ZN(n152) );
  NAND4_X1 U127 ( .A1(n162), .A2(n163), .A3(n164), .A4(n165), .ZN(\output [23]) );
  AOI222_X1 U128 ( .A1(n16), .A2(n117), .B1(n28), .B2(n86), .C1(n97), .C2(n15), 
        .ZN(n165) );
  OAI221_X1 U129 ( .B1(n79), .B2(n166), .C1(n82), .C2(n80), .A(n167), .ZN(n86)
         );
  AOI221_X1 U130 ( .B1(n84), .B2(A[7]), .C1(n168), .C2(A[31]), .A(n169), .ZN(
        n167) );
  INV_X1 U131 ( .A(A[23]), .ZN(n80) );
  AOI22_X1 U132 ( .A1(n126), .A2(n25), .B1(n3), .B2(n135), .ZN(n164) );
  AOI22_X1 U133 ( .A1(n143), .A2(n6), .B1(n116), .B2(n151), .ZN(n163) );
  AOI22_X1 U134 ( .A1(n161), .A2(n39), .B1(n41), .B2(n170), .ZN(n162) );
  NAND3_X1 U135 ( .A1(n171), .A2(n172), .A3(n173), .ZN(\output [22]) );
  AOI221_X1 U136 ( .B1(n151), .B2(n6), .C1(n116), .C2(n161), .A(n174), .ZN(
        n173) );
  OAI22_X1 U137 ( .A1(n175), .A2(n11), .B1(n8), .B2(n176), .ZN(n174) );
  AOI222_X1 U138 ( .A1(n16), .A2(n126), .B1(n28), .B2(n97), .C1(n117), .C2(n15), .ZN(n172) );
  OAI221_X1 U139 ( .B1(n79), .B2(n177), .C1(n82), .C2(n93), .A(n178), .ZN(n97)
         );
  AOI221_X1 U140 ( .B1(n84), .B2(A[6]), .C1(A[30]), .C2(n168), .A(n169), .ZN(
        n178) );
  INV_X1 U141 ( .A(A[22]), .ZN(n93) );
  AOI22_X1 U142 ( .A1(n135), .A2(n25), .B1(n3), .B2(n143), .ZN(n171) );
  NAND3_X1 U143 ( .A1(n179), .A2(n180), .A3(n181), .ZN(\output [21]) );
  AOI221_X1 U144 ( .B1(n161), .B2(n6), .C1(n116), .C2(n170), .A(n182), .ZN(
        n181) );
  OAI22_X1 U145 ( .A1(n183), .A2(n11), .B1(n8), .B2(n175), .ZN(n182) );
  AOI222_X1 U146 ( .A1(n16), .A2(n135), .B1(n28), .B2(n117), .C1(n126), .C2(
        n15), .ZN(n180) );
  OAI221_X1 U147 ( .B1(n184), .B2(n79), .C1(n82), .C2(n112), .A(n185), .ZN(
        n117) );
  AOI221_X1 U148 ( .B1(n84), .B2(A[5]), .C1(A[29]), .C2(n168), .A(n169), .ZN(
        n185) );
  INV_X1 U149 ( .A(A[21]), .ZN(n112) );
  AOI22_X1 U150 ( .A1(n143), .A2(n25), .B1(n3), .B2(n151), .ZN(n179) );
  NAND3_X1 U151 ( .A1(n186), .A2(n187), .A3(n188), .ZN(\output [20]) );
  AOI221_X1 U152 ( .B1(n189), .B2(n39), .C1(n41), .C2(n190), .A(n191), .ZN(
        n188) );
  OAI22_X1 U153 ( .A1(n175), .A2(n13), .B1(n27), .B2(n176), .ZN(n191) );
  INV_X1 U154 ( .A(n170), .ZN(n176) );
  AOI222_X1 U155 ( .A1(n16), .A2(n143), .B1(n28), .B2(n126), .C1(n135), .C2(
        n15), .ZN(n187) );
  OAI221_X1 U156 ( .B1(n192), .B2(n79), .C1(n82), .C2(n123), .A(n193), .ZN(
        n126) );
  AOI221_X1 U157 ( .B1(n84), .B2(A[4]), .C1(A[28]), .C2(n168), .A(n169), .ZN(
        n193) );
  INV_X1 U158 ( .A(A[20]), .ZN(n123) );
  AOI22_X1 U159 ( .A1(n151), .A2(n25), .B1(n3), .B2(n161), .ZN(n186) );
  OAI211_X1 U160 ( .C1(n35), .C2(n67), .A(n194), .B(n195), .ZN(\output [1]) );
  AOI221_X1 U161 ( .B1(sel[0]), .B2(n196), .C1(n28), .C2(n50), .A(n197), .ZN(
        n195) );
  OAI22_X1 U162 ( .A1(n27), .A2(n105), .B1(n43), .B2(n30), .ZN(n197) );
  INV_X1 U163 ( .A(n38), .ZN(n30) );
  OAI221_X1 U164 ( .B1(n82), .B2(n198), .C1(n199), .C2(n200), .A(n201), .ZN(
        n50) );
  OAI222_X1 U165 ( .A1(n8), .A2(n202), .B1(n198), .B2(n11), .C1(n203), .C2(n13), .ZN(n196) );
  AOI22_X1 U166 ( .A1(n40), .A2(n16), .B1(n48), .B2(n25), .ZN(n194) );
  INV_X1 U167 ( .A(n57), .ZN(n48) );
  INV_X1 U168 ( .A(n56), .ZN(n40) );
  NAND3_X1 U169 ( .A1(n204), .A2(n205), .A3(n206), .ZN(\output [19]) );
  AOI221_X1 U170 ( .B1(n190), .B2(n39), .C1(n41), .C2(n207), .A(n208), .ZN(
        n206) );
  OAI22_X1 U171 ( .A1(n183), .A2(n13), .B1(n27), .B2(n175), .ZN(n208) );
  INV_X1 U172 ( .A(n209), .ZN(n175) );
  AOI222_X1 U173 ( .A1(n16), .A2(n151), .B1(n28), .B2(n135), .C1(n143), .C2(
        n15), .ZN(n205) );
  OAI221_X1 U174 ( .B1(n210), .B2(n79), .C1(n82), .C2(n132), .A(n211), .ZN(
        n135) );
  AOI221_X1 U175 ( .B1(n84), .B2(A[3]), .C1(A[27]), .C2(n168), .A(n169), .ZN(
        n211) );
  INV_X1 U176 ( .A(A[19]), .ZN(n132) );
  AOI22_X1 U177 ( .A1(n161), .A2(n25), .B1(n3), .B2(n170), .ZN(n204) );
  NAND3_X1 U178 ( .A1(n212), .A2(n213), .A3(n214), .ZN(\output [18]) );
  AOI221_X1 U179 ( .B1(n207), .B2(n39), .C1(n41), .C2(n215), .A(n216), .ZN(
        n214) );
  OAI22_X1 U180 ( .A1(n217), .A2(n13), .B1(n27), .B2(n183), .ZN(n216) );
  INV_X1 U181 ( .A(n189), .ZN(n183) );
  AOI222_X1 U182 ( .A1(n16), .A2(n161), .B1(n28), .B2(n143), .C1(n151), .C2(
        n15), .ZN(n213) );
  OAI221_X1 U183 ( .B1(n218), .B2(n79), .C1(n82), .C2(n140), .A(n219), .ZN(
        n143) );
  AOI221_X1 U184 ( .B1(n84), .B2(A[2]), .C1(A[26]), .C2(n168), .A(n169), .ZN(
        n219) );
  INV_X1 U185 ( .A(A[18]), .ZN(n140) );
  AOI22_X1 U186 ( .A1(n170), .A2(n25), .B1(n3), .B2(n209), .ZN(n212) );
  NAND3_X1 U187 ( .A1(n220), .A2(n221), .A3(n222), .ZN(\output [17]) );
  AOI221_X1 U188 ( .B1(n215), .B2(n39), .C1(n41), .C2(n223), .A(n224), .ZN(
        n222) );
  OAI22_X1 U189 ( .A1(n225), .A2(n13), .B1(n27), .B2(n217), .ZN(n224) );
  INV_X1 U190 ( .A(n190), .ZN(n217) );
  AOI222_X1 U191 ( .A1(n16), .A2(n170), .B1(n28), .B2(n151), .C1(n161), .C2(
        n15), .ZN(n221) );
  OAI221_X1 U192 ( .B1(n200), .B2(n79), .C1(n82), .C2(n148), .A(n226), .ZN(
        n151) );
  AOI221_X1 U193 ( .B1(n84), .B2(A[1]), .C1(A[25]), .C2(n168), .A(n169), .ZN(
        n226) );
  INV_X1 U194 ( .A(A[17]), .ZN(n148) );
  AOI22_X1 U195 ( .A1(n209), .A2(n25), .B1(n3), .B2(n189), .ZN(n220) );
  NAND3_X1 U196 ( .A1(n227), .A2(n228), .A3(n229), .ZN(\output [16]) );
  AOI221_X1 U197 ( .B1(n41), .B2(n14), .C1(n223), .C2(n39), .A(n230), .ZN(n229) );
  OAI22_X1 U198 ( .A1(n231), .A2(n13), .B1(n27), .B2(n225), .ZN(n230) );
  INV_X1 U199 ( .A(n207), .ZN(n225) );
  INV_X1 U200 ( .A(n215), .ZN(n231) );
  AOI222_X1 U201 ( .A1(n16), .A2(n209), .B1(n28), .B2(n161), .C1(n170), .C2(
        n15), .ZN(n228) );
  OAI221_X1 U202 ( .B1(n79), .B2(n232), .C1(n82), .C2(n156), .A(n233), .ZN(
        n161) );
  AOI221_X1 U203 ( .B1(n84), .B2(A[0]), .C1(A[24]), .C2(n168), .A(n169), .ZN(
        n233) );
  INV_X1 U204 ( .A(n234), .ZN(n169) );
  OAI21_X1 U205 ( .B1(n235), .B2(B[3]), .A(n96), .ZN(n234) );
  AND2_X1 U206 ( .A1(n236), .A2(n160), .ZN(n168) );
  AND3_X1 U207 ( .A1(n103), .A2(n237), .A3(n235), .ZN(n84) );
  INV_X1 U208 ( .A(A[16]), .ZN(n156) );
  AOI22_X1 U209 ( .A1(n189), .A2(n25), .B1(n3), .B2(n190), .ZN(n227) );
  NAND3_X1 U210 ( .A1(n238), .A2(n239), .A3(n240), .ZN(\output [15]) );
  AOI221_X1 U211 ( .B1(n215), .B2(n6), .C1(n14), .C2(n39), .A(n241), .ZN(n240)
         );
  OAI22_X1 U212 ( .A1(n19), .A2(n13), .B1(n44), .B2(n11), .ZN(n241) );
  AOI222_X1 U213 ( .A1(n16), .A2(n189), .B1(n28), .B2(n170), .C1(n209), .C2(
        n15), .ZN(n239) );
  OAI211_X1 U214 ( .C1(n82), .C2(n166), .A(n242), .B(n243), .ZN(n170) );
  AOI22_X1 U215 ( .A1(A[7]), .A2(n244), .B1(A[23]), .B2(n236), .ZN(n243) );
  AOI22_X1 U216 ( .A1(n190), .A2(n25), .B1(n3), .B2(n207), .ZN(n238) );
  NAND4_X1 U217 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .ZN(\output [14]) );
  AOI222_X1 U218 ( .A1(n16), .A2(n190), .B1(n28), .B2(n209), .C1(n189), .C2(
        n15), .ZN(n248) );
  OAI211_X1 U219 ( .C1(n82), .C2(n177), .A(n242), .B(n249), .ZN(n209) );
  AOI22_X1 U220 ( .A1(A[6]), .A2(n244), .B1(A[22]), .B2(n236), .ZN(n249) );
  AOI22_X1 U221 ( .A1(n207), .A2(n25), .B1(n3), .B2(n215), .ZN(n247) );
  AOI22_X1 U222 ( .A1(n116), .A2(n14), .B1(n17), .B2(n39), .ZN(n246) );
  AOI22_X1 U223 ( .A1(n41), .A2(n250), .B1(n223), .B2(n6), .ZN(n245) );
  NAND3_X1 U224 ( .A1(n251), .A2(n252), .A3(n253), .ZN(\output [13]) );
  AOI221_X1 U225 ( .B1(n14), .B2(n6), .C1(n116), .C2(n17), .A(n254), .ZN(n253)
         );
  OAI22_X1 U226 ( .A1(n19), .A2(n35), .B1(n8), .B2(n22), .ZN(n254) );
  INV_X1 U227 ( .A(n250), .ZN(n22) );
  INV_X1 U228 ( .A(n3), .ZN(n35) );
  INV_X1 U229 ( .A(n223), .ZN(n19) );
  AOI222_X1 U230 ( .A1(n16), .A2(n207), .B1(n28), .B2(n189), .C1(n190), .C2(
        n15), .ZN(n252) );
  OAI211_X1 U231 ( .C1(n82), .C2(n184), .A(n242), .B(n255), .ZN(n189) );
  AOI22_X1 U232 ( .A1(n244), .A2(A[5]), .B1(A[21]), .B2(n236), .ZN(n255) );
  AOI22_X1 U233 ( .A1(n215), .A2(n25), .B1(n41), .B2(n4), .ZN(n251) );
  NAND4_X1 U234 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(\output [12]) );
  AOI222_X1 U235 ( .A1(n16), .A2(n215), .B1(n28), .B2(n190), .C1(n207), .C2(
        n15), .ZN(n259) );
  OAI211_X1 U236 ( .C1(n82), .C2(n192), .A(n242), .B(n260), .ZN(n190) );
  AOI22_X1 U237 ( .A1(n244), .A2(A[4]), .B1(A[20]), .B2(n236), .ZN(n260) );
  AOI22_X1 U238 ( .A1(n4), .A2(n39), .B1(n41), .B2(n5), .ZN(n258) );
  AOI22_X1 U239 ( .A1(n3), .A2(n14), .B1(n17), .B2(n6), .ZN(n257) );
  AOI22_X1 U240 ( .A1(n116), .A2(n250), .B1(n223), .B2(n25), .ZN(n256) );
  NAND4_X1 U241 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(\output [11]) );
  AOI222_X1 U242 ( .A1(n41), .A2(n36), .B1(n28), .B2(n207), .C1(n215), .C2(n15), .ZN(n264) );
  OAI211_X1 U243 ( .C1(n82), .C2(n210), .A(n242), .B(n265), .ZN(n207) );
  AOI22_X1 U244 ( .A1(n244), .A2(A[3]), .B1(A[19]), .B2(n236), .ZN(n265) );
  AOI22_X1 U245 ( .A1(n116), .A2(n4), .B1(n5), .B2(n39), .ZN(n263) );
  AOI22_X1 U246 ( .A1(n14), .A2(n25), .B1(n3), .B2(n17), .ZN(n262) );
  AOI22_X1 U247 ( .A1(n250), .A2(n6), .B1(n16), .B2(n223), .ZN(n261) );
  NAND3_X1 U248 ( .A1(n266), .A2(n267), .A3(n268), .ZN(\output [10]) );
  OAI22_X1 U249 ( .A1(n21), .A2(n44), .B1(n270), .B2(n31), .ZN(n269) );
  INV_X1 U250 ( .A(n14), .ZN(n270) );
  OAI211_X1 U251 ( .C1(n82), .C2(n232), .A(n242), .B(n271), .ZN(n14) );
  AOI22_X1 U252 ( .A1(A[0]), .A2(n244), .B1(A[16]), .B2(n236), .ZN(n271) );
  INV_X1 U253 ( .A(n17), .ZN(n44) );
  OAI221_X1 U254 ( .B1(n82), .B2(n272), .C1(n199), .C2(n166), .A(n201), .ZN(
        n17) );
  INV_X1 U255 ( .A(A[15]), .ZN(n166) );
  INV_X1 U256 ( .A(A[7]), .ZN(n272) );
  INV_X1 U257 ( .A(n25), .ZN(n21) );
  OAI211_X1 U258 ( .C1(n82), .C2(n200), .A(n242), .B(n273), .ZN(n223) );
  AOI22_X1 U259 ( .A1(n244), .A2(A[1]), .B1(A[17]), .B2(n236), .ZN(n273) );
  INV_X1 U260 ( .A(A[9]), .ZN(n200) );
  OAI221_X1 U261 ( .B1(n82), .B2(n274), .C1(n199), .C2(n177), .A(n201), .ZN(
        n250) );
  INV_X1 U262 ( .A(A[14]), .ZN(n177) );
  INV_X1 U263 ( .A(A[6]), .ZN(n274) );
  AOI222_X1 U264 ( .A1(n36), .A2(n39), .B1(n41), .B2(n37), .C1(n28), .C2(n215), 
        .ZN(n267) );
  OAI211_X1 U265 ( .C1(n82), .C2(n218), .A(n242), .B(n275), .ZN(n215) );
  AOI22_X1 U266 ( .A1(n244), .A2(A[2]), .B1(A[18]), .B2(n236), .ZN(n275) );
  NOR2_X1 U267 ( .A1(n103), .A2(B[4]), .ZN(n236) );
  INV_X1 U268 ( .A(n79), .ZN(n244) );
  NAND2_X1 U269 ( .A1(n276), .A2(B[3]), .ZN(n79) );
  AOI21_X1 U270 ( .B1(n96), .B2(n235), .A(n277), .ZN(n242) );
  INV_X1 U271 ( .A(n201), .ZN(n277) );
  OAI221_X1 U272 ( .B1(n82), .B2(n202), .C1(n199), .C2(n218), .A(n201), .ZN(
        n37) );
  INV_X1 U273 ( .A(A[10]), .ZN(n218) );
  INV_X1 U274 ( .A(n11), .ZN(n41) );
  OAI221_X1 U275 ( .B1(n82), .B2(n203), .C1(n199), .C2(n210), .A(n201), .ZN(
        n36) );
  INV_X1 U276 ( .A(A[11]), .ZN(n210) );
  AOI22_X1 U277 ( .A1(n4), .A2(n6), .B1(n116), .B2(n5), .ZN(n266) );
  OAI221_X1 U278 ( .B1(n82), .B2(n278), .C1(n199), .C2(n192), .A(n201), .ZN(n5) );
  INV_X1 U279 ( .A(A[12]), .ZN(n192) );
  INV_X1 U280 ( .A(A[4]), .ZN(n278) );
  OAI221_X1 U281 ( .B1(n82), .B2(n279), .C1(n199), .C2(n184), .A(n201), .ZN(n4) );
  INV_X1 U282 ( .A(A[13]), .ZN(n184) );
  INV_X1 U283 ( .A(A[5]), .ZN(n279) );
  OAI211_X1 U284 ( .C1(n43), .C2(n56), .A(n280), .B(n281), .ZN(\output [0]) );
  AOI221_X1 U285 ( .B1(sel[0]), .B2(n282), .C1(n28), .C2(n38), .A(n283), .ZN(
        n281) );
  OAI22_X1 U286 ( .A1(n31), .A2(n57), .B1(n11), .B2(n284), .ZN(n283) );
  NAND2_X1 U287 ( .A1(sel[0]), .A2(n76), .ZN(n11) );
  NAND2_X1 U288 ( .A1(A[6]), .A2(sel[0]), .ZN(n57) );
  NAND3_X1 U289 ( .A1(B[1]), .A2(n285), .A3(n286), .ZN(n31) );
  OAI221_X1 U290 ( .B1(n82), .B2(n284), .C1(n199), .C2(n232), .A(n201), .ZN(
        n38) );
  NAND3_X1 U291 ( .A1(B[3]), .A2(n96), .A3(B[4]), .ZN(n201) );
  INV_X1 U292 ( .A(sel[1]), .ZN(n237) );
  INV_X1 U293 ( .A(A[31]), .ZN(n81) );
  INV_X1 U294 ( .A(A[8]), .ZN(n232) );
  OAI21_X1 U295 ( .B1(n235), .B2(n159), .A(sel[0]), .ZN(n199) );
  NOR2_X1 U296 ( .A1(n159), .A2(B[3]), .ZN(n235) );
  INV_X1 U297 ( .A(B[4]), .ZN(n159) );
  INV_X1 U298 ( .A(A[0]), .ZN(n284) );
  INV_X1 U299 ( .A(B[3]), .ZN(n160) );
  NOR3_X1 U300 ( .A1(sel[0]), .A2(sel[1]), .A3(B[4]), .ZN(n276) );
  NAND2_X1 U301 ( .A1(n76), .A2(n103), .ZN(n20) );
  NOR2_X1 U302 ( .A1(n287), .A2(B[0]), .ZN(n76) );
  OAI222_X1 U303 ( .A1(n27), .A2(n203), .B1(n8), .B2(n198), .C1(n202), .C2(n13), .ZN(n282) );
  INV_X1 U304 ( .A(n116), .ZN(n13) );
  XOR2_X1 U305 ( .A(n289), .B(sel[0]), .Z(n286) );
  INV_X1 U306 ( .A(A[2]), .ZN(n202) );
  INV_X1 U307 ( .A(A[1]), .ZN(n198) );
  INV_X1 U308 ( .A(n39), .ZN(n8) );
  NAND3_X1 U309 ( .A1(B[1]), .A2(n292), .A3(B[2]), .ZN(n291) );
  INV_X1 U310 ( .A(A[3]), .ZN(n203) );
  INV_X1 U311 ( .A(n6), .ZN(n27) );
  NAND3_X1 U312 ( .A1(B[1]), .A2(n289), .A3(n296), .ZN(n295) );
  AOI22_X1 U313 ( .A1(n54), .A2(n25), .B1(n61), .B2(n3), .ZN(n280) );
  INV_X1 U314 ( .A(n105), .ZN(n61) );
  NAND2_X1 U315 ( .A1(A[4]), .A2(sel[0]), .ZN(n105) );
  NAND3_X1 U316 ( .A1(n292), .A2(n289), .A3(B[1]), .ZN(n297) );
  NAND2_X1 U317 ( .A1(B[2]), .A2(n288), .ZN(n294) );
  INV_X1 U318 ( .A(n296), .ZN(n290) );
  INV_X1 U319 ( .A(n67), .ZN(n54) );
  NAND2_X1 U320 ( .A1(A[5]), .A2(sel[0]), .ZN(n67) );
  NAND2_X1 U321 ( .A1(A[7]), .A2(sel[0]), .ZN(n56) );
  INV_X1 U322 ( .A(n15), .ZN(n43) );
  NAND3_X1 U323 ( .A1(B[2]), .A2(B[1]), .A3(n296), .ZN(n298) );
  NOR2_X1 U324 ( .A1(n285), .A2(n103), .ZN(n296) );
  INV_X1 U325 ( .A(sel[0]), .ZN(n103) );
  INV_X1 U326 ( .A(n292), .ZN(n293) );
  NOR2_X1 U327 ( .A1(n285), .A2(sel[0]), .ZN(n292) );
  INV_X1 U328 ( .A(B[0]), .ZN(n285) );
  NAND2_X1 U329 ( .A1(n288), .A2(n289), .ZN(n287) );
  INV_X1 U330 ( .A(B[2]), .ZN(n289) );
  INV_X1 U331 ( .A(B[1]), .ZN(n288) );
endmodule


module ND3_N32_0 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;


  NAND3_X1 U1 ( .A1(B[9]), .A2(A[9]), .A3(S), .ZN(Y[9]) );
  NAND3_X1 U2 ( .A1(A[8]), .A2(S), .A3(B[8]), .ZN(Y[8]) );
  NAND3_X1 U3 ( .A1(A[7]), .A2(S), .A3(B[7]), .ZN(Y[7]) );
  NAND3_X1 U4 ( .A1(A[6]), .A2(S), .A3(B[6]), .ZN(Y[6]) );
  NAND3_X1 U5 ( .A1(A[5]), .A2(S), .A3(B[5]), .ZN(Y[5]) );
  NAND3_X1 U6 ( .A1(A[4]), .A2(S), .A3(B[4]), .ZN(Y[4]) );
  NAND3_X1 U7 ( .A1(A[3]), .A2(S), .A3(B[3]), .ZN(Y[3]) );
  NAND3_X1 U8 ( .A1(A[31]), .A2(S), .A3(B[31]), .ZN(Y[31]) );
  NAND3_X1 U9 ( .A1(A[30]), .A2(S), .A3(B[30]), .ZN(Y[30]) );
  NAND3_X1 U10 ( .A1(A[2]), .A2(S), .A3(B[2]), .ZN(Y[2]) );
  NAND3_X1 U11 ( .A1(A[29]), .A2(S), .A3(B[29]), .ZN(Y[29]) );
  NAND3_X1 U12 ( .A1(A[28]), .A2(S), .A3(B[28]), .ZN(Y[28]) );
  NAND3_X1 U13 ( .A1(A[27]), .A2(S), .A3(B[27]), .ZN(Y[27]) );
  NAND3_X1 U14 ( .A1(A[26]), .A2(S), .A3(B[26]), .ZN(Y[26]) );
  NAND3_X1 U15 ( .A1(A[25]), .A2(S), .A3(B[25]), .ZN(Y[25]) );
  NAND3_X1 U16 ( .A1(A[24]), .A2(S), .A3(B[24]), .ZN(Y[24]) );
  NAND3_X1 U17 ( .A1(A[23]), .A2(S), .A3(B[23]), .ZN(Y[23]) );
  NAND3_X1 U18 ( .A1(A[22]), .A2(S), .A3(B[22]), .ZN(Y[22]) );
  NAND3_X1 U19 ( .A1(A[21]), .A2(S), .A3(B[21]), .ZN(Y[21]) );
  NAND3_X1 U20 ( .A1(A[20]), .A2(S), .A3(B[20]), .ZN(Y[20]) );
  NAND3_X1 U21 ( .A1(A[1]), .A2(S), .A3(B[1]), .ZN(Y[1]) );
  NAND3_X1 U22 ( .A1(A[19]), .A2(S), .A3(B[19]), .ZN(Y[19]) );
  NAND3_X1 U23 ( .A1(A[18]), .A2(S), .A3(B[18]), .ZN(Y[18]) );
  NAND3_X1 U24 ( .A1(A[17]), .A2(S), .A3(B[17]), .ZN(Y[17]) );
  NAND3_X1 U25 ( .A1(A[16]), .A2(S), .A3(B[16]), .ZN(Y[16]) );
  NAND3_X1 U26 ( .A1(A[15]), .A2(S), .A3(B[15]), .ZN(Y[15]) );
  NAND3_X1 U27 ( .A1(A[14]), .A2(S), .A3(B[14]), .ZN(Y[14]) );
  NAND3_X1 U28 ( .A1(A[13]), .A2(S), .A3(B[13]), .ZN(Y[13]) );
  NAND3_X1 U29 ( .A1(A[12]), .A2(S), .A3(B[12]), .ZN(Y[12]) );
  NAND3_X1 U30 ( .A1(A[11]), .A2(S), .A3(B[11]), .ZN(Y[11]) );
  NAND3_X1 U31 ( .A1(A[10]), .A2(S), .A3(B[10]), .ZN(Y[10]) );
  NAND3_X1 U32 ( .A1(A[0]), .A2(S), .A3(B[0]), .ZN(Y[0]) );
endmodule


module ND3_N32_3 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;


  NAND3_X1 U1 ( .A1(B[9]), .A2(A[9]), .A3(S), .ZN(Y[9]) );
  NAND3_X1 U2 ( .A1(A[8]), .A2(S), .A3(B[8]), .ZN(Y[8]) );
  NAND3_X1 U3 ( .A1(A[7]), .A2(S), .A3(B[7]), .ZN(Y[7]) );
  NAND3_X1 U4 ( .A1(A[6]), .A2(S), .A3(B[6]), .ZN(Y[6]) );
  NAND3_X1 U5 ( .A1(A[5]), .A2(S), .A3(B[5]), .ZN(Y[5]) );
  NAND3_X1 U6 ( .A1(A[4]), .A2(S), .A3(B[4]), .ZN(Y[4]) );
  NAND3_X1 U7 ( .A1(A[3]), .A2(S), .A3(B[3]), .ZN(Y[3]) );
  NAND3_X1 U8 ( .A1(A[31]), .A2(S), .A3(B[31]), .ZN(Y[31]) );
  NAND3_X1 U9 ( .A1(A[30]), .A2(S), .A3(B[30]), .ZN(Y[30]) );
  NAND3_X1 U10 ( .A1(A[2]), .A2(S), .A3(B[2]), .ZN(Y[2]) );
  NAND3_X1 U11 ( .A1(A[29]), .A2(S), .A3(B[29]), .ZN(Y[29]) );
  NAND3_X1 U12 ( .A1(A[28]), .A2(S), .A3(B[28]), .ZN(Y[28]) );
  NAND3_X1 U13 ( .A1(A[27]), .A2(S), .A3(B[27]), .ZN(Y[27]) );
  NAND3_X1 U14 ( .A1(A[26]), .A2(S), .A3(B[26]), .ZN(Y[26]) );
  NAND3_X1 U15 ( .A1(A[25]), .A2(S), .A3(B[25]), .ZN(Y[25]) );
  NAND3_X1 U16 ( .A1(A[24]), .A2(S), .A3(B[24]), .ZN(Y[24]) );
  NAND3_X1 U17 ( .A1(A[23]), .A2(S), .A3(B[23]), .ZN(Y[23]) );
  NAND3_X1 U18 ( .A1(A[22]), .A2(S), .A3(B[22]), .ZN(Y[22]) );
  NAND3_X1 U19 ( .A1(A[21]), .A2(S), .A3(B[21]), .ZN(Y[21]) );
  NAND3_X1 U20 ( .A1(A[20]), .A2(S), .A3(B[20]), .ZN(Y[20]) );
  NAND3_X1 U21 ( .A1(A[1]), .A2(S), .A3(B[1]), .ZN(Y[1]) );
  NAND3_X1 U22 ( .A1(A[19]), .A2(S), .A3(B[19]), .ZN(Y[19]) );
  NAND3_X1 U23 ( .A1(A[18]), .A2(S), .A3(B[18]), .ZN(Y[18]) );
  NAND3_X1 U24 ( .A1(A[17]), .A2(S), .A3(B[17]), .ZN(Y[17]) );
  NAND3_X1 U25 ( .A1(A[16]), .A2(S), .A3(B[16]), .ZN(Y[16]) );
  NAND3_X1 U26 ( .A1(A[15]), .A2(S), .A3(B[15]), .ZN(Y[15]) );
  NAND3_X1 U27 ( .A1(A[14]), .A2(S), .A3(B[14]), .ZN(Y[14]) );
  NAND3_X1 U28 ( .A1(A[13]), .A2(S), .A3(B[13]), .ZN(Y[13]) );
  NAND3_X1 U29 ( .A1(A[12]), .A2(S), .A3(B[12]), .ZN(Y[12]) );
  NAND3_X1 U30 ( .A1(A[11]), .A2(S), .A3(B[11]), .ZN(Y[11]) );
  NAND3_X1 U31 ( .A1(A[10]), .A2(S), .A3(B[10]), .ZN(Y[10]) );
  NAND3_X1 U32 ( .A1(A[0]), .A2(S), .A3(B[0]), .ZN(Y[0]) );
endmodule


module ND3_N32_2 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;


  NAND3_X1 U1 ( .A1(B[9]), .A2(A[9]), .A3(S), .ZN(Y[9]) );
  NAND3_X1 U2 ( .A1(A[8]), .A2(S), .A3(B[8]), .ZN(Y[8]) );
  NAND3_X1 U3 ( .A1(A[7]), .A2(S), .A3(B[7]), .ZN(Y[7]) );
  NAND3_X1 U4 ( .A1(A[6]), .A2(S), .A3(B[6]), .ZN(Y[6]) );
  NAND3_X1 U5 ( .A1(A[5]), .A2(S), .A3(B[5]), .ZN(Y[5]) );
  NAND3_X1 U6 ( .A1(A[4]), .A2(S), .A3(B[4]), .ZN(Y[4]) );
  NAND3_X1 U7 ( .A1(A[3]), .A2(S), .A3(B[3]), .ZN(Y[3]) );
  NAND3_X1 U8 ( .A1(A[31]), .A2(S), .A3(B[31]), .ZN(Y[31]) );
  NAND3_X1 U9 ( .A1(A[30]), .A2(S), .A3(B[30]), .ZN(Y[30]) );
  NAND3_X1 U10 ( .A1(A[2]), .A2(S), .A3(B[2]), .ZN(Y[2]) );
  NAND3_X1 U11 ( .A1(A[29]), .A2(S), .A3(B[29]), .ZN(Y[29]) );
  NAND3_X1 U12 ( .A1(A[28]), .A2(S), .A3(B[28]), .ZN(Y[28]) );
  NAND3_X1 U13 ( .A1(A[27]), .A2(S), .A3(B[27]), .ZN(Y[27]) );
  NAND3_X1 U14 ( .A1(A[26]), .A2(S), .A3(B[26]), .ZN(Y[26]) );
  NAND3_X1 U15 ( .A1(A[25]), .A2(S), .A3(B[25]), .ZN(Y[25]) );
  NAND3_X1 U16 ( .A1(A[24]), .A2(S), .A3(B[24]), .ZN(Y[24]) );
  NAND3_X1 U17 ( .A1(A[23]), .A2(S), .A3(B[23]), .ZN(Y[23]) );
  NAND3_X1 U18 ( .A1(A[22]), .A2(S), .A3(B[22]), .ZN(Y[22]) );
  NAND3_X1 U19 ( .A1(A[21]), .A2(S), .A3(B[21]), .ZN(Y[21]) );
  NAND3_X1 U20 ( .A1(A[20]), .A2(S), .A3(B[20]), .ZN(Y[20]) );
  NAND3_X1 U21 ( .A1(A[1]), .A2(S), .A3(B[1]), .ZN(Y[1]) );
  NAND3_X1 U22 ( .A1(A[19]), .A2(S), .A3(B[19]), .ZN(Y[19]) );
  NAND3_X1 U23 ( .A1(A[18]), .A2(S), .A3(B[18]), .ZN(Y[18]) );
  NAND3_X1 U24 ( .A1(A[17]), .A2(S), .A3(B[17]), .ZN(Y[17]) );
  NAND3_X1 U25 ( .A1(A[16]), .A2(S), .A3(B[16]), .ZN(Y[16]) );
  NAND3_X1 U26 ( .A1(A[15]), .A2(S), .A3(B[15]), .ZN(Y[15]) );
  NAND3_X1 U27 ( .A1(A[14]), .A2(S), .A3(B[14]), .ZN(Y[14]) );
  NAND3_X1 U28 ( .A1(A[13]), .A2(S), .A3(B[13]), .ZN(Y[13]) );
  NAND3_X1 U29 ( .A1(A[12]), .A2(S), .A3(B[12]), .ZN(Y[12]) );
  NAND3_X1 U30 ( .A1(A[11]), .A2(S), .A3(B[11]), .ZN(Y[11]) );
  NAND3_X1 U31 ( .A1(A[10]), .A2(S), .A3(B[10]), .ZN(Y[10]) );
  NAND3_X1 U32 ( .A1(A[0]), .A2(S), .A3(B[0]), .ZN(Y[0]) );
endmodule


module ND3_N32_1 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;


  NAND3_X1 U1 ( .A1(B[9]), .A2(A[9]), .A3(S), .ZN(Y[9]) );
  NAND3_X1 U2 ( .A1(A[8]), .A2(S), .A3(B[8]), .ZN(Y[8]) );
  NAND3_X1 U3 ( .A1(A[7]), .A2(S), .A3(B[7]), .ZN(Y[7]) );
  NAND3_X1 U4 ( .A1(A[6]), .A2(S), .A3(B[6]), .ZN(Y[6]) );
  NAND3_X1 U5 ( .A1(A[5]), .A2(S), .A3(B[5]), .ZN(Y[5]) );
  NAND3_X1 U6 ( .A1(A[4]), .A2(S), .A3(B[4]), .ZN(Y[4]) );
  NAND3_X1 U7 ( .A1(A[3]), .A2(S), .A3(B[3]), .ZN(Y[3]) );
  NAND3_X1 U8 ( .A1(A[31]), .A2(S), .A3(B[31]), .ZN(Y[31]) );
  NAND3_X1 U9 ( .A1(A[30]), .A2(S), .A3(B[30]), .ZN(Y[30]) );
  NAND3_X1 U10 ( .A1(A[2]), .A2(S), .A3(B[2]), .ZN(Y[2]) );
  NAND3_X1 U11 ( .A1(A[29]), .A2(S), .A3(B[29]), .ZN(Y[29]) );
  NAND3_X1 U12 ( .A1(A[28]), .A2(S), .A3(B[28]), .ZN(Y[28]) );
  NAND3_X1 U13 ( .A1(A[27]), .A2(S), .A3(B[27]), .ZN(Y[27]) );
  NAND3_X1 U14 ( .A1(A[26]), .A2(S), .A3(B[26]), .ZN(Y[26]) );
  NAND3_X1 U15 ( .A1(A[25]), .A2(S), .A3(B[25]), .ZN(Y[25]) );
  NAND3_X1 U16 ( .A1(A[24]), .A2(S), .A3(B[24]), .ZN(Y[24]) );
  NAND3_X1 U17 ( .A1(A[23]), .A2(S), .A3(B[23]), .ZN(Y[23]) );
  NAND3_X1 U18 ( .A1(A[22]), .A2(S), .A3(B[22]), .ZN(Y[22]) );
  NAND3_X1 U19 ( .A1(A[21]), .A2(S), .A3(B[21]), .ZN(Y[21]) );
  NAND3_X1 U20 ( .A1(A[20]), .A2(S), .A3(B[20]), .ZN(Y[20]) );
  NAND3_X1 U21 ( .A1(A[1]), .A2(S), .A3(B[1]), .ZN(Y[1]) );
  NAND3_X1 U22 ( .A1(A[19]), .A2(S), .A3(B[19]), .ZN(Y[19]) );
  NAND3_X1 U23 ( .A1(A[18]), .A2(S), .A3(B[18]), .ZN(Y[18]) );
  NAND3_X1 U24 ( .A1(A[17]), .A2(S), .A3(B[17]), .ZN(Y[17]) );
  NAND3_X1 U25 ( .A1(A[16]), .A2(S), .A3(B[16]), .ZN(Y[16]) );
  NAND3_X1 U26 ( .A1(A[15]), .A2(S), .A3(B[15]), .ZN(Y[15]) );
  NAND3_X1 U27 ( .A1(A[14]), .A2(S), .A3(B[14]), .ZN(Y[14]) );
  NAND3_X1 U28 ( .A1(A[13]), .A2(S), .A3(B[13]), .ZN(Y[13]) );
  NAND3_X1 U29 ( .A1(A[12]), .A2(S), .A3(B[12]), .ZN(Y[12]) );
  NAND3_X1 U30 ( .A1(A[11]), .A2(S), .A3(B[11]), .ZN(Y[11]) );
  NAND3_X1 U31 ( .A1(A[10]), .A2(S), .A3(B[10]), .ZN(Y[10]) );
  NAND3_X1 U32 ( .A1(A[0]), .A2(S), .A3(B[0]), .ZN(Y[0]) );
endmodule


module ND4_N32 ( L0, L1, L2, L3, Y );
  input [31:0] L0;
  input [31:0] L1;
  input [31:0] L2;
  input [31:0] L3;
  output [31:0] Y;


  NAND4_X1 U1 ( .A1(L3[9]), .A2(L2[9]), .A3(L1[9]), .A4(L0[9]), .ZN(Y[9]) );
  NAND4_X1 U2 ( .A1(L3[8]), .A2(L2[8]), .A3(L1[8]), .A4(L0[8]), .ZN(Y[8]) );
  NAND4_X1 U3 ( .A1(L3[7]), .A2(L2[7]), .A3(L1[7]), .A4(L0[7]), .ZN(Y[7]) );
  NAND4_X1 U4 ( .A1(L3[6]), .A2(L2[6]), .A3(L1[6]), .A4(L0[6]), .ZN(Y[6]) );
  NAND4_X1 U5 ( .A1(L3[5]), .A2(L2[5]), .A3(L1[5]), .A4(L0[5]), .ZN(Y[5]) );
  NAND4_X1 U6 ( .A1(L3[4]), .A2(L2[4]), .A3(L1[4]), .A4(L0[4]), .ZN(Y[4]) );
  NAND4_X1 U7 ( .A1(L3[3]), .A2(L2[3]), .A3(L1[3]), .A4(L0[3]), .ZN(Y[3]) );
  NAND4_X1 U8 ( .A1(L3[31]), .A2(L2[31]), .A3(L1[31]), .A4(L0[31]), .ZN(Y[31])
         );
  NAND4_X1 U9 ( .A1(L3[30]), .A2(L2[30]), .A3(L1[30]), .A4(L0[30]), .ZN(Y[30])
         );
  NAND4_X1 U10 ( .A1(L3[2]), .A2(L2[2]), .A3(L1[2]), .A4(L0[2]), .ZN(Y[2]) );
  NAND4_X1 U11 ( .A1(L3[29]), .A2(L2[29]), .A3(L1[29]), .A4(L0[29]), .ZN(Y[29]) );
  NAND4_X1 U12 ( .A1(L3[28]), .A2(L2[28]), .A3(L1[28]), .A4(L0[28]), .ZN(Y[28]) );
  NAND4_X1 U13 ( .A1(L3[27]), .A2(L2[27]), .A3(L1[27]), .A4(L0[27]), .ZN(Y[27]) );
  NAND4_X1 U14 ( .A1(L3[26]), .A2(L2[26]), .A3(L1[26]), .A4(L0[26]), .ZN(Y[26]) );
  NAND4_X1 U15 ( .A1(L3[25]), .A2(L2[25]), .A3(L1[25]), .A4(L0[25]), .ZN(Y[25]) );
  NAND4_X1 U16 ( .A1(L3[24]), .A2(L2[24]), .A3(L1[24]), .A4(L0[24]), .ZN(Y[24]) );
  NAND4_X1 U17 ( .A1(L3[23]), .A2(L2[23]), .A3(L1[23]), .A4(L0[23]), .ZN(Y[23]) );
  NAND4_X1 U18 ( .A1(L3[22]), .A2(L2[22]), .A3(L1[22]), .A4(L0[22]), .ZN(Y[22]) );
  NAND4_X1 U19 ( .A1(L3[21]), .A2(L2[21]), .A3(L1[21]), .A4(L0[21]), .ZN(Y[21]) );
  NAND4_X1 U20 ( .A1(L3[20]), .A2(L2[20]), .A3(L1[20]), .A4(L0[20]), .ZN(Y[20]) );
  NAND4_X1 U21 ( .A1(L3[1]), .A2(L2[1]), .A3(L1[1]), .A4(L0[1]), .ZN(Y[1]) );
  NAND4_X1 U22 ( .A1(L3[19]), .A2(L2[19]), .A3(L1[19]), .A4(L0[19]), .ZN(Y[19]) );
  NAND4_X1 U23 ( .A1(L3[18]), .A2(L2[18]), .A3(L1[18]), .A4(L0[18]), .ZN(Y[18]) );
  NAND4_X1 U24 ( .A1(L3[17]), .A2(L2[17]), .A3(L1[17]), .A4(L0[17]), .ZN(Y[17]) );
  NAND4_X1 U25 ( .A1(L3[16]), .A2(L2[16]), .A3(L1[16]), .A4(L0[16]), .ZN(Y[16]) );
  NAND4_X1 U26 ( .A1(L3[15]), .A2(L2[15]), .A3(L1[15]), .A4(L0[15]), .ZN(Y[15]) );
  NAND4_X1 U27 ( .A1(L3[14]), .A2(L2[14]), .A3(L1[14]), .A4(L0[14]), .ZN(Y[14]) );
  NAND4_X1 U28 ( .A1(L3[13]), .A2(L2[13]), .A3(L1[13]), .A4(L0[13]), .ZN(Y[13]) );
  NAND4_X1 U29 ( .A1(L3[12]), .A2(L2[12]), .A3(L1[12]), .A4(L0[12]), .ZN(Y[12]) );
  NAND4_X1 U30 ( .A1(L3[11]), .A2(L2[11]), .A3(L1[11]), .A4(L0[11]), .ZN(Y[11]) );
  NAND4_X1 U31 ( .A1(L3[10]), .A2(L2[10]), .A3(L1[10]), .A4(L0[10]), .ZN(Y[10]) );
  NAND4_X1 U32 ( .A1(L3[0]), .A2(L2[0]), .A3(L1[0]), .A4(L0[0]), .ZN(Y[0]) );
endmodule


module LogicalT2_N32 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [3:0] S;
  output [31:0] Y;
  wire   \L[0][31] , \L[0][30] , \L[0][29] , \L[0][28] , \L[0][27] ,
         \L[0][26] , \L[0][25] , \L[0][24] , \L[0][23] , \L[0][22] ,
         \L[0][21] , \L[0][20] , \L[0][19] , \L[0][18] , \L[0][17] ,
         \L[0][16] , \L[0][15] , \L[0][14] , \L[0][13] , \L[0][12] ,
         \L[0][11] , \L[0][10] , \L[0][9] , \L[0][8] , \L[0][7] , \L[0][6] ,
         \L[0][5] , \L[0][4] , \L[0][3] , \L[0][2] , \L[0][1] , \L[0][0] ,
         \L[1][31] , \L[1][30] , \L[1][29] , \L[1][28] , \L[1][27] ,
         \L[1][26] , \L[1][25] , \L[1][24] , \L[1][23] , \L[1][22] ,
         \L[1][21] , \L[1][20] , \L[1][19] , \L[1][18] , \L[1][17] ,
         \L[1][16] , \L[1][15] , \L[1][14] , \L[1][13] , \L[1][12] ,
         \L[1][11] , \L[1][10] , \L[1][9] , \L[1][8] , \L[1][7] , \L[1][6] ,
         \L[1][5] , \L[1][4] , \L[1][3] , \L[1][2] , \L[1][1] , \L[1][0] ,
         \L[2][31] , \L[2][30] , \L[2][29] , \L[2][28] , \L[2][27] ,
         \L[2][26] , \L[2][25] , \L[2][24] , \L[2][23] , \L[2][22] ,
         \L[2][21] , \L[2][20] , \L[2][19] , \L[2][18] , \L[2][17] ,
         \L[2][16] , \L[2][15] , \L[2][14] , \L[2][13] , \L[2][12] ,
         \L[2][11] , \L[2][10] , \L[2][9] , \L[2][8] , \L[2][7] , \L[2][6] ,
         \L[2][5] , \L[2][4] , \L[2][3] , \L[2][2] , \L[2][1] , \L[2][0] ,
         \L[3][31] , \L[3][30] , \L[3][29] , \L[3][28] , \L[3][27] ,
         \L[3][26] , \L[3][25] , \L[3][24] , \L[3][23] , \L[3][22] ,
         \L[3][21] , \L[3][20] , \L[3][19] , \L[3][18] , \L[3][17] ,
         \L[3][16] , \L[3][15] , \L[3][14] , \L[3][13] , \L[3][12] ,
         \L[3][11] , \L[3][10] , \L[3][9] , \L[3][8] , \L[3][7] , \L[3][6] ,
         \L[3][5] , \L[3][4] , \L[3][3] , \L[3][2] , \L[3][1] , \L[3][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;

  ND3_N32_0 nand0 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, 
        n6, n5, n4, n3, n2, n1}), .B({n64, n63, n62, n61, n60, n59, n58, n57, 
        n56, n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, 
        n42, n41, n40, n39, n38, n37, n36, n35, n34, n33}), .S(S[3]), .Y({
        \L[0][31] , \L[0][30] , \L[0][29] , \L[0][28] , \L[0][27] , \L[0][26] , 
        \L[0][25] , \L[0][24] , \L[0][23] , \L[0][22] , \L[0][21] , \L[0][20] , 
        \L[0][19] , \L[0][18] , \L[0][17] , \L[0][16] , \L[0][15] , \L[0][14] , 
        \L[0][13] , \L[0][12] , \L[0][11] , \L[0][10] , \L[0][9] , \L[0][8] , 
        \L[0][7] , \L[0][6] , \L[0][5] , \L[0][4] , \L[0][3] , \L[0][2] , 
        \L[0][1] , \L[0][0] }) );
  ND3_N32_3 nand1 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, 
        n6, n5, n4, n3, n2, n1}), .B(B), .S(S[2]), .Y({\L[1][31] , \L[1][30] , 
        \L[1][29] , \L[1][28] , \L[1][27] , \L[1][26] , \L[1][25] , \L[1][24] , 
        \L[1][23] , \L[1][22] , \L[1][21] , \L[1][20] , \L[1][19] , \L[1][18] , 
        \L[1][17] , \L[1][16] , \L[1][15] , \L[1][14] , \L[1][13] , \L[1][12] , 
        \L[1][11] , \L[1][10] , \L[1][9] , \L[1][8] , \L[1][7] , \L[1][6] , 
        \L[1][5] , \L[1][4] , \L[1][3] , \L[1][2] , \L[1][1] , \L[1][0] }) );
  ND3_N32_2 nand2 ( .A(A), .B({n64, n63, n62, n61, n60, n59, n58, n57, n56, 
        n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, n42, 
        n41, n40, n39, n38, n37, n36, n35, n34, n33}), .S(S[1]), .Y({
        \L[2][31] , \L[2][30] , \L[2][29] , \L[2][28] , \L[2][27] , \L[2][26] , 
        \L[2][25] , \L[2][24] , \L[2][23] , \L[2][22] , \L[2][21] , \L[2][20] , 
        \L[2][19] , \L[2][18] , \L[2][17] , \L[2][16] , \L[2][15] , \L[2][14] , 
        \L[2][13] , \L[2][12] , \L[2][11] , \L[2][10] , \L[2][9] , \L[2][8] , 
        \L[2][7] , \L[2][6] , \L[2][5] , \L[2][4] , \L[2][3] , \L[2][2] , 
        \L[2][1] , \L[2][0] }) );
  ND3_N32_1 nand3 ( .A(A), .B(B), .S(S[0]), .Y({\L[3][31] , \L[3][30] , 
        \L[3][29] , \L[3][28] , \L[3][27] , \L[3][26] , \L[3][25] , \L[3][24] , 
        \L[3][23] , \L[3][22] , \L[3][21] , \L[3][20] , \L[3][19] , \L[3][18] , 
        \L[3][17] , \L[3][16] , \L[3][15] , \L[3][14] , \L[3][13] , \L[3][12] , 
        \L[3][11] , \L[3][10] , \L[3][9] , \L[3][8] , \L[3][7] , \L[3][6] , 
        \L[3][5] , \L[3][4] , \L[3][3] , \L[3][2] , \L[3][1] , \L[3][0] }) );
  ND4_N32 level2 ( .L0({\L[0][31] , \L[0][30] , \L[0][29] , \L[0][28] , 
        \L[0][27] , \L[0][26] , \L[0][25] , \L[0][24] , \L[0][23] , \L[0][22] , 
        \L[0][21] , \L[0][20] , \L[0][19] , \L[0][18] , \L[0][17] , \L[0][16] , 
        \L[0][15] , \L[0][14] , \L[0][13] , \L[0][12] , \L[0][11] , \L[0][10] , 
        \L[0][9] , \L[0][8] , \L[0][7] , \L[0][6] , \L[0][5] , \L[0][4] , 
        \L[0][3] , \L[0][2] , \L[0][1] , \L[0][0] }), .L1({\L[1][31] , 
        \L[1][30] , \L[1][29] , \L[1][28] , \L[1][27] , \L[1][26] , \L[1][25] , 
        \L[1][24] , \L[1][23] , \L[1][22] , \L[1][21] , \L[1][20] , \L[1][19] , 
        \L[1][18] , \L[1][17] , \L[1][16] , \L[1][15] , \L[1][14] , \L[1][13] , 
        \L[1][12] , \L[1][11] , \L[1][10] , \L[1][9] , \L[1][8] , \L[1][7] , 
        \L[1][6] , \L[1][5] , \L[1][4] , \L[1][3] , \L[1][2] , \L[1][1] , 
        \L[1][0] }), .L2({\L[2][31] , \L[2][30] , \L[2][29] , \L[2][28] , 
        \L[2][27] , \L[2][26] , \L[2][25] , \L[2][24] , \L[2][23] , \L[2][22] , 
        \L[2][21] , \L[2][20] , \L[2][19] , \L[2][18] , \L[2][17] , \L[2][16] , 
        \L[2][15] , \L[2][14] , \L[2][13] , \L[2][12] , \L[2][11] , \L[2][10] , 
        \L[2][9] , \L[2][8] , \L[2][7] , \L[2][6] , \L[2][5] , \L[2][4] , 
        \L[2][3] , \L[2][2] , \L[2][1] , \L[2][0] }), .L3({\L[3][31] , 
        \L[3][30] , \L[3][29] , \L[3][28] , \L[3][27] , \L[3][26] , \L[3][25] , 
        \L[3][24] , \L[3][23] , \L[3][22] , \L[3][21] , \L[3][20] , \L[3][19] , 
        \L[3][18] , \L[3][17] , \L[3][16] , \L[3][15] , \L[3][14] , \L[3][13] , 
        \L[3][12] , \L[3][11] , \L[3][10] , \L[3][9] , \L[3][8] , \L[3][7] , 
        \L[3][6] , \L[3][5] , \L[3][4] , \L[3][3] , \L[3][2] , \L[3][1] , 
        \L[3][0] }), .Y(Y) );
  INV_X1 U1 ( .A(A[0]), .ZN(n1) );
  INV_X1 U2 ( .A(A[1]), .ZN(n2) );
  INV_X1 U3 ( .A(A[2]), .ZN(n3) );
  INV_X1 U4 ( .A(A[3]), .ZN(n4) );
  INV_X1 U5 ( .A(A[4]), .ZN(n5) );
  INV_X1 U6 ( .A(A[5]), .ZN(n6) );
  INV_X1 U7 ( .A(A[6]), .ZN(n7) );
  INV_X1 U8 ( .A(A[7]), .ZN(n8) );
  INV_X1 U9 ( .A(A[8]), .ZN(n9) );
  INV_X1 U10 ( .A(A[9]), .ZN(n10) );
  INV_X1 U11 ( .A(A[10]), .ZN(n11) );
  INV_X1 U12 ( .A(A[11]), .ZN(n12) );
  INV_X1 U13 ( .A(A[12]), .ZN(n13) );
  INV_X1 U14 ( .A(A[13]), .ZN(n14) );
  INV_X1 U15 ( .A(A[14]), .ZN(n15) );
  INV_X1 U16 ( .A(A[15]), .ZN(n16) );
  INV_X1 U17 ( .A(A[16]), .ZN(n17) );
  INV_X1 U18 ( .A(A[17]), .ZN(n18) );
  INV_X1 U19 ( .A(A[18]), .ZN(n19) );
  INV_X1 U20 ( .A(A[19]), .ZN(n20) );
  INV_X1 U21 ( .A(A[20]), .ZN(n21) );
  INV_X1 U22 ( .A(A[21]), .ZN(n22) );
  INV_X1 U23 ( .A(A[22]), .ZN(n23) );
  INV_X1 U24 ( .A(A[23]), .ZN(n24) );
  INV_X1 U25 ( .A(A[24]), .ZN(n25) );
  INV_X1 U26 ( .A(A[25]), .ZN(n26) );
  INV_X1 U27 ( .A(A[26]), .ZN(n27) );
  INV_X1 U28 ( .A(A[27]), .ZN(n28) );
  INV_X1 U29 ( .A(A[28]), .ZN(n29) );
  INV_X1 U30 ( .A(A[29]), .ZN(n30) );
  INV_X1 U31 ( .A(A[30]), .ZN(n31) );
  INV_X1 U32 ( .A(A[31]), .ZN(n32) );
  INV_X1 U33 ( .A(B[0]), .ZN(n33) );
  INV_X1 U34 ( .A(B[1]), .ZN(n34) );
  INV_X1 U35 ( .A(B[2]), .ZN(n35) );
  INV_X1 U36 ( .A(B[3]), .ZN(n36) );
  INV_X1 U37 ( .A(B[4]), .ZN(n37) );
  INV_X1 U38 ( .A(B[5]), .ZN(n38) );
  INV_X1 U39 ( .A(B[6]), .ZN(n39) );
  INV_X1 U40 ( .A(B[7]), .ZN(n40) );
  INV_X1 U41 ( .A(B[8]), .ZN(n41) );
  INV_X1 U42 ( .A(B[9]), .ZN(n42) );
  INV_X1 U43 ( .A(B[10]), .ZN(n43) );
  INV_X1 U44 ( .A(B[11]), .ZN(n44) );
  INV_X1 U45 ( .A(B[12]), .ZN(n45) );
  INV_X1 U46 ( .A(B[13]), .ZN(n46) );
  INV_X1 U47 ( .A(B[14]), .ZN(n47) );
  INV_X1 U48 ( .A(B[15]), .ZN(n48) );
  INV_X1 U49 ( .A(B[16]), .ZN(n49) );
  INV_X1 U50 ( .A(B[17]), .ZN(n50) );
  INV_X1 U51 ( .A(B[18]), .ZN(n51) );
  INV_X1 U52 ( .A(B[19]), .ZN(n52) );
  INV_X1 U53 ( .A(B[20]), .ZN(n53) );
  INV_X1 U54 ( .A(B[21]), .ZN(n54) );
  INV_X1 U55 ( .A(B[22]), .ZN(n55) );
  INV_X1 U56 ( .A(B[23]), .ZN(n56) );
  INV_X1 U57 ( .A(B[24]), .ZN(n57) );
  INV_X1 U58 ( .A(B[25]), .ZN(n58) );
  INV_X1 U59 ( .A(B[26]), .ZN(n59) );
  INV_X1 U60 ( .A(B[27]), .ZN(n60) );
  INV_X1 U61 ( .A(B[28]), .ZN(n61) );
  INV_X1 U62 ( .A(B[29]), .ZN(n62) );
  INV_X1 U63 ( .A(B[30]), .ZN(n63) );
  INV_X1 U64 ( .A(B[31]), .ZN(n64) );
endmodule


module NOR2_0 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_15 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_14 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_13 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_12 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_11 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_10 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_9 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_8 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_7 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_6 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_5 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_4 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_3 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_2 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR2_1 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_15 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_14 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_13 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_12 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_11 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_10 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_9 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_8 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_7 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_6 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_5 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_4 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_3 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_2 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND2_1 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NORN_N32 ( A, Z );
  input [31:0] A;
  output Z;
  wire   \M[3][1] , \M[3][0] , \M[2][3] , \M[2][2] , \M[2][1] , \M[2][0] ,
         \M[1][7] , \M[1][6] , \M[1][5] , \M[1][4] , \M[1][3] , \M[1][2] ,
         \M[1][1] , \M[1][0] , \M[0][15] , \M[0][14] , \M[0][13] , \M[0][12] ,
         \M[0][11] , \M[0][10] , \M[0][9] , \M[0][8] , \M[0][7] , \M[0][6] ,
         \M[0][5] , \M[0][4] , \M[0][3] , \M[0][2] , \M[0][1] , \M[0][0] ;

  NOR2_0 NOR0i_0_0 ( .A(A[0]), .B(A[1]), .Y(\M[0][0] ) );
  NOR2_15 NOR0i_0_1 ( .A(A[2]), .B(A[3]), .Y(\M[0][1] ) );
  NOR2_14 NOR0i_0_2 ( .A(A[4]), .B(A[5]), .Y(\M[0][2] ) );
  NOR2_13 NOR0i_0_3 ( .A(A[6]), .B(A[7]), .Y(\M[0][3] ) );
  NOR2_12 NOR0i_0_4 ( .A(A[8]), .B(A[9]), .Y(\M[0][4] ) );
  NOR2_11 NOR0i_0_5 ( .A(A[10]), .B(A[11]), .Y(\M[0][5] ) );
  NOR2_10 NOR0i_0_6 ( .A(A[12]), .B(A[13]), .Y(\M[0][6] ) );
  NOR2_9 NOR0i_0_7 ( .A(A[14]), .B(A[15]), .Y(\M[0][7] ) );
  NOR2_8 NOR0i_0_8 ( .A(A[16]), .B(A[17]), .Y(\M[0][8] ) );
  NOR2_7 NOR0i_0_9 ( .A(A[18]), .B(A[19]), .Y(\M[0][9] ) );
  NOR2_6 NOR0i_0_10 ( .A(A[20]), .B(A[21]), .Y(\M[0][10] ) );
  NOR2_5 NOR0i_0_11 ( .A(A[22]), .B(A[23]), .Y(\M[0][11] ) );
  NOR2_4 NOR0i_0_12 ( .A(A[24]), .B(A[25]), .Y(\M[0][12] ) );
  NOR2_3 NOR0i_0_13 ( .A(A[26]), .B(A[27]), .Y(\M[0][13] ) );
  NOR2_2 NOR0i_0_14 ( .A(A[28]), .B(A[29]), .Y(\M[0][14] ) );
  NOR2_1 NOR0i_0_15 ( .A(A[30]), .B(A[31]), .Y(\M[0][15] ) );
  AND2_15 ANDi_1_0 ( .A(\M[0][0] ), .B(\M[0][1] ), .Y(\M[1][0] ) );
  AND2_14 ANDi_1_1 ( .A(\M[0][2] ), .B(\M[0][3] ), .Y(\M[1][1] ) );
  AND2_13 ANDi_1_2 ( .A(\M[0][4] ), .B(\M[0][5] ), .Y(\M[1][2] ) );
  AND2_12 ANDi_1_3 ( .A(\M[0][6] ), .B(\M[0][7] ), .Y(\M[1][3] ) );
  AND2_11 ANDi_1_4 ( .A(\M[0][8] ), .B(\M[0][9] ), .Y(\M[1][4] ) );
  AND2_10 ANDi_1_5 ( .A(\M[0][10] ), .B(\M[0][11] ), .Y(\M[1][5] ) );
  AND2_9 ANDi_1_6 ( .A(\M[0][12] ), .B(\M[0][13] ), .Y(\M[1][6] ) );
  AND2_8 ANDi_1_7 ( .A(\M[0][14] ), .B(\M[0][15] ), .Y(\M[1][7] ) );
  AND2_7 ANDi_2_0 ( .A(\M[1][0] ), .B(\M[1][1] ), .Y(\M[2][0] ) );
  AND2_6 ANDi_2_1 ( .A(\M[1][2] ), .B(\M[1][3] ), .Y(\M[2][1] ) );
  AND2_5 ANDi_2_2 ( .A(\M[1][4] ), .B(\M[1][5] ), .Y(\M[2][2] ) );
  AND2_4 ANDi_2_3 ( .A(\M[1][6] ), .B(\M[1][7] ), .Y(\M[2][3] ) );
  AND2_3 ANDi_3_0 ( .A(\M[2][0] ), .B(\M[2][1] ), .Y(\M[3][0] ) );
  AND2_2 ANDi_3_1 ( .A(\M[2][2] ), .B(\M[2][3] ), .Y(\M[3][1] ) );
  AND2_1 ANDi_4_0 ( .A(\M[3][0] ), .B(\M[3][1] ), .Y(Z) );
endmodule


module comparator ( C, Z, result );
  output [5:0] result;
  input C, Z;
  wire   C, Z;
  assign result[2] = C;
  assign result[1] = Z;

  INV_X1 U1 ( .A(result[5]), .ZN(result[3]) );
  NAND2_X1 U2 ( .A1(C), .A2(result[0]), .ZN(result[5]) );
  INV_X1 U3 ( .A(Z), .ZN(result[0]) );
  INV_X1 U4 ( .A(C), .ZN(result[4]) );
endmodule


module MUX6_1 ( NEQ_LINE, EQ_LINE, GEQ_LINE, G_LINE, L_LINE, LEQ_LINE, SEL, 
        RES_LINE );
  input [2:0] SEL;
  input NEQ_LINE, EQ_LINE, GEQ_LINE, G_LINE, L_LINE, LEQ_LINE;
  output RES_LINE;
  wire   n1, n2, n3, n4, n5;

  MUX2_X1 U1 ( .A(n1), .B(n2), .S(SEL[2]), .Z(RES_LINE) );
  MUX2_X1 U2 ( .A(LEQ_LINE), .B(L_LINE), .S(n3), .Z(n2) );
  NOR2_X1 U3 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n3) );
  MUX2_X1 U4 ( .A(n4), .B(n5), .S(SEL[1]), .Z(n1) );
  MUX2_X1 U5 ( .A(GEQ_LINE), .B(G_LINE), .S(SEL[0]), .Z(n5) );
  MUX2_X1 U6 ( .A(NEQ_LINE), .B(EQ_LINE), .S(SEL[0]), .Z(n4) );
endmodule


module topLevelCMP_N32 ( SUB, Cout, Sel, res );
  input [31:0] SUB;
  input [2:0] Sel;
  output [31:0] res;
  input Cout;
  wire   Z_s;
  wire   [5:0] cmp_res_6bit;
  assign res[1] = 1'b0;
  assign res[2] = 1'b0;
  assign res[3] = 1'b0;
  assign res[4] = 1'b0;
  assign res[5] = 1'b0;
  assign res[6] = 1'b0;
  assign res[7] = 1'b0;
  assign res[8] = 1'b0;
  assign res[9] = 1'b0;
  assign res[10] = 1'b0;
  assign res[11] = 1'b0;
  assign res[12] = 1'b0;
  assign res[13] = 1'b0;
  assign res[14] = 1'b0;
  assign res[15] = 1'b0;
  assign res[16] = 1'b0;
  assign res[17] = 1'b0;
  assign res[18] = 1'b0;
  assign res[19] = 1'b0;
  assign res[20] = 1'b0;
  assign res[21] = 1'b0;
  assign res[22] = 1'b0;
  assign res[23] = 1'b0;
  assign res[24] = 1'b0;
  assign res[25] = 1'b0;
  assign res[26] = 1'b0;
  assign res[27] = 1'b0;
  assign res[28] = 1'b0;
  assign res[29] = 1'b0;
  assign res[30] = 1'b0;
  assign res[31] = 1'b0;

  NORN_N32 compNORN ( .A(SUB), .Z(Z_s) );
  comparator compComparator ( .C(Cout), .Z(Z_s), .result(cmp_res_6bit) );
  MUX6_1 mpx ( .NEQ_LINE(cmp_res_6bit[0]), .EQ_LINE(cmp_res_6bit[1]), 
        .GEQ_LINE(cmp_res_6bit[2]), .G_LINE(cmp_res_6bit[3]), .L_LINE(
        cmp_res_6bit[4]), .LEQ_LINE(cmp_res_6bit[5]), .SEL(Sel), .RES_LINE(
        res[0]) );
endmodule


module MUX41_GENERIC_N32_1 ( SHIFTER_OUT, ADD_OUT, CMP_OUT, LOGICALS_OUT, SEL, 
        Y );
  input [31:0] SHIFTER_OUT;
  input [31:0] ADD_OUT;
  input [31:0] CMP_OUT;
  input [31:0] LOGICALS_OUT;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;

  AND2_X2 U1 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n4) );
  AND2_X2 U2 ( .A1(SEL[1]), .A2(n69), .ZN(n3) );
  NOR2_X4 U3 ( .A1(n69), .A2(SEL[1]), .ZN(n6) );
  NOR2_X4 U4 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n1), .A2(n2), .ZN(Y[9]) );
  AOI22_X1 U6 ( .A1(CMP_OUT[9]), .A2(n3), .B1(LOGICALS_OUT[9]), .B2(n4), .ZN(
        n2) );
  AOI22_X1 U7 ( .A1(SHIFTER_OUT[9]), .A2(n5), .B1(ADD_OUT[9]), .B2(n6), .ZN(n1) );
  NAND2_X1 U8 ( .A1(n7), .A2(n8), .ZN(Y[8]) );
  AOI22_X1 U9 ( .A1(CMP_OUT[8]), .A2(n3), .B1(LOGICALS_OUT[8]), .B2(n4), .ZN(
        n8) );
  AOI22_X1 U10 ( .A1(SHIFTER_OUT[8]), .A2(n5), .B1(ADD_OUT[8]), .B2(n6), .ZN(
        n7) );
  NAND2_X1 U11 ( .A1(n9), .A2(n10), .ZN(Y[7]) );
  AOI22_X1 U12 ( .A1(CMP_OUT[7]), .A2(n3), .B1(LOGICALS_OUT[7]), .B2(n4), .ZN(
        n10) );
  AOI22_X1 U13 ( .A1(SHIFTER_OUT[7]), .A2(n5), .B1(ADD_OUT[7]), .B2(n6), .ZN(
        n9) );
  NAND2_X1 U14 ( .A1(n11), .A2(n12), .ZN(Y[6]) );
  AOI22_X1 U15 ( .A1(CMP_OUT[6]), .A2(n3), .B1(LOGICALS_OUT[6]), .B2(n4), .ZN(
        n12) );
  AOI22_X1 U16 ( .A1(SHIFTER_OUT[6]), .A2(n5), .B1(ADD_OUT[6]), .B2(n6), .ZN(
        n11) );
  NAND2_X1 U17 ( .A1(n13), .A2(n14), .ZN(Y[5]) );
  AOI22_X1 U18 ( .A1(CMP_OUT[5]), .A2(n3), .B1(LOGICALS_OUT[5]), .B2(n4), .ZN(
        n14) );
  AOI22_X1 U19 ( .A1(SHIFTER_OUT[5]), .A2(n5), .B1(ADD_OUT[5]), .B2(n6), .ZN(
        n13) );
  NAND2_X1 U20 ( .A1(n15), .A2(n16), .ZN(Y[4]) );
  AOI22_X1 U21 ( .A1(CMP_OUT[4]), .A2(n3), .B1(LOGICALS_OUT[4]), .B2(n4), .ZN(
        n16) );
  AOI22_X1 U22 ( .A1(SHIFTER_OUT[4]), .A2(n5), .B1(ADD_OUT[4]), .B2(n6), .ZN(
        n15) );
  NAND2_X1 U23 ( .A1(n17), .A2(n18), .ZN(Y[3]) );
  AOI22_X1 U24 ( .A1(CMP_OUT[3]), .A2(n3), .B1(LOGICALS_OUT[3]), .B2(n4), .ZN(
        n18) );
  AOI22_X1 U25 ( .A1(SHIFTER_OUT[3]), .A2(n5), .B1(ADD_OUT[3]), .B2(n6), .ZN(
        n17) );
  NAND2_X1 U26 ( .A1(n19), .A2(n20), .ZN(Y[31]) );
  AOI22_X1 U27 ( .A1(CMP_OUT[31]), .A2(n3), .B1(LOGICALS_OUT[31]), .B2(n4), 
        .ZN(n20) );
  AOI22_X1 U28 ( .A1(SHIFTER_OUT[31]), .A2(n5), .B1(ADD_OUT[31]), .B2(n6), 
        .ZN(n19) );
  NAND2_X1 U29 ( .A1(n21), .A2(n22), .ZN(Y[30]) );
  AOI22_X1 U30 ( .A1(CMP_OUT[30]), .A2(n3), .B1(LOGICALS_OUT[30]), .B2(n4), 
        .ZN(n22) );
  AOI22_X1 U31 ( .A1(SHIFTER_OUT[30]), .A2(n5), .B1(ADD_OUT[30]), .B2(n6), 
        .ZN(n21) );
  NAND2_X1 U32 ( .A1(n23), .A2(n24), .ZN(Y[2]) );
  AOI22_X1 U33 ( .A1(CMP_OUT[2]), .A2(n3), .B1(LOGICALS_OUT[2]), .B2(n4), .ZN(
        n24) );
  AOI22_X1 U34 ( .A1(SHIFTER_OUT[2]), .A2(n5), .B1(ADD_OUT[2]), .B2(n6), .ZN(
        n23) );
  NAND2_X1 U35 ( .A1(n25), .A2(n26), .ZN(Y[29]) );
  AOI22_X1 U36 ( .A1(CMP_OUT[29]), .A2(n3), .B1(LOGICALS_OUT[29]), .B2(n4), 
        .ZN(n26) );
  AOI22_X1 U37 ( .A1(SHIFTER_OUT[29]), .A2(n5), .B1(ADD_OUT[29]), .B2(n6), 
        .ZN(n25) );
  NAND2_X1 U38 ( .A1(n27), .A2(n28), .ZN(Y[28]) );
  AOI22_X1 U39 ( .A1(CMP_OUT[28]), .A2(n3), .B1(LOGICALS_OUT[28]), .B2(n4), 
        .ZN(n28) );
  AOI22_X1 U40 ( .A1(SHIFTER_OUT[28]), .A2(n5), .B1(ADD_OUT[28]), .B2(n6), 
        .ZN(n27) );
  NAND2_X1 U41 ( .A1(n29), .A2(n30), .ZN(Y[27]) );
  AOI22_X1 U42 ( .A1(CMP_OUT[27]), .A2(n3), .B1(LOGICALS_OUT[27]), .B2(n4), 
        .ZN(n30) );
  AOI22_X1 U43 ( .A1(SHIFTER_OUT[27]), .A2(n5), .B1(ADD_OUT[27]), .B2(n6), 
        .ZN(n29) );
  NAND2_X1 U44 ( .A1(n31), .A2(n32), .ZN(Y[26]) );
  AOI22_X1 U45 ( .A1(CMP_OUT[26]), .A2(n3), .B1(LOGICALS_OUT[26]), .B2(n4), 
        .ZN(n32) );
  AOI22_X1 U46 ( .A1(SHIFTER_OUT[26]), .A2(n5), .B1(ADD_OUT[26]), .B2(n6), 
        .ZN(n31) );
  NAND2_X1 U47 ( .A1(n33), .A2(n34), .ZN(Y[25]) );
  AOI22_X1 U48 ( .A1(CMP_OUT[25]), .A2(n3), .B1(LOGICALS_OUT[25]), .B2(n4), 
        .ZN(n34) );
  AOI22_X1 U49 ( .A1(SHIFTER_OUT[25]), .A2(n5), .B1(ADD_OUT[25]), .B2(n6), 
        .ZN(n33) );
  NAND2_X1 U50 ( .A1(n35), .A2(n36), .ZN(Y[24]) );
  AOI22_X1 U51 ( .A1(CMP_OUT[24]), .A2(n3), .B1(LOGICALS_OUT[24]), .B2(n4), 
        .ZN(n36) );
  AOI22_X1 U52 ( .A1(SHIFTER_OUT[24]), .A2(n5), .B1(ADD_OUT[24]), .B2(n6), 
        .ZN(n35) );
  NAND2_X1 U53 ( .A1(n37), .A2(n38), .ZN(Y[23]) );
  AOI22_X1 U54 ( .A1(CMP_OUT[23]), .A2(n3), .B1(LOGICALS_OUT[23]), .B2(n4), 
        .ZN(n38) );
  AOI22_X1 U55 ( .A1(SHIFTER_OUT[23]), .A2(n5), .B1(ADD_OUT[23]), .B2(n6), 
        .ZN(n37) );
  NAND2_X1 U56 ( .A1(n39), .A2(n40), .ZN(Y[22]) );
  AOI22_X1 U57 ( .A1(CMP_OUT[22]), .A2(n3), .B1(LOGICALS_OUT[22]), .B2(n4), 
        .ZN(n40) );
  AOI22_X1 U58 ( .A1(SHIFTER_OUT[22]), .A2(n5), .B1(ADD_OUT[22]), .B2(n6), 
        .ZN(n39) );
  NAND2_X1 U59 ( .A1(n41), .A2(n42), .ZN(Y[21]) );
  AOI22_X1 U60 ( .A1(CMP_OUT[21]), .A2(n3), .B1(LOGICALS_OUT[21]), .B2(n4), 
        .ZN(n42) );
  AOI22_X1 U61 ( .A1(SHIFTER_OUT[21]), .A2(n5), .B1(ADD_OUT[21]), .B2(n6), 
        .ZN(n41) );
  NAND2_X1 U62 ( .A1(n43), .A2(n44), .ZN(Y[20]) );
  AOI22_X1 U63 ( .A1(CMP_OUT[20]), .A2(n3), .B1(LOGICALS_OUT[20]), .B2(n4), 
        .ZN(n44) );
  AOI22_X1 U64 ( .A1(SHIFTER_OUT[20]), .A2(n5), .B1(ADD_OUT[20]), .B2(n6), 
        .ZN(n43) );
  NAND2_X1 U65 ( .A1(n45), .A2(n46), .ZN(Y[1]) );
  AOI22_X1 U66 ( .A1(CMP_OUT[1]), .A2(n3), .B1(LOGICALS_OUT[1]), .B2(n4), .ZN(
        n46) );
  AOI22_X1 U67 ( .A1(SHIFTER_OUT[1]), .A2(n5), .B1(ADD_OUT[1]), .B2(n6), .ZN(
        n45) );
  NAND2_X1 U68 ( .A1(n47), .A2(n48), .ZN(Y[19]) );
  AOI22_X1 U69 ( .A1(CMP_OUT[19]), .A2(n3), .B1(LOGICALS_OUT[19]), .B2(n4), 
        .ZN(n48) );
  AOI22_X1 U70 ( .A1(SHIFTER_OUT[19]), .A2(n5), .B1(ADD_OUT[19]), .B2(n6), 
        .ZN(n47) );
  NAND2_X1 U71 ( .A1(n49), .A2(n50), .ZN(Y[18]) );
  AOI22_X1 U72 ( .A1(CMP_OUT[18]), .A2(n3), .B1(LOGICALS_OUT[18]), .B2(n4), 
        .ZN(n50) );
  AOI22_X1 U73 ( .A1(SHIFTER_OUT[18]), .A2(n5), .B1(ADD_OUT[18]), .B2(n6), 
        .ZN(n49) );
  NAND2_X1 U74 ( .A1(n51), .A2(n52), .ZN(Y[17]) );
  AOI22_X1 U75 ( .A1(CMP_OUT[17]), .A2(n3), .B1(LOGICALS_OUT[17]), .B2(n4), 
        .ZN(n52) );
  AOI22_X1 U76 ( .A1(SHIFTER_OUT[17]), .A2(n5), .B1(ADD_OUT[17]), .B2(n6), 
        .ZN(n51) );
  NAND2_X1 U77 ( .A1(n53), .A2(n54), .ZN(Y[16]) );
  AOI22_X1 U78 ( .A1(CMP_OUT[16]), .A2(n3), .B1(LOGICALS_OUT[16]), .B2(n4), 
        .ZN(n54) );
  AOI22_X1 U79 ( .A1(SHIFTER_OUT[16]), .A2(n5), .B1(ADD_OUT[16]), .B2(n6), 
        .ZN(n53) );
  NAND2_X1 U80 ( .A1(n55), .A2(n56), .ZN(Y[15]) );
  AOI22_X1 U81 ( .A1(CMP_OUT[15]), .A2(n3), .B1(LOGICALS_OUT[15]), .B2(n4), 
        .ZN(n56) );
  AOI22_X1 U82 ( .A1(SHIFTER_OUT[15]), .A2(n5), .B1(ADD_OUT[15]), .B2(n6), 
        .ZN(n55) );
  NAND2_X1 U83 ( .A1(n57), .A2(n58), .ZN(Y[14]) );
  AOI22_X1 U84 ( .A1(CMP_OUT[14]), .A2(n3), .B1(LOGICALS_OUT[14]), .B2(n4), 
        .ZN(n58) );
  AOI22_X1 U85 ( .A1(SHIFTER_OUT[14]), .A2(n5), .B1(ADD_OUT[14]), .B2(n6), 
        .ZN(n57) );
  NAND2_X1 U86 ( .A1(n59), .A2(n60), .ZN(Y[13]) );
  AOI22_X1 U87 ( .A1(CMP_OUT[13]), .A2(n3), .B1(LOGICALS_OUT[13]), .B2(n4), 
        .ZN(n60) );
  AOI22_X1 U88 ( .A1(SHIFTER_OUT[13]), .A2(n5), .B1(ADD_OUT[13]), .B2(n6), 
        .ZN(n59) );
  NAND2_X1 U89 ( .A1(n61), .A2(n62), .ZN(Y[12]) );
  AOI22_X1 U90 ( .A1(CMP_OUT[12]), .A2(n3), .B1(LOGICALS_OUT[12]), .B2(n4), 
        .ZN(n62) );
  AOI22_X1 U91 ( .A1(SHIFTER_OUT[12]), .A2(n5), .B1(ADD_OUT[12]), .B2(n6), 
        .ZN(n61) );
  NAND2_X1 U92 ( .A1(n63), .A2(n64), .ZN(Y[11]) );
  AOI22_X1 U93 ( .A1(CMP_OUT[11]), .A2(n3), .B1(LOGICALS_OUT[11]), .B2(n4), 
        .ZN(n64) );
  AOI22_X1 U94 ( .A1(SHIFTER_OUT[11]), .A2(n5), .B1(ADD_OUT[11]), .B2(n6), 
        .ZN(n63) );
  NAND2_X1 U95 ( .A1(n65), .A2(n66), .ZN(Y[10]) );
  AOI22_X1 U96 ( .A1(CMP_OUT[10]), .A2(n3), .B1(LOGICALS_OUT[10]), .B2(n4), 
        .ZN(n66) );
  AOI22_X1 U97 ( .A1(SHIFTER_OUT[10]), .A2(n5), .B1(ADD_OUT[10]), .B2(n6), 
        .ZN(n65) );
  NAND2_X1 U98 ( .A1(n67), .A2(n68), .ZN(Y[0]) );
  AOI22_X1 U99 ( .A1(CMP_OUT[0]), .A2(n3), .B1(LOGICALS_OUT[0]), .B2(n4), .ZN(
        n68) );
  AOI22_X1 U100 ( .A1(SHIFTER_OUT[0]), .A2(n5), .B1(ADD_OUT[0]), .B2(n6), .ZN(
        n67) );
  INV_X1 U101 ( .A(SEL[0]), .ZN(n69) );
endmodule


module ALU_N32_NBLOCK4 ( OPCODE, OPERANDA, OPERANDB, RESULT );
  input [5:0] OPCODE;
  input [31:0] OPERANDA;
  input [31:0] OPERANDB;
  output [31:0] RESULT;
  wire   cout, sign_delta, n1;
  wire   [31:0] add_result;
  wire   [31:0] shifter_result;
  wire   [31:0] logical_result;
  wire   [31:0] cmp_result;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  P4Adder_N32_K4 ADD_SUB ( .A(OPERANDA), .B(OPERANDB), .CIN(OPCODE[0]), .Cout(
        cout), .SUM(add_result) );
  ShifterT2_N32 SHIFTER ( .A(OPERANDA), .B(OPERANDB[4:0]), .sel(OPCODE[1:0]), 
        .\output (shifter_result) );
  LogicalT2_N32 LOGICAL_OP ( .A(OPERANDA), .B(OPERANDB), .S({OPCODE[0], 
        OPCODE[1], OPCODE[2], OPCODE[3]}), .Y(logical_result) );
  topLevelCMP_N32 COMPARATOR ( .SUB(add_result), .Cout(sign_delta), .Sel(
        OPCODE[3:1]), .res({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, cmp_result[0]}) );
  MUX41_GENERIC_N32_1 OUT_SELECT ( .SHIFTER_OUT(shifter_result), .ADD_OUT(
        add_result), .CMP_OUT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        cmp_result[0]}), .LOGICALS_OUT(logical_result), .SEL(OPCODE[5:4]), .Y(
        RESULT) );
  XOR2_X1 U1 ( .A(OPERANDA[31]), .B(n1), .Z(sign_delta) );
  XOR2_X1 U2 ( .A(cout), .B(OPERANDB[31]), .Z(n1) );
endmodule


module ffd_69 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_68 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_67 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_66 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_65 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_64 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_63 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_62 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_61 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_60 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_59 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_58 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_57 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_56 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_55 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_54 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_53 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_52 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_51 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_50 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_49 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_48 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_47 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_46 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_45 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_44 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_43 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_42 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_41 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_40 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_39 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X2 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_38 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n2, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n6), .CK(CK), .QN(n5) );
  INV_X4 U3 ( .A(n5), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n6) );
  MUX2_X1 U5 ( .A(n5), .B(n4), .S(En), .Z(n2) );
  INV_X1 U6 ( .A(D), .ZN(n4) );
endmodule


module regN_N32_2 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_69 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_68 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_67 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_66 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_65 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_64 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_63 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_62 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_61 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_60 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_59 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_58 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_57 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_56 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_55 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_54 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_53 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_52 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_51 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_50 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_49 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_48 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_47 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_46 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_45 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_44 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_43 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_42 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_41 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_40 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_39 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_38 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_37 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_36 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_35 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_34 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_33 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_32 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_31 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_30 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_29 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_28 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_27 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_26 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_25 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_24 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_23 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_22 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_21 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_20 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_19 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_18 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_17 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_16 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_15 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_14 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_13 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_12 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_11 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_10 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_9 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_8 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_7 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_6 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N32_1 ( regIn, Clk, Reset, Enable, regOut );
  input [31:0] regIn;
  output [31:0] regOut;
  input Clk, Reset, Enable;


  ffd_37 ffi_31 ( .D(regIn[31]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[31]) );
  ffd_36 ffi_30 ( .D(regIn[30]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[30]) );
  ffd_35 ffi_29 ( .D(regIn[29]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[29]) );
  ffd_34 ffi_28 ( .D(regIn[28]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[28]) );
  ffd_33 ffi_27 ( .D(regIn[27]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[27]) );
  ffd_32 ffi_26 ( .D(regIn[26]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[26]) );
  ffd_31 ffi_25 ( .D(regIn[25]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[25]) );
  ffd_30 ffi_24 ( .D(regIn[24]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[24]) );
  ffd_29 ffi_23 ( .D(regIn[23]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[23]) );
  ffd_28 ffi_22 ( .D(regIn[22]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[22]) );
  ffd_27 ffi_21 ( .D(regIn[21]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[21]) );
  ffd_26 ffi_20 ( .D(regIn[20]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[20]) );
  ffd_25 ffi_19 ( .D(regIn[19]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[19]) );
  ffd_24 ffi_18 ( .D(regIn[18]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[18]) );
  ffd_23 ffi_17 ( .D(regIn[17]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[17]) );
  ffd_22 ffi_16 ( .D(regIn[16]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[16]) );
  ffd_21 ffi_15 ( .D(regIn[15]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[15]) );
  ffd_20 ffi_14 ( .D(regIn[14]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[14]) );
  ffd_19 ffi_13 ( .D(regIn[13]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[13]) );
  ffd_18 ffi_12 ( .D(regIn[12]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[12]) );
  ffd_17 ffi_11 ( .D(regIn[11]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[11]) );
  ffd_16 ffi_10 ( .D(regIn[10]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[10]) );
  ffd_15 ffi_9 ( .D(regIn[9]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[9]) );
  ffd_14 ffi_8 ( .D(regIn[8]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[8]) );
  ffd_13 ffi_7 ( .D(regIn[7]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[7]) );
  ffd_12 ffi_6 ( .D(regIn[6]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[6]) );
  ffd_11 ffi_5 ( .D(regIn[5]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[5]) );
  ffd_10 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_9 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_8 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_7 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_6 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module ffd_5 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_4 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_3 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_2 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module ffd_1 ( D, CK, RESET, En, Q );
  input D, CK, RESET, En;
  output Q;
  wire   n1, n2, n4, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CK), .Q(Q), .QN(n4) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(n5) );
  MUX2_X1 U4 ( .A(n4), .B(n2), .S(En), .Z(n1) );
  INV_X1 U5 ( .A(D), .ZN(n2) );
endmodule


module regN_N5_1 ( regIn, Clk, Reset, Enable, regOut );
  input [4:0] regIn;
  output [4:0] regOut;
  input Clk, Reset, Enable;


  ffd_5 ffi_4 ( .D(regIn[4]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[4]) );
  ffd_4 ffi_3 ( .D(regIn[3]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[3]) );
  ffd_3 ffi_2 ( .D(regIn[2]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[2]) );
  ffd_2 ffi_1 ( .D(regIn[1]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[1]) );
  ffd_1 ffi_0 ( .D(regIn[0]), .CK(Clk), .RESET(Reset), .En(Enable), .Q(
        regOut[0]) );
endmodule


module EXUNIT_N32 ( NPC1, RD1, A, B, IMM, S1_A_NPC, S2_IMM_B, ALU_OPCODE, CLK, 
        RST, JUMP_EN, EN_REGN_ALU_OUT, JUMP, ALUOUT, ALU_OUT_REGN, B_OUT_REGN, 
        NPC2, RD2_OUT_REGN );
  input [31:0] NPC1;
  input [4:0] RD1;
  input [31:0] A;
  input [31:0] B;
  input [31:0] IMM;
  input [5:0] ALU_OPCODE;
  input [1:0] JUMP_EN;
  output [31:0] ALUOUT;
  output [31:0] ALU_OUT_REGN;
  output [31:0] B_OUT_REGN;
  output [31:0] NPC2;
  output [4:0] RD2_OUT_REGN;
  input S1_A_NPC, S2_IMM_B, CLK, RST, EN_REGN_ALU_OUT;
  output JUMP;
  wire   ZERO_CMP, n1;
  wire   [31:0] A_prime;
  wire   [31:0] B_prime;

  MUX21_GENERIC_NBIT32_4 COMP_MPX21_1 ( .A(NPC1), .B(A), .SEL(S1_A_NPC), .Y(
        A_prime) );
  MUX21_GENERIC_NBIT32_3 COMP_MPX21_2 ( .A(B), .B(IMM), .SEL(S2_IMM_B), .Y(
        B_prime) );
  ZERODET_N32 COMP_ZERO_CMP ( .A(A), .Y(ZERO_CMP) );
  MUX4_1 COMP_41_1MPX ( .ZERO(1'b0), .ONE(1'b1), .INV_CMP(n1), .CMP(ZERO_CMP), 
        .Sel(JUMP_EN), .Y(JUMP) );
  regN_N32_3 COMP_NPC2 ( .regIn(NPC1), .Clk(CLK), .Reset(RST), .Enable(
        EN_REGN_ALU_OUT), .regOut(NPC2) );
  ALU_N32_NBLOCK4 COMP_ALU ( .OPCODE(ALU_OPCODE), .OPERANDA(A_prime), 
        .OPERANDB(B_prime), .RESULT(ALUOUT) );
  regN_N32_2 COMP_REGN_ALUOUT ( .regIn(ALUOUT), .Clk(CLK), .Reset(RST), 
        .Enable(EN_REGN_ALU_OUT), .regOut(ALU_OUT_REGN) );
  regN_N32_1 COMP_REGN_BOUT ( .regIn(B), .Clk(CLK), .Reset(RST), .Enable(
        EN_REGN_ALU_OUT), .regOut(B_OUT_REGN) );
  regN_N5_1 COMP_REG5_RD2OUT ( .regIn(RD1), .Clk(CLK), .Reset(RST), .Enable(
        EN_REGN_ALU_OUT), .regOut(RD2_OUT_REGN) );
  INV_X1 U3 ( .A(ZERO_CMP), .ZN(n1) );
endmodule


module DataMemory_RAM_DEPTH32_WORD_SIZE32 ( Rst, Addr, Din, Dout, Sel, RM, WM, 
        EN, CLK );
  input [31:0] Addr;
  input [31:0] Din;
  output [31:0] Dout;
  input [2:0] Sel;
  input Rst, RM, WM, EN, CLK;
  wire   \DRAM_mem[0][31] , \DRAM_mem[0][30] , \DRAM_mem[0][29] ,
         \DRAM_mem[0][28] , \DRAM_mem[0][27] , \DRAM_mem[0][26] ,
         \DRAM_mem[0][25] , \DRAM_mem[0][24] , \DRAM_mem[0][23] ,
         \DRAM_mem[0][22] , \DRAM_mem[0][21] , \DRAM_mem[0][20] ,
         \DRAM_mem[0][19] , \DRAM_mem[0][18] , \DRAM_mem[0][17] ,
         \DRAM_mem[0][16] , \DRAM_mem[0][15] , \DRAM_mem[0][14] ,
         \DRAM_mem[0][13] , \DRAM_mem[0][12] , \DRAM_mem[0][11] ,
         \DRAM_mem[0][10] , \DRAM_mem[0][9] , \DRAM_mem[0][8] ,
         \DRAM_mem[0][7] , \DRAM_mem[0][6] , \DRAM_mem[0][5] ,
         \DRAM_mem[0][4] , \DRAM_mem[0][3] , \DRAM_mem[0][2] ,
         \DRAM_mem[0][1] , \DRAM_mem[0][0] , \DRAM_mem[1][31] ,
         \DRAM_mem[1][30] , \DRAM_mem[1][29] , \DRAM_mem[1][28] ,
         \DRAM_mem[1][27] , \DRAM_mem[1][26] , \DRAM_mem[1][25] ,
         \DRAM_mem[1][24] , \DRAM_mem[1][23] , \DRAM_mem[1][22] ,
         \DRAM_mem[1][21] , \DRAM_mem[1][20] , \DRAM_mem[1][19] ,
         \DRAM_mem[1][18] , \DRAM_mem[1][17] , \DRAM_mem[1][16] ,
         \DRAM_mem[1][15] , \DRAM_mem[1][14] , \DRAM_mem[1][13] ,
         \DRAM_mem[1][12] , \DRAM_mem[1][11] , \DRAM_mem[1][10] ,
         \DRAM_mem[1][9] , \DRAM_mem[1][8] , \DRAM_mem[1][7] ,
         \DRAM_mem[1][6] , \DRAM_mem[1][5] , \DRAM_mem[1][4] ,
         \DRAM_mem[1][3] , \DRAM_mem[1][2] , \DRAM_mem[1][1] ,
         \DRAM_mem[1][0] , \DRAM_mem[2][31] , \DRAM_mem[2][30] ,
         \DRAM_mem[2][29] , \DRAM_mem[2][28] , \DRAM_mem[2][27] ,
         \DRAM_mem[2][26] , \DRAM_mem[2][25] , \DRAM_mem[2][24] ,
         \DRAM_mem[2][23] , \DRAM_mem[2][22] , \DRAM_mem[2][21] ,
         \DRAM_mem[2][20] , \DRAM_mem[2][19] , \DRAM_mem[2][18] ,
         \DRAM_mem[2][17] , \DRAM_mem[2][16] , \DRAM_mem[2][15] ,
         \DRAM_mem[2][14] , \DRAM_mem[2][13] , \DRAM_mem[2][12] ,
         \DRAM_mem[2][11] , \DRAM_mem[2][10] , \DRAM_mem[2][9] ,
         \DRAM_mem[2][8] , \DRAM_mem[2][7] , \DRAM_mem[2][6] ,
         \DRAM_mem[2][5] , \DRAM_mem[2][4] , \DRAM_mem[2][3] ,
         \DRAM_mem[2][2] , \DRAM_mem[2][1] , \DRAM_mem[2][0] ,
         \DRAM_mem[3][31] , \DRAM_mem[3][30] , \DRAM_mem[3][29] ,
         \DRAM_mem[3][28] , \DRAM_mem[3][27] , \DRAM_mem[3][26] ,
         \DRAM_mem[3][25] , \DRAM_mem[3][24] , \DRAM_mem[3][23] ,
         \DRAM_mem[3][22] , \DRAM_mem[3][21] , \DRAM_mem[3][20] ,
         \DRAM_mem[3][19] , \DRAM_mem[3][18] , \DRAM_mem[3][17] ,
         \DRAM_mem[3][16] , \DRAM_mem[3][15] , \DRAM_mem[3][14] ,
         \DRAM_mem[3][13] , \DRAM_mem[3][12] , \DRAM_mem[3][11] ,
         \DRAM_mem[3][10] , \DRAM_mem[3][9] , \DRAM_mem[3][8] ,
         \DRAM_mem[3][7] , \DRAM_mem[3][6] , \DRAM_mem[3][5] ,
         \DRAM_mem[3][4] , \DRAM_mem[3][3] , \DRAM_mem[3][2] ,
         \DRAM_mem[3][1] , \DRAM_mem[3][0] , \DRAM_mem[4][31] ,
         \DRAM_mem[4][30] , \DRAM_mem[4][29] , \DRAM_mem[4][28] ,
         \DRAM_mem[4][27] , \DRAM_mem[4][26] , \DRAM_mem[4][25] ,
         \DRAM_mem[4][24] , \DRAM_mem[4][23] , \DRAM_mem[4][22] ,
         \DRAM_mem[4][21] , \DRAM_mem[4][20] , \DRAM_mem[4][19] ,
         \DRAM_mem[4][18] , \DRAM_mem[4][17] , \DRAM_mem[4][16] ,
         \DRAM_mem[4][15] , \DRAM_mem[4][14] , \DRAM_mem[4][13] ,
         \DRAM_mem[4][12] , \DRAM_mem[4][11] , \DRAM_mem[4][10] ,
         \DRAM_mem[4][9] , \DRAM_mem[4][8] , \DRAM_mem[4][7] ,
         \DRAM_mem[4][6] , \DRAM_mem[4][5] , \DRAM_mem[4][4] ,
         \DRAM_mem[4][3] , \DRAM_mem[4][2] , \DRAM_mem[4][1] ,
         \DRAM_mem[4][0] , \DRAM_mem[5][31] , \DRAM_mem[5][30] ,
         \DRAM_mem[5][29] , \DRAM_mem[5][28] , \DRAM_mem[5][27] ,
         \DRAM_mem[5][26] , \DRAM_mem[5][25] , \DRAM_mem[5][24] ,
         \DRAM_mem[5][23] , \DRAM_mem[5][22] , \DRAM_mem[5][21] ,
         \DRAM_mem[5][20] , \DRAM_mem[5][19] , \DRAM_mem[5][18] ,
         \DRAM_mem[5][17] , \DRAM_mem[5][16] , \DRAM_mem[5][15] ,
         \DRAM_mem[5][14] , \DRAM_mem[5][13] , \DRAM_mem[5][12] ,
         \DRAM_mem[5][11] , \DRAM_mem[5][10] , \DRAM_mem[5][9] ,
         \DRAM_mem[5][8] , \DRAM_mem[5][7] , \DRAM_mem[5][6] ,
         \DRAM_mem[5][5] , \DRAM_mem[5][4] , \DRAM_mem[5][3] ,
         \DRAM_mem[5][2] , \DRAM_mem[5][1] , \DRAM_mem[5][0] ,
         \DRAM_mem[6][31] , \DRAM_mem[6][30] , \DRAM_mem[6][29] ,
         \DRAM_mem[6][28] , \DRAM_mem[6][27] , \DRAM_mem[6][26] ,
         \DRAM_mem[6][25] , \DRAM_mem[6][24] , \DRAM_mem[6][23] ,
         \DRAM_mem[6][22] , \DRAM_mem[6][21] , \DRAM_mem[6][20] ,
         \DRAM_mem[6][19] , \DRAM_mem[6][18] , \DRAM_mem[6][17] ,
         \DRAM_mem[6][16] , \DRAM_mem[6][15] , \DRAM_mem[6][14] ,
         \DRAM_mem[6][13] , \DRAM_mem[6][12] , \DRAM_mem[6][11] ,
         \DRAM_mem[6][10] , \DRAM_mem[6][9] , \DRAM_mem[6][8] ,
         \DRAM_mem[6][7] , \DRAM_mem[6][6] , \DRAM_mem[6][5] ,
         \DRAM_mem[6][4] , \DRAM_mem[6][3] , \DRAM_mem[6][2] ,
         \DRAM_mem[6][1] , \DRAM_mem[6][0] , \DRAM_mem[7][31] ,
         \DRAM_mem[7][30] , \DRAM_mem[7][29] , \DRAM_mem[7][28] ,
         \DRAM_mem[7][27] , \DRAM_mem[7][26] , \DRAM_mem[7][25] ,
         \DRAM_mem[7][24] , \DRAM_mem[7][23] , \DRAM_mem[7][22] ,
         \DRAM_mem[7][21] , \DRAM_mem[7][20] , \DRAM_mem[7][19] ,
         \DRAM_mem[7][18] , \DRAM_mem[7][17] , \DRAM_mem[7][16] ,
         \DRAM_mem[7][15] , \DRAM_mem[7][14] , \DRAM_mem[7][13] ,
         \DRAM_mem[7][12] , \DRAM_mem[7][11] , \DRAM_mem[7][10] ,
         \DRAM_mem[7][9] , \DRAM_mem[7][8] , \DRAM_mem[7][7] ,
         \DRAM_mem[7][6] , \DRAM_mem[7][5] , \DRAM_mem[7][4] ,
         \DRAM_mem[7][3] , \DRAM_mem[7][2] , \DRAM_mem[7][1] ,
         \DRAM_mem[7][0] , \DRAM_mem[8][31] , \DRAM_mem[8][30] ,
         \DRAM_mem[8][29] , \DRAM_mem[8][28] , \DRAM_mem[8][27] ,
         \DRAM_mem[8][26] , \DRAM_mem[8][25] , \DRAM_mem[8][24] ,
         \DRAM_mem[8][23] , \DRAM_mem[8][22] , \DRAM_mem[8][21] ,
         \DRAM_mem[8][20] , \DRAM_mem[8][19] , \DRAM_mem[8][18] ,
         \DRAM_mem[8][17] , \DRAM_mem[8][16] , \DRAM_mem[8][15] ,
         \DRAM_mem[8][14] , \DRAM_mem[8][13] , \DRAM_mem[8][12] ,
         \DRAM_mem[8][11] , \DRAM_mem[8][10] , \DRAM_mem[8][9] ,
         \DRAM_mem[8][8] , \DRAM_mem[8][7] , \DRAM_mem[8][6] ,
         \DRAM_mem[8][5] , \DRAM_mem[8][4] , \DRAM_mem[8][3] ,
         \DRAM_mem[8][2] , \DRAM_mem[8][1] , \DRAM_mem[8][0] ,
         \DRAM_mem[9][31] , \DRAM_mem[9][30] , \DRAM_mem[9][29] ,
         \DRAM_mem[9][28] , \DRAM_mem[9][27] , \DRAM_mem[9][26] ,
         \DRAM_mem[9][25] , \DRAM_mem[9][24] , \DRAM_mem[9][23] ,
         \DRAM_mem[9][22] , \DRAM_mem[9][21] , \DRAM_mem[9][20] ,
         \DRAM_mem[9][19] , \DRAM_mem[9][18] , \DRAM_mem[9][17] ,
         \DRAM_mem[9][16] , \DRAM_mem[9][15] , \DRAM_mem[9][14] ,
         \DRAM_mem[9][13] , \DRAM_mem[9][12] , \DRAM_mem[9][11] ,
         \DRAM_mem[9][10] , \DRAM_mem[9][9] , \DRAM_mem[9][8] ,
         \DRAM_mem[9][7] , \DRAM_mem[9][6] , \DRAM_mem[9][5] ,
         \DRAM_mem[9][4] , \DRAM_mem[9][3] , \DRAM_mem[9][2] ,
         \DRAM_mem[9][1] , \DRAM_mem[9][0] , \DRAM_mem[10][31] ,
         \DRAM_mem[10][30] , \DRAM_mem[10][29] , \DRAM_mem[10][28] ,
         \DRAM_mem[10][27] , \DRAM_mem[10][26] , \DRAM_mem[10][25] ,
         \DRAM_mem[10][24] , \DRAM_mem[10][23] , \DRAM_mem[10][22] ,
         \DRAM_mem[10][21] , \DRAM_mem[10][20] , \DRAM_mem[10][19] ,
         \DRAM_mem[10][18] , \DRAM_mem[10][17] , \DRAM_mem[10][16] ,
         \DRAM_mem[10][15] , \DRAM_mem[10][14] , \DRAM_mem[10][13] ,
         \DRAM_mem[10][12] , \DRAM_mem[10][11] , \DRAM_mem[10][10] ,
         \DRAM_mem[10][9] , \DRAM_mem[10][8] , \DRAM_mem[10][7] ,
         \DRAM_mem[10][6] , \DRAM_mem[10][5] , \DRAM_mem[10][4] ,
         \DRAM_mem[10][3] , \DRAM_mem[10][2] , \DRAM_mem[10][1] ,
         \DRAM_mem[10][0] , \DRAM_mem[11][31] , \DRAM_mem[11][30] ,
         \DRAM_mem[11][29] , \DRAM_mem[11][28] , \DRAM_mem[11][27] ,
         \DRAM_mem[11][26] , \DRAM_mem[11][25] , \DRAM_mem[11][24] ,
         \DRAM_mem[11][23] , \DRAM_mem[11][22] , \DRAM_mem[11][21] ,
         \DRAM_mem[11][20] , \DRAM_mem[11][19] , \DRAM_mem[11][18] ,
         \DRAM_mem[11][17] , \DRAM_mem[11][16] , \DRAM_mem[11][15] ,
         \DRAM_mem[11][14] , \DRAM_mem[11][13] , \DRAM_mem[11][12] ,
         \DRAM_mem[11][11] , \DRAM_mem[11][10] , \DRAM_mem[11][9] ,
         \DRAM_mem[11][8] , \DRAM_mem[11][7] , \DRAM_mem[11][6] ,
         \DRAM_mem[11][5] , \DRAM_mem[11][4] , \DRAM_mem[11][3] ,
         \DRAM_mem[11][2] , \DRAM_mem[11][1] , \DRAM_mem[11][0] ,
         \DRAM_mem[12][31] , \DRAM_mem[12][30] , \DRAM_mem[12][29] ,
         \DRAM_mem[12][28] , \DRAM_mem[12][27] , \DRAM_mem[12][26] ,
         \DRAM_mem[12][25] , \DRAM_mem[12][24] , \DRAM_mem[12][23] ,
         \DRAM_mem[12][22] , \DRAM_mem[12][21] , \DRAM_mem[12][20] ,
         \DRAM_mem[12][19] , \DRAM_mem[12][18] , \DRAM_mem[12][17] ,
         \DRAM_mem[12][16] , \DRAM_mem[12][15] , \DRAM_mem[12][14] ,
         \DRAM_mem[12][13] , \DRAM_mem[12][12] , \DRAM_mem[12][11] ,
         \DRAM_mem[12][10] , \DRAM_mem[12][9] , \DRAM_mem[12][8] ,
         \DRAM_mem[12][7] , \DRAM_mem[12][6] , \DRAM_mem[12][5] ,
         \DRAM_mem[12][4] , \DRAM_mem[12][3] , \DRAM_mem[12][2] ,
         \DRAM_mem[12][1] , \DRAM_mem[12][0] , \DRAM_mem[13][31] ,
         \DRAM_mem[13][30] , \DRAM_mem[13][29] , \DRAM_mem[13][28] ,
         \DRAM_mem[13][27] , \DRAM_mem[13][26] , \DRAM_mem[13][25] ,
         \DRAM_mem[13][24] , \DRAM_mem[13][23] , \DRAM_mem[13][22] ,
         \DRAM_mem[13][21] , \DRAM_mem[13][20] , \DRAM_mem[13][19] ,
         \DRAM_mem[13][18] , \DRAM_mem[13][17] , \DRAM_mem[13][16] ,
         \DRAM_mem[13][15] , \DRAM_mem[13][14] , \DRAM_mem[13][13] ,
         \DRAM_mem[13][12] , \DRAM_mem[13][11] , \DRAM_mem[13][10] ,
         \DRAM_mem[13][9] , \DRAM_mem[13][8] , \DRAM_mem[13][7] ,
         \DRAM_mem[13][6] , \DRAM_mem[13][5] , \DRAM_mem[13][4] ,
         \DRAM_mem[13][3] , \DRAM_mem[13][2] , \DRAM_mem[13][1] ,
         \DRAM_mem[13][0] , \DRAM_mem[14][31] , \DRAM_mem[14][30] ,
         \DRAM_mem[14][29] , \DRAM_mem[14][28] , \DRAM_mem[14][27] ,
         \DRAM_mem[14][26] , \DRAM_mem[14][25] , \DRAM_mem[14][24] ,
         \DRAM_mem[14][23] , \DRAM_mem[14][22] , \DRAM_mem[14][21] ,
         \DRAM_mem[14][20] , \DRAM_mem[14][19] , \DRAM_mem[14][18] ,
         \DRAM_mem[14][17] , \DRAM_mem[14][16] , \DRAM_mem[14][15] ,
         \DRAM_mem[14][14] , \DRAM_mem[14][13] , \DRAM_mem[14][12] ,
         \DRAM_mem[14][11] , \DRAM_mem[14][10] , \DRAM_mem[14][9] ,
         \DRAM_mem[14][8] , \DRAM_mem[14][7] , \DRAM_mem[14][6] ,
         \DRAM_mem[14][5] , \DRAM_mem[14][4] , \DRAM_mem[14][3] ,
         \DRAM_mem[14][2] , \DRAM_mem[14][1] , \DRAM_mem[14][0] ,
         \DRAM_mem[15][31] , \DRAM_mem[15][30] , \DRAM_mem[15][29] ,
         \DRAM_mem[15][28] , \DRAM_mem[15][27] , \DRAM_mem[15][26] ,
         \DRAM_mem[15][25] , \DRAM_mem[15][24] , \DRAM_mem[15][23] ,
         \DRAM_mem[15][22] , \DRAM_mem[15][21] , \DRAM_mem[15][20] ,
         \DRAM_mem[15][19] , \DRAM_mem[15][18] , \DRAM_mem[15][17] ,
         \DRAM_mem[15][16] , \DRAM_mem[15][15] , \DRAM_mem[15][14] ,
         \DRAM_mem[15][13] , \DRAM_mem[15][12] , \DRAM_mem[15][11] ,
         \DRAM_mem[15][10] , \DRAM_mem[15][9] , \DRAM_mem[15][8] ,
         \DRAM_mem[15][7] , \DRAM_mem[15][6] , \DRAM_mem[15][5] ,
         \DRAM_mem[15][4] , \DRAM_mem[15][3] , \DRAM_mem[15][2] ,
         \DRAM_mem[15][1] , \DRAM_mem[15][0] , \DRAM_mem[16][31] ,
         \DRAM_mem[16][30] , \DRAM_mem[16][29] , \DRAM_mem[16][28] ,
         \DRAM_mem[16][27] , \DRAM_mem[16][26] , \DRAM_mem[16][25] ,
         \DRAM_mem[16][24] , \DRAM_mem[16][23] , \DRAM_mem[16][22] ,
         \DRAM_mem[16][21] , \DRAM_mem[16][20] , \DRAM_mem[16][19] ,
         \DRAM_mem[16][18] , \DRAM_mem[16][17] , \DRAM_mem[16][16] ,
         \DRAM_mem[16][15] , \DRAM_mem[16][14] , \DRAM_mem[16][13] ,
         \DRAM_mem[16][12] , \DRAM_mem[16][11] , \DRAM_mem[16][10] ,
         \DRAM_mem[16][9] , \DRAM_mem[16][8] , \DRAM_mem[16][7] ,
         \DRAM_mem[16][6] , \DRAM_mem[16][5] , \DRAM_mem[16][4] ,
         \DRAM_mem[16][3] , \DRAM_mem[16][2] , \DRAM_mem[16][1] ,
         \DRAM_mem[16][0] , \DRAM_mem[17][31] , \DRAM_mem[17][30] ,
         \DRAM_mem[17][29] , \DRAM_mem[17][28] , \DRAM_mem[17][27] ,
         \DRAM_mem[17][26] , \DRAM_mem[17][25] , \DRAM_mem[17][24] ,
         \DRAM_mem[17][23] , \DRAM_mem[17][22] , \DRAM_mem[17][21] ,
         \DRAM_mem[17][20] , \DRAM_mem[17][19] , \DRAM_mem[17][18] ,
         \DRAM_mem[17][17] , \DRAM_mem[17][16] , \DRAM_mem[17][15] ,
         \DRAM_mem[17][14] , \DRAM_mem[17][13] , \DRAM_mem[17][12] ,
         \DRAM_mem[17][11] , \DRAM_mem[17][10] , \DRAM_mem[17][9] ,
         \DRAM_mem[17][8] , \DRAM_mem[17][7] , \DRAM_mem[17][6] ,
         \DRAM_mem[17][5] , \DRAM_mem[17][4] , \DRAM_mem[17][3] ,
         \DRAM_mem[17][2] , \DRAM_mem[17][1] , \DRAM_mem[17][0] ,
         \DRAM_mem[18][31] , \DRAM_mem[18][30] , \DRAM_mem[18][29] ,
         \DRAM_mem[18][28] , \DRAM_mem[18][27] , \DRAM_mem[18][26] ,
         \DRAM_mem[18][25] , \DRAM_mem[18][24] , \DRAM_mem[18][23] ,
         \DRAM_mem[18][22] , \DRAM_mem[18][21] , \DRAM_mem[18][20] ,
         \DRAM_mem[18][19] , \DRAM_mem[18][18] , \DRAM_mem[18][17] ,
         \DRAM_mem[18][16] , \DRAM_mem[18][15] , \DRAM_mem[18][14] ,
         \DRAM_mem[18][13] , \DRAM_mem[18][12] , \DRAM_mem[18][11] ,
         \DRAM_mem[18][10] , \DRAM_mem[18][9] , \DRAM_mem[18][8] ,
         \DRAM_mem[18][7] , \DRAM_mem[18][6] , \DRAM_mem[18][5] ,
         \DRAM_mem[18][4] , \DRAM_mem[18][3] , \DRAM_mem[18][2] ,
         \DRAM_mem[18][1] , \DRAM_mem[18][0] , \DRAM_mem[19][31] ,
         \DRAM_mem[19][30] , \DRAM_mem[19][29] , \DRAM_mem[19][28] ,
         \DRAM_mem[19][27] , \DRAM_mem[19][26] , \DRAM_mem[19][25] ,
         \DRAM_mem[19][24] , \DRAM_mem[19][23] , \DRAM_mem[19][22] ,
         \DRAM_mem[19][21] , \DRAM_mem[19][20] , \DRAM_mem[19][19] ,
         \DRAM_mem[19][18] , \DRAM_mem[19][17] , \DRAM_mem[19][16] ,
         \DRAM_mem[19][15] , \DRAM_mem[19][14] , \DRAM_mem[19][13] ,
         \DRAM_mem[19][12] , \DRAM_mem[19][11] , \DRAM_mem[19][10] ,
         \DRAM_mem[19][9] , \DRAM_mem[19][8] , \DRAM_mem[19][7] ,
         \DRAM_mem[19][6] , \DRAM_mem[19][5] , \DRAM_mem[19][4] ,
         \DRAM_mem[19][3] , \DRAM_mem[19][2] , \DRAM_mem[19][1] ,
         \DRAM_mem[19][0] , \DRAM_mem[20][31] , \DRAM_mem[20][30] ,
         \DRAM_mem[20][29] , \DRAM_mem[20][28] , \DRAM_mem[20][27] ,
         \DRAM_mem[20][26] , \DRAM_mem[20][25] , \DRAM_mem[20][24] ,
         \DRAM_mem[20][23] , \DRAM_mem[20][22] , \DRAM_mem[20][21] ,
         \DRAM_mem[20][20] , \DRAM_mem[20][19] , \DRAM_mem[20][18] ,
         \DRAM_mem[20][17] , \DRAM_mem[20][16] , \DRAM_mem[20][15] ,
         \DRAM_mem[20][14] , \DRAM_mem[20][13] , \DRAM_mem[20][12] ,
         \DRAM_mem[20][11] , \DRAM_mem[20][10] , \DRAM_mem[20][9] ,
         \DRAM_mem[20][8] , \DRAM_mem[20][7] , \DRAM_mem[20][6] ,
         \DRAM_mem[20][5] , \DRAM_mem[20][4] , \DRAM_mem[20][3] ,
         \DRAM_mem[20][2] , \DRAM_mem[20][1] , \DRAM_mem[20][0] ,
         \DRAM_mem[21][31] , \DRAM_mem[21][30] , \DRAM_mem[21][29] ,
         \DRAM_mem[21][28] , \DRAM_mem[21][27] , \DRAM_mem[21][26] ,
         \DRAM_mem[21][25] , \DRAM_mem[21][24] , \DRAM_mem[21][23] ,
         \DRAM_mem[21][22] , \DRAM_mem[21][21] , \DRAM_mem[21][20] ,
         \DRAM_mem[21][19] , \DRAM_mem[21][18] , \DRAM_mem[21][17] ,
         \DRAM_mem[21][16] , \DRAM_mem[21][15] , \DRAM_mem[21][14] ,
         \DRAM_mem[21][13] , \DRAM_mem[21][12] , \DRAM_mem[21][11] ,
         \DRAM_mem[21][10] , \DRAM_mem[21][9] , \DRAM_mem[21][8] ,
         \DRAM_mem[21][7] , \DRAM_mem[21][6] , \DRAM_mem[21][5] ,
         \DRAM_mem[21][4] , \DRAM_mem[21][3] , \DRAM_mem[21][2] ,
         \DRAM_mem[21][1] , \DRAM_mem[21][0] , \DRAM_mem[22][31] ,
         \DRAM_mem[22][30] , \DRAM_mem[22][29] , \DRAM_mem[22][28] ,
         \DRAM_mem[22][27] , \DRAM_mem[22][26] , \DRAM_mem[22][25] ,
         \DRAM_mem[22][24] , \DRAM_mem[22][23] , \DRAM_mem[22][22] ,
         \DRAM_mem[22][21] , \DRAM_mem[22][20] , \DRAM_mem[22][19] ,
         \DRAM_mem[22][18] , \DRAM_mem[22][17] , \DRAM_mem[22][16] ,
         \DRAM_mem[22][15] , \DRAM_mem[22][14] , \DRAM_mem[22][13] ,
         \DRAM_mem[22][12] , \DRAM_mem[22][11] , \DRAM_mem[22][10] ,
         \DRAM_mem[22][9] , \DRAM_mem[22][8] , \DRAM_mem[22][7] ,
         \DRAM_mem[22][6] , \DRAM_mem[22][5] , \DRAM_mem[22][4] ,
         \DRAM_mem[22][3] , \DRAM_mem[22][2] , \DRAM_mem[22][1] ,
         \DRAM_mem[22][0] , \DRAM_mem[23][31] , \DRAM_mem[23][30] ,
         \DRAM_mem[23][29] , \DRAM_mem[23][28] , \DRAM_mem[23][27] ,
         \DRAM_mem[23][26] , \DRAM_mem[23][25] , \DRAM_mem[23][24] ,
         \DRAM_mem[23][23] , \DRAM_mem[23][22] , \DRAM_mem[23][21] ,
         \DRAM_mem[23][20] , \DRAM_mem[23][19] , \DRAM_mem[23][18] ,
         \DRAM_mem[23][17] , \DRAM_mem[23][16] , \DRAM_mem[23][15] ,
         \DRAM_mem[23][14] , \DRAM_mem[23][13] , \DRAM_mem[23][12] ,
         \DRAM_mem[23][11] , \DRAM_mem[23][10] , \DRAM_mem[23][9] ,
         \DRAM_mem[23][8] , \DRAM_mem[23][7] , \DRAM_mem[23][6] ,
         \DRAM_mem[23][5] , \DRAM_mem[23][4] , \DRAM_mem[23][3] ,
         \DRAM_mem[23][2] , \DRAM_mem[23][1] , \DRAM_mem[23][0] ,
         \DRAM_mem[24][31] , \DRAM_mem[24][30] , \DRAM_mem[24][29] ,
         \DRAM_mem[24][28] , \DRAM_mem[24][27] , \DRAM_mem[24][26] ,
         \DRAM_mem[24][25] , \DRAM_mem[24][24] , \DRAM_mem[24][23] ,
         \DRAM_mem[24][22] , \DRAM_mem[24][21] , \DRAM_mem[24][20] ,
         \DRAM_mem[24][19] , \DRAM_mem[24][18] , \DRAM_mem[24][17] ,
         \DRAM_mem[24][16] , \DRAM_mem[24][15] , \DRAM_mem[24][14] ,
         \DRAM_mem[24][13] , \DRAM_mem[24][12] , \DRAM_mem[24][11] ,
         \DRAM_mem[24][10] , \DRAM_mem[24][9] , \DRAM_mem[24][8] ,
         \DRAM_mem[24][7] , \DRAM_mem[24][6] , \DRAM_mem[24][5] ,
         \DRAM_mem[24][4] , \DRAM_mem[24][3] , \DRAM_mem[24][2] ,
         \DRAM_mem[24][1] , \DRAM_mem[24][0] , \DRAM_mem[25][31] ,
         \DRAM_mem[25][30] , \DRAM_mem[25][29] , \DRAM_mem[25][28] ,
         \DRAM_mem[25][27] , \DRAM_mem[25][26] , \DRAM_mem[25][25] ,
         \DRAM_mem[25][24] , \DRAM_mem[25][23] , \DRAM_mem[25][22] ,
         \DRAM_mem[25][21] , \DRAM_mem[25][20] , \DRAM_mem[25][19] ,
         \DRAM_mem[25][18] , \DRAM_mem[25][17] , \DRAM_mem[25][16] ,
         \DRAM_mem[25][15] , \DRAM_mem[25][14] , \DRAM_mem[25][13] ,
         \DRAM_mem[25][12] , \DRAM_mem[25][11] , \DRAM_mem[25][10] ,
         \DRAM_mem[25][9] , \DRAM_mem[25][8] , \DRAM_mem[25][7] ,
         \DRAM_mem[25][6] , \DRAM_mem[25][5] , \DRAM_mem[25][4] ,
         \DRAM_mem[25][3] , \DRAM_mem[25][2] , \DRAM_mem[25][1] ,
         \DRAM_mem[25][0] , \DRAM_mem[26][31] , \DRAM_mem[26][30] ,
         \DRAM_mem[26][29] , \DRAM_mem[26][28] , \DRAM_mem[26][27] ,
         \DRAM_mem[26][26] , \DRAM_mem[26][25] , \DRAM_mem[26][24] ,
         \DRAM_mem[26][23] , \DRAM_mem[26][22] , \DRAM_mem[26][21] ,
         \DRAM_mem[26][20] , \DRAM_mem[26][19] , \DRAM_mem[26][18] ,
         \DRAM_mem[26][17] , \DRAM_mem[26][16] , \DRAM_mem[26][15] ,
         \DRAM_mem[26][14] , \DRAM_mem[26][13] , \DRAM_mem[26][12] ,
         \DRAM_mem[26][11] , \DRAM_mem[26][10] , \DRAM_mem[26][9] ,
         \DRAM_mem[26][8] , \DRAM_mem[26][7] , \DRAM_mem[26][6] ,
         \DRAM_mem[26][5] , \DRAM_mem[26][4] , \DRAM_mem[26][3] ,
         \DRAM_mem[26][2] , \DRAM_mem[26][1] , \DRAM_mem[26][0] ,
         \DRAM_mem[27][31] , \DRAM_mem[27][30] , \DRAM_mem[27][29] ,
         \DRAM_mem[27][28] , \DRAM_mem[27][27] , \DRAM_mem[27][26] ,
         \DRAM_mem[27][25] , \DRAM_mem[27][24] , \DRAM_mem[27][23] ,
         \DRAM_mem[27][22] , \DRAM_mem[27][21] , \DRAM_mem[27][20] ,
         \DRAM_mem[27][19] , \DRAM_mem[27][18] , \DRAM_mem[27][17] ,
         \DRAM_mem[27][16] , \DRAM_mem[27][15] , \DRAM_mem[27][14] ,
         \DRAM_mem[27][13] , \DRAM_mem[27][12] , \DRAM_mem[27][11] ,
         \DRAM_mem[27][10] , \DRAM_mem[27][9] , \DRAM_mem[27][8] ,
         \DRAM_mem[27][7] , \DRAM_mem[27][6] , \DRAM_mem[27][5] ,
         \DRAM_mem[27][4] , \DRAM_mem[27][3] , \DRAM_mem[27][2] ,
         \DRAM_mem[27][1] , \DRAM_mem[27][0] , \DRAM_mem[28][31] ,
         \DRAM_mem[28][30] , \DRAM_mem[28][29] , \DRAM_mem[28][28] ,
         \DRAM_mem[28][27] , \DRAM_mem[28][26] , \DRAM_mem[28][25] ,
         \DRAM_mem[28][24] , \DRAM_mem[28][23] , \DRAM_mem[28][22] ,
         \DRAM_mem[28][21] , \DRAM_mem[28][20] , \DRAM_mem[28][19] ,
         \DRAM_mem[28][18] , \DRAM_mem[28][17] , \DRAM_mem[28][16] ,
         \DRAM_mem[28][15] , \DRAM_mem[28][14] , \DRAM_mem[28][13] ,
         \DRAM_mem[28][12] , \DRAM_mem[28][11] , \DRAM_mem[28][10] ,
         \DRAM_mem[28][9] , \DRAM_mem[28][8] , \DRAM_mem[28][7] ,
         \DRAM_mem[28][6] , \DRAM_mem[28][5] , \DRAM_mem[28][4] ,
         \DRAM_mem[28][3] , \DRAM_mem[28][2] , \DRAM_mem[28][1] ,
         \DRAM_mem[28][0] , \DRAM_mem[29][31] , \DRAM_mem[29][30] ,
         \DRAM_mem[29][29] , \DRAM_mem[29][28] , \DRAM_mem[29][27] ,
         \DRAM_mem[29][26] , \DRAM_mem[29][25] , \DRAM_mem[29][24] ,
         \DRAM_mem[29][23] , \DRAM_mem[29][22] , \DRAM_mem[29][21] ,
         \DRAM_mem[29][20] , \DRAM_mem[29][19] , \DRAM_mem[29][18] ,
         \DRAM_mem[29][17] , \DRAM_mem[29][16] , \DRAM_mem[29][15] ,
         \DRAM_mem[29][14] , \DRAM_mem[29][13] , \DRAM_mem[29][12] ,
         \DRAM_mem[29][11] , \DRAM_mem[29][10] , \DRAM_mem[29][9] ,
         \DRAM_mem[29][8] , \DRAM_mem[29][7] , \DRAM_mem[29][6] ,
         \DRAM_mem[29][5] , \DRAM_mem[29][4] , \DRAM_mem[29][3] ,
         \DRAM_mem[29][2] , \DRAM_mem[29][1] , \DRAM_mem[29][0] ,
         \DRAM_mem[30][31] , \DRAM_mem[30][30] , \DRAM_mem[30][29] ,
         \DRAM_mem[30][28] , \DRAM_mem[30][27] , \DRAM_mem[30][26] ,
         \DRAM_mem[30][25] , \DRAM_mem[30][24] , \DRAM_mem[30][23] ,
         \DRAM_mem[30][22] , \DRAM_mem[30][21] , \DRAM_mem[30][20] ,
         \DRAM_mem[30][19] , \DRAM_mem[30][18] , \DRAM_mem[30][17] ,
         \DRAM_mem[30][16] , \DRAM_mem[30][15] , \DRAM_mem[30][14] ,
         \DRAM_mem[30][13] , \DRAM_mem[30][12] , \DRAM_mem[30][11] ,
         \DRAM_mem[30][10] , \DRAM_mem[30][9] , \DRAM_mem[30][8] ,
         \DRAM_mem[30][7] , \DRAM_mem[30][6] , \DRAM_mem[30][5] ,
         \DRAM_mem[30][4] , \DRAM_mem[30][3] , \DRAM_mem[30][2] ,
         \DRAM_mem[30][1] , \DRAM_mem[30][0] , \DRAM_mem[31][31] ,
         \DRAM_mem[31][30] , \DRAM_mem[31][29] , \DRAM_mem[31][28] ,
         \DRAM_mem[31][27] , \DRAM_mem[31][26] , \DRAM_mem[31][25] ,
         \DRAM_mem[31][24] , \DRAM_mem[31][23] , \DRAM_mem[31][22] ,
         \DRAM_mem[31][21] , \DRAM_mem[31][20] , \DRAM_mem[31][19] ,
         \DRAM_mem[31][18] , \DRAM_mem[31][17] , \DRAM_mem[31][16] ,
         \DRAM_mem[31][15] , \DRAM_mem[31][14] , \DRAM_mem[31][13] ,
         \DRAM_mem[31][12] , \DRAM_mem[31][11] , \DRAM_mem[31][10] ,
         \DRAM_mem[31][9] , \DRAM_mem[31][8] , \DRAM_mem[31][7] ,
         \DRAM_mem[31][6] , \DRAM_mem[31][5] , \DRAM_mem[31][4] ,
         \DRAM_mem[31][3] , \DRAM_mem[31][2] , \DRAM_mem[31][1] ,
         \DRAM_mem[31][0] , N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;

  DFFR_X1 \DRAM_mem_reg[0][31]  ( .D(n2180), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[0][31] ) );
  DFFR_X1 \DRAM_mem_reg[0][30]  ( .D(n2179), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[0][30] ) );
  DFFR_X1 \DRAM_mem_reg[0][29]  ( .D(n2178), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[0][29] ) );
  DFFR_X1 \DRAM_mem_reg[0][28]  ( .D(n2177), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[0][28] ) );
  DFFR_X1 \DRAM_mem_reg[0][27]  ( .D(n2176), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[0][27] ) );
  DFFR_X1 \DRAM_mem_reg[0][26]  ( .D(n2175), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[0][26] ) );
  DFFR_X1 \DRAM_mem_reg[0][25]  ( .D(n2174), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[0][25] ) );
  DFFR_X1 \DRAM_mem_reg[0][24]  ( .D(n2173), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[0][24] ) );
  DFFR_X1 \DRAM_mem_reg[0][23]  ( .D(n2172), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[0][23] ) );
  DFFR_X1 \DRAM_mem_reg[0][22]  ( .D(n2171), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[0][22] ) );
  DFFR_X1 \DRAM_mem_reg[0][21]  ( .D(n2170), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[0][21] ) );
  DFFR_X1 \DRAM_mem_reg[0][20]  ( .D(n2169), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[0][20] ) );
  DFFR_X1 \DRAM_mem_reg[0][19]  ( .D(n2168), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[0][19] ) );
  DFFR_X1 \DRAM_mem_reg[0][18]  ( .D(n2167), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[0][18] ) );
  DFFR_X1 \DRAM_mem_reg[0][17]  ( .D(n2166), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[0][17] ) );
  DFFR_X1 \DRAM_mem_reg[0][16]  ( .D(n2165), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[0][16] ) );
  DFFR_X1 \DRAM_mem_reg[0][15]  ( .D(n2164), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[0][15] ) );
  DFFR_X1 \DRAM_mem_reg[0][14]  ( .D(n2163), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[0][14] ) );
  DFFR_X1 \DRAM_mem_reg[0][13]  ( .D(n2162), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[0][13] ) );
  DFFR_X1 \DRAM_mem_reg[0][12]  ( .D(n2161), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[0][12] ) );
  DFFR_X1 \DRAM_mem_reg[0][11]  ( .D(n2160), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[0][11] ) );
  DFFR_X1 \DRAM_mem_reg[0][10]  ( .D(n2159), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[0][10] ) );
  DFFR_X1 \DRAM_mem_reg[0][9]  ( .D(n2158), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[0][9] ) );
  DFFR_X1 \DRAM_mem_reg[0][8]  ( .D(n2157), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[0][8] ) );
  DFFR_X1 \DRAM_mem_reg[0][7]  ( .D(n2156), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[0][7] ) );
  DFFR_X1 \DRAM_mem_reg[0][6]  ( .D(n2155), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[0][6] ) );
  DFFR_X1 \DRAM_mem_reg[0][5]  ( .D(n2154), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[0][5] ) );
  DFFR_X1 \DRAM_mem_reg[0][4]  ( .D(n2153), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[0][4] ) );
  DFFR_X1 \DRAM_mem_reg[0][3]  ( .D(n2152), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[0][3] ) );
  DFFR_X1 \DRAM_mem_reg[0][2]  ( .D(n2151), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[0][2] ) );
  DFFR_X1 \DRAM_mem_reg[0][1]  ( .D(n2150), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[0][1] ) );
  DFFR_X1 \DRAM_mem_reg[0][0]  ( .D(n2149), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[0][0] ) );
  DFFR_X1 \DRAM_mem_reg[1][31]  ( .D(n2148), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[1][31] ) );
  DFFR_X1 \DRAM_mem_reg[1][30]  ( .D(n2147), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[1][30] ) );
  DFFR_X1 \DRAM_mem_reg[1][29]  ( .D(n2146), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[1][29] ) );
  DFFR_X1 \DRAM_mem_reg[1][28]  ( .D(n2145), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[1][28] ) );
  DFFR_X1 \DRAM_mem_reg[1][27]  ( .D(n2144), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[1][27] ) );
  DFFR_X1 \DRAM_mem_reg[1][26]  ( .D(n2143), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[1][26] ) );
  DFFR_X1 \DRAM_mem_reg[1][25]  ( .D(n2142), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[1][25] ) );
  DFFR_X1 \DRAM_mem_reg[1][24]  ( .D(n2141), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[1][24] ) );
  DFFR_X1 \DRAM_mem_reg[1][23]  ( .D(n2140), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[1][23] ) );
  DFFR_X1 \DRAM_mem_reg[1][22]  ( .D(n2139), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[1][22] ) );
  DFFR_X1 \DRAM_mem_reg[1][21]  ( .D(n2138), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[1][21] ) );
  DFFR_X1 \DRAM_mem_reg[1][20]  ( .D(n2137), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[1][20] ) );
  DFFR_X1 \DRAM_mem_reg[1][19]  ( .D(n2136), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[1][19] ) );
  DFFR_X1 \DRAM_mem_reg[1][18]  ( .D(n2135), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[1][18] ) );
  DFFR_X1 \DRAM_mem_reg[1][17]  ( .D(n2134), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[1][17] ) );
  DFFR_X1 \DRAM_mem_reg[1][16]  ( .D(n2133), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[1][16] ) );
  DFFR_X1 \DRAM_mem_reg[1][15]  ( .D(n2132), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[1][15] ) );
  DFFR_X1 \DRAM_mem_reg[1][14]  ( .D(n2131), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[1][14] ) );
  DFFR_X1 \DRAM_mem_reg[1][13]  ( .D(n2130), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[1][13] ) );
  DFFR_X1 \DRAM_mem_reg[1][12]  ( .D(n2129), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[1][12] ) );
  DFFR_X1 \DRAM_mem_reg[1][11]  ( .D(n2128), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[1][11] ) );
  DFFR_X1 \DRAM_mem_reg[1][10]  ( .D(n2127), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[1][10] ) );
  DFFR_X1 \DRAM_mem_reg[1][9]  ( .D(n2126), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[1][9] ) );
  DFFR_X1 \DRAM_mem_reg[1][8]  ( .D(n2125), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[1][8] ) );
  DFFR_X1 \DRAM_mem_reg[1][7]  ( .D(n2124), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[1][7] ) );
  DFFR_X1 \DRAM_mem_reg[1][6]  ( .D(n2123), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[1][6] ) );
  DFFR_X1 \DRAM_mem_reg[1][5]  ( .D(n2122), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[1][5] ) );
  DFFR_X1 \DRAM_mem_reg[1][4]  ( .D(n2121), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[1][4] ) );
  DFFR_X1 \DRAM_mem_reg[1][3]  ( .D(n2120), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[1][3] ) );
  DFFR_X1 \DRAM_mem_reg[1][2]  ( .D(n2119), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[1][2] ) );
  DFFR_X1 \DRAM_mem_reg[1][1]  ( .D(n2118), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[1][1] ) );
  DFFR_X1 \DRAM_mem_reg[1][0]  ( .D(n2117), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[1][0] ) );
  DFFR_X1 \DRAM_mem_reg[2][31]  ( .D(n2116), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[2][31] ) );
  DFFR_X1 \DRAM_mem_reg[2][30]  ( .D(n2115), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[2][30] ) );
  DFFR_X1 \DRAM_mem_reg[2][29]  ( .D(n2114), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[2][29] ) );
  DFFR_X1 \DRAM_mem_reg[2][28]  ( .D(n2113), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[2][28] ) );
  DFFR_X1 \DRAM_mem_reg[2][27]  ( .D(n2112), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[2][27] ) );
  DFFR_X1 \DRAM_mem_reg[2][26]  ( .D(n2111), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[2][26] ) );
  DFFR_X1 \DRAM_mem_reg[2][25]  ( .D(n2110), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[2][25] ) );
  DFFR_X1 \DRAM_mem_reg[2][24]  ( .D(n2109), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[2][24] ) );
  DFFR_X1 \DRAM_mem_reg[2][23]  ( .D(n2108), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[2][23] ) );
  DFFR_X1 \DRAM_mem_reg[2][22]  ( .D(n2107), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[2][22] ) );
  DFFR_X1 \DRAM_mem_reg[2][21]  ( .D(n2106), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[2][21] ) );
  DFFR_X1 \DRAM_mem_reg[2][20]  ( .D(n2105), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[2][20] ) );
  DFFR_X1 \DRAM_mem_reg[2][19]  ( .D(n2104), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[2][19] ) );
  DFFR_X1 \DRAM_mem_reg[2][18]  ( .D(n2103), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[2][18] ) );
  DFFR_X1 \DRAM_mem_reg[2][17]  ( .D(n2102), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[2][17] ) );
  DFFR_X1 \DRAM_mem_reg[2][16]  ( .D(n2101), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[2][16] ) );
  DFFR_X1 \DRAM_mem_reg[2][15]  ( .D(n2100), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[2][15] ) );
  DFFR_X1 \DRAM_mem_reg[2][14]  ( .D(n2099), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[2][14] ) );
  DFFR_X1 \DRAM_mem_reg[2][13]  ( .D(n2098), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[2][13] ) );
  DFFR_X1 \DRAM_mem_reg[2][12]  ( .D(n2097), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[2][12] ) );
  DFFR_X1 \DRAM_mem_reg[2][11]  ( .D(n2096), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[2][11] ) );
  DFFR_X1 \DRAM_mem_reg[2][10]  ( .D(n2095), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[2][10] ) );
  DFFR_X1 \DRAM_mem_reg[2][9]  ( .D(n2094), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[2][9] ) );
  DFFR_X1 \DRAM_mem_reg[2][8]  ( .D(n2093), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[2][8] ) );
  DFFR_X1 \DRAM_mem_reg[2][7]  ( .D(n2092), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[2][7] ) );
  DFFR_X1 \DRAM_mem_reg[2][6]  ( .D(n2091), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[2][6] ) );
  DFFR_X1 \DRAM_mem_reg[2][5]  ( .D(n2090), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[2][5] ) );
  DFFR_X1 \DRAM_mem_reg[2][4]  ( .D(n2089), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[2][4] ) );
  DFFR_X1 \DRAM_mem_reg[2][3]  ( .D(n2088), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[2][3] ) );
  DFFR_X1 \DRAM_mem_reg[2][2]  ( .D(n2087), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[2][2] ) );
  DFFR_X1 \DRAM_mem_reg[2][1]  ( .D(n2086), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[2][1] ) );
  DFFR_X1 \DRAM_mem_reg[2][0]  ( .D(n2085), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[2][0] ) );
  DFFR_X1 \DRAM_mem_reg[3][31]  ( .D(n2084), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[3][31] ) );
  DFFR_X1 \DRAM_mem_reg[3][30]  ( .D(n2083), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[3][30] ) );
  DFFR_X1 \DRAM_mem_reg[3][29]  ( .D(n2082), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[3][29] ) );
  DFFR_X1 \DRAM_mem_reg[3][28]  ( .D(n2081), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[3][28] ) );
  DFFR_X1 \DRAM_mem_reg[3][27]  ( .D(n2080), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[3][27] ) );
  DFFR_X1 \DRAM_mem_reg[3][26]  ( .D(n2079), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[3][26] ) );
  DFFR_X1 \DRAM_mem_reg[3][25]  ( .D(n2078), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[3][25] ) );
  DFFR_X1 \DRAM_mem_reg[3][24]  ( .D(n2077), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[3][24] ) );
  DFFR_X1 \DRAM_mem_reg[3][23]  ( .D(n2076), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[3][23] ) );
  DFFR_X1 \DRAM_mem_reg[3][22]  ( .D(n2075), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[3][22] ) );
  DFFR_X1 \DRAM_mem_reg[3][21]  ( .D(n2074), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[3][21] ) );
  DFFR_X1 \DRAM_mem_reg[3][20]  ( .D(n2073), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[3][20] ) );
  DFFR_X1 \DRAM_mem_reg[3][19]  ( .D(n2072), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[3][19] ) );
  DFFR_X1 \DRAM_mem_reg[3][18]  ( .D(n2071), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[3][18] ) );
  DFFR_X1 \DRAM_mem_reg[3][17]  ( .D(n2070), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[3][17] ) );
  DFFR_X1 \DRAM_mem_reg[3][16]  ( .D(n2069), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[3][16] ) );
  DFFR_X1 \DRAM_mem_reg[3][15]  ( .D(n2068), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[3][15] ) );
  DFFR_X1 \DRAM_mem_reg[3][14]  ( .D(n2067), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[3][14] ) );
  DFFR_X1 \DRAM_mem_reg[3][13]  ( .D(n2066), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[3][13] ) );
  DFFR_X1 \DRAM_mem_reg[3][12]  ( .D(n2065), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[3][12] ) );
  DFFR_X1 \DRAM_mem_reg[3][11]  ( .D(n2064), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[3][11] ) );
  DFFR_X1 \DRAM_mem_reg[3][10]  ( .D(n2063), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[3][10] ) );
  DFFR_X1 \DRAM_mem_reg[3][9]  ( .D(n2062), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[3][9] ) );
  DFFR_X1 \DRAM_mem_reg[3][8]  ( .D(n2061), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[3][8] ) );
  DFFR_X1 \DRAM_mem_reg[3][7]  ( .D(n2060), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[3][7] ) );
  DFFR_X1 \DRAM_mem_reg[3][6]  ( .D(n2059), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[3][6] ) );
  DFFR_X1 \DRAM_mem_reg[3][5]  ( .D(n2058), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[3][5] ) );
  DFFR_X1 \DRAM_mem_reg[3][4]  ( .D(n2057), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[3][4] ) );
  DFFR_X1 \DRAM_mem_reg[3][3]  ( .D(n2056), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[3][3] ) );
  DFFR_X1 \DRAM_mem_reg[3][2]  ( .D(n2055), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[3][2] ) );
  DFFR_X1 \DRAM_mem_reg[3][1]  ( .D(n2054), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[3][1] ) );
  DFFR_X1 \DRAM_mem_reg[3][0]  ( .D(n2053), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[3][0] ) );
  DFFR_X1 \DRAM_mem_reg[4][31]  ( .D(n2052), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[4][31] ) );
  DFFR_X1 \DRAM_mem_reg[4][30]  ( .D(n2051), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[4][30] ) );
  DFFR_X1 \DRAM_mem_reg[4][29]  ( .D(n2050), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[4][29] ) );
  DFFR_X1 \DRAM_mem_reg[4][28]  ( .D(n2049), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[4][28] ) );
  DFFR_X1 \DRAM_mem_reg[4][27]  ( .D(n2048), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[4][27] ) );
  DFFR_X1 \DRAM_mem_reg[4][26]  ( .D(n2047), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[4][26] ) );
  DFFR_X1 \DRAM_mem_reg[4][25]  ( .D(n2046), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[4][25] ) );
  DFFR_X1 \DRAM_mem_reg[4][24]  ( .D(n2045), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[4][24] ) );
  DFFR_X1 \DRAM_mem_reg[4][23]  ( .D(n2044), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[4][23] ) );
  DFFR_X1 \DRAM_mem_reg[4][22]  ( .D(n2043), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[4][22] ) );
  DFFR_X1 \DRAM_mem_reg[4][21]  ( .D(n2042), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[4][21] ) );
  DFFR_X1 \DRAM_mem_reg[4][20]  ( .D(n2041), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[4][20] ) );
  DFFR_X1 \DRAM_mem_reg[4][19]  ( .D(n2040), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[4][19] ) );
  DFFR_X1 \DRAM_mem_reg[4][18]  ( .D(n2039), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[4][18] ) );
  DFFR_X1 \DRAM_mem_reg[4][17]  ( .D(n2038), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[4][17] ) );
  DFFR_X1 \DRAM_mem_reg[4][16]  ( .D(n2037), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[4][16] ) );
  DFFR_X1 \DRAM_mem_reg[4][15]  ( .D(n2036), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[4][15] ) );
  DFFR_X1 \DRAM_mem_reg[4][14]  ( .D(n2035), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[4][14] ) );
  DFFR_X1 \DRAM_mem_reg[4][13]  ( .D(n2034), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[4][13] ) );
  DFFR_X1 \DRAM_mem_reg[4][12]  ( .D(n2033), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[4][12] ) );
  DFFR_X1 \DRAM_mem_reg[4][11]  ( .D(n2032), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[4][11] ) );
  DFFR_X1 \DRAM_mem_reg[4][10]  ( .D(n2031), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[4][10] ) );
  DFFR_X1 \DRAM_mem_reg[4][9]  ( .D(n2030), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[4][9] ) );
  DFFR_X1 \DRAM_mem_reg[4][8]  ( .D(n2029), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[4][8] ) );
  DFFR_X1 \DRAM_mem_reg[4][7]  ( .D(n2028), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[4][7] ) );
  DFFR_X1 \DRAM_mem_reg[4][6]  ( .D(n2027), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[4][6] ) );
  DFFR_X1 \DRAM_mem_reg[4][5]  ( .D(n2026), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[4][5] ) );
  DFFR_X1 \DRAM_mem_reg[4][4]  ( .D(n2025), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[4][4] ) );
  DFFR_X1 \DRAM_mem_reg[4][3]  ( .D(n2024), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[4][3] ) );
  DFFR_X1 \DRAM_mem_reg[4][2]  ( .D(n2023), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[4][2] ) );
  DFFR_X1 \DRAM_mem_reg[4][1]  ( .D(n2022), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[4][1] ) );
  DFFR_X1 \DRAM_mem_reg[4][0]  ( .D(n2021), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[4][0] ) );
  DFFR_X1 \DRAM_mem_reg[5][31]  ( .D(n2020), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[5][31] ) );
  DFFR_X1 \DRAM_mem_reg[5][30]  ( .D(n2019), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[5][30] ) );
  DFFR_X1 \DRAM_mem_reg[5][29]  ( .D(n2018), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[5][29] ) );
  DFFR_X1 \DRAM_mem_reg[5][28]  ( .D(n2017), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[5][28] ) );
  DFFR_X1 \DRAM_mem_reg[5][27]  ( .D(n2016), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[5][27] ) );
  DFFR_X1 \DRAM_mem_reg[5][26]  ( .D(n2015), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[5][26] ) );
  DFFR_X1 \DRAM_mem_reg[5][25]  ( .D(n2014), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[5][25] ) );
  DFFR_X1 \DRAM_mem_reg[5][24]  ( .D(n2013), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[5][24] ) );
  DFFR_X1 \DRAM_mem_reg[5][23]  ( .D(n2012), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[5][23] ) );
  DFFR_X1 \DRAM_mem_reg[5][22]  ( .D(n2011), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[5][22] ) );
  DFFR_X1 \DRAM_mem_reg[5][21]  ( .D(n2010), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[5][21] ) );
  DFFR_X1 \DRAM_mem_reg[5][20]  ( .D(n2009), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[5][20] ) );
  DFFR_X1 \DRAM_mem_reg[5][19]  ( .D(n2008), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[5][19] ) );
  DFFR_X1 \DRAM_mem_reg[5][18]  ( .D(n2007), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[5][18] ) );
  DFFR_X1 \DRAM_mem_reg[5][17]  ( .D(n2006), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[5][17] ) );
  DFFR_X1 \DRAM_mem_reg[5][16]  ( .D(n2005), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[5][16] ) );
  DFFR_X1 \DRAM_mem_reg[5][15]  ( .D(n2004), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[5][15] ) );
  DFFR_X1 \DRAM_mem_reg[5][14]  ( .D(n2003), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[5][14] ) );
  DFFR_X1 \DRAM_mem_reg[5][13]  ( .D(n2002), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[5][13] ) );
  DFFR_X1 \DRAM_mem_reg[5][12]  ( .D(n2001), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[5][12] ) );
  DFFR_X1 \DRAM_mem_reg[5][11]  ( .D(n2000), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[5][11] ) );
  DFFR_X1 \DRAM_mem_reg[5][10]  ( .D(n1999), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[5][10] ) );
  DFFR_X1 \DRAM_mem_reg[5][9]  ( .D(n1998), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[5][9] ) );
  DFFR_X1 \DRAM_mem_reg[5][8]  ( .D(n1997), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[5][8] ) );
  DFFR_X1 \DRAM_mem_reg[5][7]  ( .D(n1996), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[5][7] ) );
  DFFR_X1 \DRAM_mem_reg[5][6]  ( .D(n1995), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[5][6] ) );
  DFFR_X1 \DRAM_mem_reg[5][5]  ( .D(n1994), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[5][5] ) );
  DFFR_X1 \DRAM_mem_reg[5][4]  ( .D(n1993), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[5][4] ) );
  DFFR_X1 \DRAM_mem_reg[5][3]  ( .D(n1992), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[5][3] ) );
  DFFR_X1 \DRAM_mem_reg[5][2]  ( .D(n1991), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[5][2] ) );
  DFFR_X1 \DRAM_mem_reg[5][1]  ( .D(n1990), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[5][1] ) );
  DFFR_X1 \DRAM_mem_reg[5][0]  ( .D(n1989), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[5][0] ) );
  DFFR_X1 \DRAM_mem_reg[6][31]  ( .D(n1988), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[6][31] ) );
  DFFR_X1 \DRAM_mem_reg[6][30]  ( .D(n1987), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[6][30] ) );
  DFFR_X1 \DRAM_mem_reg[6][29]  ( .D(n1986), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[6][29] ) );
  DFFR_X1 \DRAM_mem_reg[6][28]  ( .D(n1985), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[6][28] ) );
  DFFR_X1 \DRAM_mem_reg[6][27]  ( .D(n1984), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[6][27] ) );
  DFFR_X1 \DRAM_mem_reg[6][26]  ( .D(n1983), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[6][26] ) );
  DFFR_X1 \DRAM_mem_reg[6][25]  ( .D(n1982), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[6][25] ) );
  DFFR_X1 \DRAM_mem_reg[6][24]  ( .D(n1981), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[6][24] ) );
  DFFR_X1 \DRAM_mem_reg[6][23]  ( .D(n1980), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[6][23] ) );
  DFFR_X1 \DRAM_mem_reg[6][22]  ( .D(n1979), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[6][22] ) );
  DFFR_X1 \DRAM_mem_reg[6][21]  ( .D(n1978), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[6][21] ) );
  DFFR_X1 \DRAM_mem_reg[6][20]  ( .D(n1977), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[6][20] ) );
  DFFR_X1 \DRAM_mem_reg[6][19]  ( .D(n1976), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[6][19] ) );
  DFFR_X1 \DRAM_mem_reg[6][18]  ( .D(n1975), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[6][18] ) );
  DFFR_X1 \DRAM_mem_reg[6][17]  ( .D(n1974), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[6][17] ) );
  DFFR_X1 \DRAM_mem_reg[6][16]  ( .D(n1973), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[6][16] ) );
  DFFR_X1 \DRAM_mem_reg[6][15]  ( .D(n1972), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[6][15] ) );
  DFFR_X1 \DRAM_mem_reg[6][14]  ( .D(n1971), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[6][14] ) );
  DFFR_X1 \DRAM_mem_reg[6][13]  ( .D(n1970), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[6][13] ) );
  DFFR_X1 \DRAM_mem_reg[6][12]  ( .D(n1969), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[6][12] ) );
  DFFR_X1 \DRAM_mem_reg[6][11]  ( .D(n1968), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[6][11] ) );
  DFFR_X1 \DRAM_mem_reg[6][10]  ( .D(n1967), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[6][10] ) );
  DFFR_X1 \DRAM_mem_reg[6][9]  ( .D(n1966), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[6][9] ) );
  DFFR_X1 \DRAM_mem_reg[6][8]  ( .D(n1965), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[6][8] ) );
  DFFR_X1 \DRAM_mem_reg[6][7]  ( .D(n1964), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[6][7] ) );
  DFFR_X1 \DRAM_mem_reg[6][6]  ( .D(n1963), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[6][6] ) );
  DFFR_X1 \DRAM_mem_reg[6][5]  ( .D(n1962), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[6][5] ) );
  DFFR_X1 \DRAM_mem_reg[6][4]  ( .D(n1961), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[6][4] ) );
  DFFR_X1 \DRAM_mem_reg[6][3]  ( .D(n1960), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[6][3] ) );
  DFFR_X1 \DRAM_mem_reg[6][2]  ( .D(n1959), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[6][2] ) );
  DFFR_X1 \DRAM_mem_reg[6][1]  ( .D(n1958), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[6][1] ) );
  DFFR_X1 \DRAM_mem_reg[6][0]  ( .D(n1957), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[6][0] ) );
  DFFR_X1 \DRAM_mem_reg[7][31]  ( .D(n1956), .CK(CLK), .RN(n86), .Q(
        \DRAM_mem[7][31] ) );
  DFFR_X1 \DRAM_mem_reg[7][30]  ( .D(n1955), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[7][30] ) );
  DFFR_X1 \DRAM_mem_reg[7][29]  ( .D(n1954), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[7][29] ) );
  DFFR_X1 \DRAM_mem_reg[7][28]  ( .D(n1953), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[7][28] ) );
  DFFR_X1 \DRAM_mem_reg[7][27]  ( .D(n1952), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[7][27] ) );
  DFFR_X1 \DRAM_mem_reg[7][26]  ( .D(n1951), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[7][26] ) );
  DFFR_X1 \DRAM_mem_reg[7][25]  ( .D(n1950), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[7][25] ) );
  DFFR_X1 \DRAM_mem_reg[7][24]  ( .D(n1949), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[7][24] ) );
  DFFR_X1 \DRAM_mem_reg[7][23]  ( .D(n1948), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[7][23] ) );
  DFFR_X1 \DRAM_mem_reg[7][22]  ( .D(n1947), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[7][22] ) );
  DFFR_X1 \DRAM_mem_reg[7][21]  ( .D(n1946), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[7][21] ) );
  DFFR_X1 \DRAM_mem_reg[7][20]  ( .D(n1945), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[7][20] ) );
  DFFR_X1 \DRAM_mem_reg[7][19]  ( .D(n1944), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[7][19] ) );
  DFFR_X1 \DRAM_mem_reg[7][18]  ( .D(n1943), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[7][18] ) );
  DFFR_X1 \DRAM_mem_reg[7][17]  ( .D(n1942), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[7][17] ) );
  DFFR_X1 \DRAM_mem_reg[7][16]  ( .D(n1941), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[7][16] ) );
  DFFR_X1 \DRAM_mem_reg[7][15]  ( .D(n1940), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[7][15] ) );
  DFFR_X1 \DRAM_mem_reg[7][14]  ( .D(n1939), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[7][14] ) );
  DFFR_X1 \DRAM_mem_reg[7][13]  ( .D(n1938), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[7][13] ) );
  DFFR_X1 \DRAM_mem_reg[7][12]  ( .D(n1937), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[7][12] ) );
  DFFR_X1 \DRAM_mem_reg[7][11]  ( .D(n1936), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[7][11] ) );
  DFFR_X1 \DRAM_mem_reg[7][10]  ( .D(n1935), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[7][10] ) );
  DFFR_X1 \DRAM_mem_reg[7][9]  ( .D(n1934), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[7][9] ) );
  DFFR_X1 \DRAM_mem_reg[7][8]  ( .D(n1933), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[7][8] ) );
  DFFR_X1 \DRAM_mem_reg[7][7]  ( .D(n1932), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[7][7] ) );
  DFFR_X1 \DRAM_mem_reg[7][6]  ( .D(n1931), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[7][6] ) );
  DFFR_X1 \DRAM_mem_reg[7][5]  ( .D(n1930), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[7][5] ) );
  DFFR_X1 \DRAM_mem_reg[7][4]  ( .D(n1929), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[7][4] ) );
  DFFR_X1 \DRAM_mem_reg[7][3]  ( .D(n1928), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[7][3] ) );
  DFFR_X1 \DRAM_mem_reg[7][2]  ( .D(n1927), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[7][2] ) );
  DFFR_X1 \DRAM_mem_reg[7][1]  ( .D(n1926), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[7][1] ) );
  DFFR_X1 \DRAM_mem_reg[7][0]  ( .D(n1925), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[7][0] ) );
  DFFR_X1 \DRAM_mem_reg[8][31]  ( .D(n1924), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[8][31] ) );
  DFFR_X1 \DRAM_mem_reg[8][30]  ( .D(n1923), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[8][30] ) );
  DFFR_X1 \DRAM_mem_reg[8][29]  ( .D(n1922), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[8][29] ) );
  DFFR_X1 \DRAM_mem_reg[8][28]  ( .D(n1921), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[8][28] ) );
  DFFR_X1 \DRAM_mem_reg[8][27]  ( .D(n1920), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[8][27] ) );
  DFFR_X1 \DRAM_mem_reg[8][26]  ( .D(n1919), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[8][26] ) );
  DFFR_X1 \DRAM_mem_reg[8][25]  ( .D(n1918), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[8][25] ) );
  DFFR_X1 \DRAM_mem_reg[8][24]  ( .D(n1917), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[8][24] ) );
  DFFR_X1 \DRAM_mem_reg[8][23]  ( .D(n1916), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[8][23] ) );
  DFFR_X1 \DRAM_mem_reg[8][22]  ( .D(n1915), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[8][22] ) );
  DFFR_X1 \DRAM_mem_reg[8][21]  ( .D(n1914), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[8][21] ) );
  DFFR_X1 \DRAM_mem_reg[8][20]  ( .D(n1913), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[8][20] ) );
  DFFR_X1 \DRAM_mem_reg[8][19]  ( .D(n1912), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[8][19] ) );
  DFFR_X1 \DRAM_mem_reg[8][18]  ( .D(n1911), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[8][18] ) );
  DFFR_X1 \DRAM_mem_reg[8][17]  ( .D(n1910), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[8][17] ) );
  DFFR_X1 \DRAM_mem_reg[8][16]  ( .D(n1909), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[8][16] ) );
  DFFR_X1 \DRAM_mem_reg[8][15]  ( .D(n1908), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[8][15] ) );
  DFFR_X1 \DRAM_mem_reg[8][14]  ( .D(n1907), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[8][14] ) );
  DFFR_X1 \DRAM_mem_reg[8][13]  ( .D(n1906), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[8][13] ) );
  DFFR_X1 \DRAM_mem_reg[8][12]  ( .D(n1905), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[8][12] ) );
  DFFR_X1 \DRAM_mem_reg[8][11]  ( .D(n1904), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[8][11] ) );
  DFFR_X1 \DRAM_mem_reg[8][10]  ( .D(n1903), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[8][10] ) );
  DFFR_X1 \DRAM_mem_reg[8][9]  ( .D(n1902), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[8][9] ) );
  DFFR_X1 \DRAM_mem_reg[8][8]  ( .D(n1901), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[8][8] ) );
  DFFR_X1 \DRAM_mem_reg[8][7]  ( .D(n1900), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[8][7] ) );
  DFFR_X1 \DRAM_mem_reg[8][6]  ( .D(n1899), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[8][6] ) );
  DFFR_X1 \DRAM_mem_reg[8][5]  ( .D(n1898), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[8][5] ) );
  DFFR_X1 \DRAM_mem_reg[8][4]  ( .D(n1897), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[8][4] ) );
  DFFR_X1 \DRAM_mem_reg[8][3]  ( .D(n1896), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[8][3] ) );
  DFFR_X1 \DRAM_mem_reg[8][2]  ( .D(n1895), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[8][2] ) );
  DFFR_X1 \DRAM_mem_reg[8][1]  ( .D(n1894), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[8][1] ) );
  DFFR_X1 \DRAM_mem_reg[8][0]  ( .D(n1893), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[8][0] ) );
  DFFR_X1 \DRAM_mem_reg[9][31]  ( .D(n1892), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[9][31] ) );
  DFFR_X1 \DRAM_mem_reg[9][30]  ( .D(n1891), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[9][30] ) );
  DFFR_X1 \DRAM_mem_reg[9][29]  ( .D(n1890), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[9][29] ) );
  DFFR_X1 \DRAM_mem_reg[9][28]  ( .D(n1889), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[9][28] ) );
  DFFR_X1 \DRAM_mem_reg[9][27]  ( .D(n1888), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[9][27] ) );
  DFFR_X1 \DRAM_mem_reg[9][26]  ( .D(n1887), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[9][26] ) );
  DFFR_X1 \DRAM_mem_reg[9][25]  ( .D(n1886), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[9][25] ) );
  DFFR_X1 \DRAM_mem_reg[9][24]  ( .D(n1885), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[9][24] ) );
  DFFR_X1 \DRAM_mem_reg[9][23]  ( .D(n1884), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[9][23] ) );
  DFFR_X1 \DRAM_mem_reg[9][22]  ( .D(n1883), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[9][22] ) );
  DFFR_X1 \DRAM_mem_reg[9][21]  ( .D(n1882), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[9][21] ) );
  DFFR_X1 \DRAM_mem_reg[9][20]  ( .D(n1881), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[9][20] ) );
  DFFR_X1 \DRAM_mem_reg[9][19]  ( .D(n1880), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[9][19] ) );
  DFFR_X1 \DRAM_mem_reg[9][18]  ( .D(n1879), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[9][18] ) );
  DFFR_X1 \DRAM_mem_reg[9][17]  ( .D(n1878), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[9][17] ) );
  DFFR_X1 \DRAM_mem_reg[9][16]  ( .D(n1877), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[9][16] ) );
  DFFR_X1 \DRAM_mem_reg[9][15]  ( .D(n1876), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[9][15] ) );
  DFFR_X1 \DRAM_mem_reg[9][14]  ( .D(n1875), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[9][14] ) );
  DFFR_X1 \DRAM_mem_reg[9][13]  ( .D(n1874), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[9][13] ) );
  DFFR_X1 \DRAM_mem_reg[9][12]  ( .D(n1873), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[9][12] ) );
  DFFR_X1 \DRAM_mem_reg[9][11]  ( .D(n1872), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[9][11] ) );
  DFFR_X1 \DRAM_mem_reg[9][10]  ( .D(n1871), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[9][10] ) );
  DFFR_X1 \DRAM_mem_reg[9][9]  ( .D(n1870), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[9][9] ) );
  DFFR_X1 \DRAM_mem_reg[9][8]  ( .D(n1869), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[9][8] ) );
  DFFR_X1 \DRAM_mem_reg[9][7]  ( .D(n1868), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[9][7] ) );
  DFFR_X1 \DRAM_mem_reg[9][6]  ( .D(n1867), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[9][6] ) );
  DFFR_X1 \DRAM_mem_reg[9][5]  ( .D(n1866), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[9][5] ) );
  DFFR_X1 \DRAM_mem_reg[9][4]  ( .D(n1865), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[9][4] ) );
  DFFR_X1 \DRAM_mem_reg[9][3]  ( .D(n1864), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[9][3] ) );
  DFFR_X1 \DRAM_mem_reg[9][2]  ( .D(n1863), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[9][2] ) );
  DFFR_X1 \DRAM_mem_reg[9][1]  ( .D(n1862), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[9][1] ) );
  DFFR_X1 \DRAM_mem_reg[9][0]  ( .D(n1861), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[9][0] ) );
  DFFR_X1 \DRAM_mem_reg[10][31]  ( .D(n1860), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[10][31] ) );
  DFFR_X1 \DRAM_mem_reg[10][30]  ( .D(n1859), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[10][30] ) );
  DFFR_X1 \DRAM_mem_reg[10][29]  ( .D(n1858), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[10][29] ) );
  DFFR_X1 \DRAM_mem_reg[10][28]  ( .D(n1857), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[10][28] ) );
  DFFR_X1 \DRAM_mem_reg[10][27]  ( .D(n1856), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[10][27] ) );
  DFFR_X1 \DRAM_mem_reg[10][26]  ( .D(n1855), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[10][26] ) );
  DFFR_X1 \DRAM_mem_reg[10][25]  ( .D(n1854), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[10][25] ) );
  DFFR_X1 \DRAM_mem_reg[10][24]  ( .D(n1853), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[10][24] ) );
  DFFR_X1 \DRAM_mem_reg[10][23]  ( .D(n1852), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[10][23] ) );
  DFFR_X1 \DRAM_mem_reg[10][22]  ( .D(n1851), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[10][22] ) );
  DFFR_X1 \DRAM_mem_reg[10][21]  ( .D(n1850), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[10][21] ) );
  DFFR_X1 \DRAM_mem_reg[10][20]  ( .D(n1849), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[10][20] ) );
  DFFR_X1 \DRAM_mem_reg[10][19]  ( .D(n1848), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[10][19] ) );
  DFFR_X1 \DRAM_mem_reg[10][18]  ( .D(n1847), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[10][18] ) );
  DFFR_X1 \DRAM_mem_reg[10][17]  ( .D(n1846), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[10][17] ) );
  DFFR_X1 \DRAM_mem_reg[10][16]  ( .D(n1845), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[10][16] ) );
  DFFR_X1 \DRAM_mem_reg[10][15]  ( .D(n1844), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[10][15] ) );
  DFFR_X1 \DRAM_mem_reg[10][14]  ( .D(n1843), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[10][14] ) );
  DFFR_X1 \DRAM_mem_reg[10][13]  ( .D(n1842), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[10][13] ) );
  DFFR_X1 \DRAM_mem_reg[10][12]  ( .D(n1841), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[10][12] ) );
  DFFR_X1 \DRAM_mem_reg[10][11]  ( .D(n1840), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[10][11] ) );
  DFFR_X1 \DRAM_mem_reg[10][10]  ( .D(n1839), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[10][10] ) );
  DFFR_X1 \DRAM_mem_reg[10][9]  ( .D(n1838), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[10][9] ) );
  DFFR_X1 \DRAM_mem_reg[10][8]  ( .D(n1837), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[10][8] ) );
  DFFR_X1 \DRAM_mem_reg[10][7]  ( .D(n1836), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[10][7] ) );
  DFFR_X1 \DRAM_mem_reg[10][6]  ( .D(n1835), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[10][6] ) );
  DFFR_X1 \DRAM_mem_reg[10][5]  ( .D(n1834), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[10][5] ) );
  DFFR_X1 \DRAM_mem_reg[10][4]  ( .D(n1833), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[10][4] ) );
  DFFR_X1 \DRAM_mem_reg[10][3]  ( .D(n1832), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[10][3] ) );
  DFFR_X1 \DRAM_mem_reg[10][2]  ( .D(n1831), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[10][2] ) );
  DFFR_X1 \DRAM_mem_reg[10][1]  ( .D(n1830), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[10][1] ) );
  DFFR_X1 \DRAM_mem_reg[10][0]  ( .D(n1829), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[10][0] ) );
  DFFR_X1 \DRAM_mem_reg[11][31]  ( .D(n1828), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[11][31] ) );
  DFFR_X1 \DRAM_mem_reg[11][30]  ( .D(n1827), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[11][30] ) );
  DFFR_X1 \DRAM_mem_reg[11][29]  ( .D(n1826), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[11][29] ) );
  DFFR_X1 \DRAM_mem_reg[11][28]  ( .D(n1825), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[11][28] ) );
  DFFR_X1 \DRAM_mem_reg[11][27]  ( .D(n1824), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[11][27] ) );
  DFFR_X1 \DRAM_mem_reg[11][26]  ( .D(n1823), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[11][26] ) );
  DFFR_X1 \DRAM_mem_reg[11][25]  ( .D(n1822), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[11][25] ) );
  DFFR_X1 \DRAM_mem_reg[11][24]  ( .D(n1821), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[11][24] ) );
  DFFR_X1 \DRAM_mem_reg[11][23]  ( .D(n1820), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[11][23] ) );
  DFFR_X1 \DRAM_mem_reg[11][22]  ( .D(n1819), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[11][22] ) );
  DFFR_X1 \DRAM_mem_reg[11][21]  ( .D(n1818), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[11][21] ) );
  DFFR_X1 \DRAM_mem_reg[11][20]  ( .D(n1817), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[11][20] ) );
  DFFR_X1 \DRAM_mem_reg[11][19]  ( .D(n1816), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[11][19] ) );
  DFFR_X1 \DRAM_mem_reg[11][18]  ( .D(n1815), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[11][18] ) );
  DFFR_X1 \DRAM_mem_reg[11][17]  ( .D(n1814), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[11][17] ) );
  DFFR_X1 \DRAM_mem_reg[11][16]  ( .D(n1813), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[11][16] ) );
  DFFR_X1 \DRAM_mem_reg[11][15]  ( .D(n1812), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[11][15] ) );
  DFFR_X1 \DRAM_mem_reg[11][14]  ( .D(n1811), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[11][14] ) );
  DFFR_X1 \DRAM_mem_reg[11][13]  ( .D(n1810), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[11][13] ) );
  DFFR_X1 \DRAM_mem_reg[11][12]  ( .D(n1809), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[11][12] ) );
  DFFR_X1 \DRAM_mem_reg[11][11]  ( .D(n1808), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[11][11] ) );
  DFFR_X1 \DRAM_mem_reg[11][10]  ( .D(n1807), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[11][10] ) );
  DFFR_X1 \DRAM_mem_reg[11][9]  ( .D(n1806), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[11][9] ) );
  DFFR_X1 \DRAM_mem_reg[11][8]  ( .D(n1805), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[11][8] ) );
  DFFR_X1 \DRAM_mem_reg[11][7]  ( .D(n1804), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[11][7] ) );
  DFFR_X1 \DRAM_mem_reg[11][6]  ( .D(n1803), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[11][6] ) );
  DFFR_X1 \DRAM_mem_reg[11][5]  ( .D(n1802), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[11][5] ) );
  DFFR_X1 \DRAM_mem_reg[11][4]  ( .D(n1801), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[11][4] ) );
  DFFR_X1 \DRAM_mem_reg[11][3]  ( .D(n1800), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[11][3] ) );
  DFFR_X1 \DRAM_mem_reg[11][2]  ( .D(n1799), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[11][2] ) );
  DFFR_X1 \DRAM_mem_reg[11][1]  ( .D(n1798), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[11][1] ) );
  DFFR_X1 \DRAM_mem_reg[11][0]  ( .D(n1797), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[11][0] ) );
  DFFR_X1 \DRAM_mem_reg[12][31]  ( .D(n1796), .CK(CLK), .RN(n1), .Q(
        \DRAM_mem[12][31] ) );
  DFFR_X1 \DRAM_mem_reg[12][30]  ( .D(n1795), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[12][30] ) );
  DFFR_X1 \DRAM_mem_reg[12][29]  ( .D(n1794), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[12][29] ) );
  DFFR_X1 \DRAM_mem_reg[12][28]  ( .D(n1793), .CK(CLK), .RN(n9), .Q(
        \DRAM_mem[12][28] ) );
  DFFR_X1 \DRAM_mem_reg[12][27]  ( .D(n1792), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[12][27] ) );
  DFFR_X1 \DRAM_mem_reg[12][26]  ( .D(n1791), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[12][26] ) );
  DFFR_X1 \DRAM_mem_reg[12][25]  ( .D(n1790), .CK(CLK), .RN(n17), .Q(
        \DRAM_mem[12][25] ) );
  DFFR_X1 \DRAM_mem_reg[12][24]  ( .D(n1789), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[12][24] ) );
  DFFR_X1 \DRAM_mem_reg[12][23]  ( .D(n1788), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[12][23] ) );
  DFFR_X1 \DRAM_mem_reg[12][22]  ( .D(n1787), .CK(CLK), .RN(n25), .Q(
        \DRAM_mem[12][22] ) );
  DFFR_X1 \DRAM_mem_reg[12][21]  ( .D(n1786), .CK(CLK), .RN(n33), .Q(
        \DRAM_mem[12][21] ) );
  DFFR_X1 \DRAM_mem_reg[12][20]  ( .D(n1785), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[12][20] ) );
  DFFR_X1 \DRAM_mem_reg[12][19]  ( .D(n1784), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[12][19] ) );
  DFFR_X1 \DRAM_mem_reg[12][18]  ( .D(n1783), .CK(CLK), .RN(n41), .Q(
        \DRAM_mem[12][18] ) );
  DFFR_X1 \DRAM_mem_reg[12][17]  ( .D(n1782), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[12][17] ) );
  DFFR_X1 \DRAM_mem_reg[12][16]  ( .D(n1781), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[12][16] ) );
  DFFR_X1 \DRAM_mem_reg[12][15]  ( .D(n1780), .CK(CLK), .RN(n49), .Q(
        \DRAM_mem[12][15] ) );
  DFFR_X1 \DRAM_mem_reg[12][14]  ( .D(n1779), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[12][14] ) );
  DFFR_X1 \DRAM_mem_reg[12][13]  ( .D(n1778), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[12][13] ) );
  DFFR_X1 \DRAM_mem_reg[12][12]  ( .D(n1777), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[12][12] ) );
  DFFR_X1 \DRAM_mem_reg[12][11]  ( .D(n1776), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[12][11] ) );
  DFFR_X1 \DRAM_mem_reg[12][10]  ( .D(n1775), .CK(CLK), .RN(n57), .Q(
        \DRAM_mem[12][10] ) );
  DFFR_X1 \DRAM_mem_reg[12][9]  ( .D(n1774), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[12][9] ) );
  DFFR_X1 \DRAM_mem_reg[12][8]  ( .D(n1773), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[12][8] ) );
  DFFR_X1 \DRAM_mem_reg[12][7]  ( .D(n1772), .CK(CLK), .RN(n81), .Q(
        \DRAM_mem[12][7] ) );
  DFFR_X1 \DRAM_mem_reg[12][6]  ( .D(n1771), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[12][6] ) );
  DFFR_X1 \DRAM_mem_reg[12][5]  ( .D(n1770), .CK(CLK), .RN(n73), .Q(
        \DRAM_mem[12][5] ) );
  DFFR_X1 \DRAM_mem_reg[12][4]  ( .D(n1769), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[12][4] ) );
  DFFR_X1 \DRAM_mem_reg[12][3]  ( .D(n1768), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[12][3] ) );
  DFFR_X1 \DRAM_mem_reg[12][2]  ( .D(n1767), .CK(CLK), .RN(n65), .Q(
        \DRAM_mem[12][2] ) );
  DFFR_X1 \DRAM_mem_reg[12][1]  ( .D(n1766), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[12][1] ) );
  DFFR_X1 \DRAM_mem_reg[12][0]  ( .D(n1765), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[12][0] ) );
  DFFR_X1 \DRAM_mem_reg[13][31]  ( .D(n1764), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[13][31] ) );
  DFFR_X1 \DRAM_mem_reg[13][30]  ( .D(n1763), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[13][30] ) );
  DFFR_X1 \DRAM_mem_reg[13][29]  ( .D(n1762), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[13][29] ) );
  DFFR_X1 \DRAM_mem_reg[13][28]  ( .D(n1761), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[13][28] ) );
  DFFR_X1 \DRAM_mem_reg[13][27]  ( .D(n1760), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[13][27] ) );
  DFFR_X1 \DRAM_mem_reg[13][26]  ( .D(n1759), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[13][26] ) );
  DFFR_X1 \DRAM_mem_reg[13][25]  ( .D(n1758), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[13][25] ) );
  DFFR_X1 \DRAM_mem_reg[13][24]  ( .D(n1757), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[13][24] ) );
  DFFR_X1 \DRAM_mem_reg[13][23]  ( .D(n1756), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[13][23] ) );
  DFFR_X1 \DRAM_mem_reg[13][22]  ( .D(n1755), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[13][22] ) );
  DFFR_X1 \DRAM_mem_reg[13][21]  ( .D(n1754), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[13][21] ) );
  DFFR_X1 \DRAM_mem_reg[13][20]  ( .D(n1753), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[13][20] ) );
  DFFR_X1 \DRAM_mem_reg[13][19]  ( .D(n1752), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[13][19] ) );
  DFFR_X1 \DRAM_mem_reg[13][18]  ( .D(n1751), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[13][18] ) );
  DFFR_X1 \DRAM_mem_reg[13][17]  ( .D(n1750), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[13][17] ) );
  DFFR_X1 \DRAM_mem_reg[13][16]  ( .D(n1749), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[13][16] ) );
  DFFR_X1 \DRAM_mem_reg[13][15]  ( .D(n1748), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[13][15] ) );
  DFFR_X1 \DRAM_mem_reg[13][14]  ( .D(n1747), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[13][14] ) );
  DFFR_X1 \DRAM_mem_reg[13][13]  ( .D(n1746), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[13][13] ) );
  DFFR_X1 \DRAM_mem_reg[13][12]  ( .D(n1745), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[13][12] ) );
  DFFR_X1 \DRAM_mem_reg[13][11]  ( .D(n1744), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[13][11] ) );
  DFFR_X1 \DRAM_mem_reg[13][10]  ( .D(n1743), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[13][10] ) );
  DFFR_X1 \DRAM_mem_reg[13][9]  ( .D(n1742), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[13][9] ) );
  DFFR_X1 \DRAM_mem_reg[13][8]  ( .D(n1741), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[13][8] ) );
  DFFR_X1 \DRAM_mem_reg[13][7]  ( .D(n1740), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[13][7] ) );
  DFFR_X1 \DRAM_mem_reg[13][6]  ( .D(n1739), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[13][6] ) );
  DFFR_X1 \DRAM_mem_reg[13][5]  ( .D(n1738), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[13][5] ) );
  DFFR_X1 \DRAM_mem_reg[13][4]  ( .D(n1737), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[13][4] ) );
  DFFR_X1 \DRAM_mem_reg[13][3]  ( .D(n1736), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[13][3] ) );
  DFFR_X1 \DRAM_mem_reg[13][2]  ( .D(n1735), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[13][2] ) );
  DFFR_X1 \DRAM_mem_reg[13][1]  ( .D(n1734), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[13][1] ) );
  DFFR_X1 \DRAM_mem_reg[13][0]  ( .D(n1733), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[13][0] ) );
  DFFR_X1 \DRAM_mem_reg[14][31]  ( .D(n1732), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[14][31] ) );
  DFFR_X1 \DRAM_mem_reg[14][30]  ( .D(n1731), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[14][30] ) );
  DFFR_X1 \DRAM_mem_reg[14][29]  ( .D(n1730), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[14][29] ) );
  DFFR_X1 \DRAM_mem_reg[14][28]  ( .D(n1729), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[14][28] ) );
  DFFR_X1 \DRAM_mem_reg[14][27]  ( .D(n1728), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[14][27] ) );
  DFFR_X1 \DRAM_mem_reg[14][26]  ( .D(n1727), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[14][26] ) );
  DFFR_X1 \DRAM_mem_reg[14][25]  ( .D(n1726), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[14][25] ) );
  DFFR_X1 \DRAM_mem_reg[14][24]  ( .D(n1725), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[14][24] ) );
  DFFR_X1 \DRAM_mem_reg[14][23]  ( .D(n1724), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[14][23] ) );
  DFFR_X1 \DRAM_mem_reg[14][22]  ( .D(n1723), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[14][22] ) );
  DFFR_X1 \DRAM_mem_reg[14][21]  ( .D(n1722), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[14][21] ) );
  DFFR_X1 \DRAM_mem_reg[14][20]  ( .D(n1721), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[14][20] ) );
  DFFR_X1 \DRAM_mem_reg[14][19]  ( .D(n1720), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[14][19] ) );
  DFFR_X1 \DRAM_mem_reg[14][18]  ( .D(n1719), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[14][18] ) );
  DFFR_X1 \DRAM_mem_reg[14][17]  ( .D(n1718), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[14][17] ) );
  DFFR_X1 \DRAM_mem_reg[14][16]  ( .D(n1717), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[14][16] ) );
  DFFR_X1 \DRAM_mem_reg[14][15]  ( .D(n1716), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[14][15] ) );
  DFFR_X1 \DRAM_mem_reg[14][14]  ( .D(n1715), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[14][14] ) );
  DFFR_X1 \DRAM_mem_reg[14][13]  ( .D(n1714), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[14][13] ) );
  DFFR_X1 \DRAM_mem_reg[14][12]  ( .D(n1713), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[14][12] ) );
  DFFR_X1 \DRAM_mem_reg[14][11]  ( .D(n1712), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[14][11] ) );
  DFFR_X1 \DRAM_mem_reg[14][10]  ( .D(n1711), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[14][10] ) );
  DFFR_X1 \DRAM_mem_reg[14][9]  ( .D(n1710), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[14][9] ) );
  DFFR_X1 \DRAM_mem_reg[14][8]  ( .D(n1709), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[14][8] ) );
  DFFR_X1 \DRAM_mem_reg[14][7]  ( .D(n1708), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[14][7] ) );
  DFFR_X1 \DRAM_mem_reg[14][6]  ( .D(n1707), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[14][6] ) );
  DFFR_X1 \DRAM_mem_reg[14][5]  ( .D(n1706), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[14][5] ) );
  DFFR_X1 \DRAM_mem_reg[14][4]  ( .D(n1705), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[14][4] ) );
  DFFR_X1 \DRAM_mem_reg[14][3]  ( .D(n1704), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[14][3] ) );
  DFFR_X1 \DRAM_mem_reg[14][2]  ( .D(n1703), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[14][2] ) );
  DFFR_X1 \DRAM_mem_reg[14][1]  ( .D(n1702), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[14][1] ) );
  DFFR_X1 \DRAM_mem_reg[14][0]  ( .D(n1701), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[14][0] ) );
  DFFR_X1 \DRAM_mem_reg[15][31]  ( .D(n1700), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[15][31] ) );
  DFFR_X1 \DRAM_mem_reg[15][30]  ( .D(n1699), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[15][30] ) );
  DFFR_X1 \DRAM_mem_reg[15][29]  ( .D(n1698), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[15][29] ) );
  DFFR_X1 \DRAM_mem_reg[15][28]  ( .D(n1697), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[15][28] ) );
  DFFR_X1 \DRAM_mem_reg[15][27]  ( .D(n1696), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[15][27] ) );
  DFFR_X1 \DRAM_mem_reg[15][26]  ( .D(n1695), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[15][26] ) );
  DFFR_X1 \DRAM_mem_reg[15][25]  ( .D(n1694), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[15][25] ) );
  DFFR_X1 \DRAM_mem_reg[15][24]  ( .D(n1693), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[15][24] ) );
  DFFR_X1 \DRAM_mem_reg[15][23]  ( .D(n1692), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[15][23] ) );
  DFFR_X1 \DRAM_mem_reg[15][22]  ( .D(n1691), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[15][22] ) );
  DFFR_X1 \DRAM_mem_reg[15][21]  ( .D(n1690), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[15][21] ) );
  DFFR_X1 \DRAM_mem_reg[15][20]  ( .D(n1689), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[15][20] ) );
  DFFR_X1 \DRAM_mem_reg[15][19]  ( .D(n1688), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[15][19] ) );
  DFFR_X1 \DRAM_mem_reg[15][18]  ( .D(n1687), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[15][18] ) );
  DFFR_X1 \DRAM_mem_reg[15][17]  ( .D(n1686), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[15][17] ) );
  DFFR_X1 \DRAM_mem_reg[15][16]  ( .D(n1685), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[15][16] ) );
  DFFR_X1 \DRAM_mem_reg[15][15]  ( .D(n1684), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[15][15] ) );
  DFFR_X1 \DRAM_mem_reg[15][14]  ( .D(n1683), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[15][14] ) );
  DFFR_X1 \DRAM_mem_reg[15][13]  ( .D(n1682), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[15][13] ) );
  DFFR_X1 \DRAM_mem_reg[15][12]  ( .D(n1681), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[15][12] ) );
  DFFR_X1 \DRAM_mem_reg[15][11]  ( .D(n1680), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[15][11] ) );
  DFFR_X1 \DRAM_mem_reg[15][10]  ( .D(n1679), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[15][10] ) );
  DFFR_X1 \DRAM_mem_reg[15][9]  ( .D(n1678), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[15][9] ) );
  DFFR_X1 \DRAM_mem_reg[15][8]  ( .D(n1677), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[15][8] ) );
  DFFR_X1 \DRAM_mem_reg[15][7]  ( .D(n1676), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[15][7] ) );
  DFFR_X1 \DRAM_mem_reg[15][6]  ( .D(n1675), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[15][6] ) );
  DFFR_X1 \DRAM_mem_reg[15][5]  ( .D(n1674), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[15][5] ) );
  DFFR_X1 \DRAM_mem_reg[15][4]  ( .D(n1673), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[15][4] ) );
  DFFR_X1 \DRAM_mem_reg[15][3]  ( .D(n1672), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[15][3] ) );
  DFFR_X1 \DRAM_mem_reg[15][2]  ( .D(n1671), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[15][2] ) );
  DFFR_X1 \DRAM_mem_reg[15][1]  ( .D(n1670), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[15][1] ) );
  DFFR_X1 \DRAM_mem_reg[15][0]  ( .D(n1669), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[15][0] ) );
  DFFR_X1 \DRAM_mem_reg[16][31]  ( .D(n1668), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[16][31] ) );
  DFFR_X1 \DRAM_mem_reg[16][30]  ( .D(n1667), .CK(CLK), .RN(n4), .Q(
        \DRAM_mem[16][30] ) );
  DFFR_X1 \DRAM_mem_reg[16][29]  ( .D(n1666), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[16][29] ) );
  DFFR_X1 \DRAM_mem_reg[16][28]  ( .D(n1665), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[16][28] ) );
  DFFR_X1 \DRAM_mem_reg[16][27]  ( .D(n1664), .CK(CLK), .RN(n12), .Q(
        \DRAM_mem[16][27] ) );
  DFFR_X1 \DRAM_mem_reg[16][26]  ( .D(n1663), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[16][26] ) );
  DFFR_X1 \DRAM_mem_reg[16][25]  ( .D(n1662), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[16][25] ) );
  DFFR_X1 \DRAM_mem_reg[16][24]  ( .D(n1661), .CK(CLK), .RN(n20), .Q(
        \DRAM_mem[16][24] ) );
  DFFR_X1 \DRAM_mem_reg[16][23]  ( .D(n1660), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[16][23] ) );
  DFFR_X1 \DRAM_mem_reg[16][22]  ( .D(n1659), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[16][22] ) );
  DFFR_X1 \DRAM_mem_reg[16][21]  ( .D(n1658), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[16][21] ) );
  DFFR_X1 \DRAM_mem_reg[16][20]  ( .D(n1657), .CK(CLK), .RN(n36), .Q(
        \DRAM_mem[16][20] ) );
  DFFR_X1 \DRAM_mem_reg[16][19]  ( .D(n1656), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[16][19] ) );
  DFFR_X1 \DRAM_mem_reg[16][18]  ( .D(n1655), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[16][18] ) );
  DFFR_X1 \DRAM_mem_reg[16][17]  ( .D(n1654), .CK(CLK), .RN(n44), .Q(
        \DRAM_mem[16][17] ) );
  DFFR_X1 \DRAM_mem_reg[16][16]  ( .D(n1653), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[16][16] ) );
  DFFR_X1 \DRAM_mem_reg[16][15]  ( .D(n1652), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[16][15] ) );
  DFFR_X1 \DRAM_mem_reg[16][14]  ( .D(n1651), .CK(CLK), .RN(n52), .Q(
        \DRAM_mem[16][14] ) );
  DFFR_X1 \DRAM_mem_reg[16][13]  ( .D(n1650), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[16][13] ) );
  DFFR_X1 \DRAM_mem_reg[16][12]  ( .D(n1649), .CK(CLK), .RN(n28), .Q(
        \DRAM_mem[16][12] ) );
  DFFR_X1 \DRAM_mem_reg[16][11]  ( .D(n1648), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[16][11] ) );
  DFFR_X1 \DRAM_mem_reg[16][10]  ( .D(n1647), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[16][10] ) );
  DFFR_X1 \DRAM_mem_reg[16][9]  ( .D(n1646), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[16][9] ) );
  DFFR_X1 \DRAM_mem_reg[16][8]  ( .D(n1645), .CK(CLK), .RN(n84), .Q(
        \DRAM_mem[16][8] ) );
  DFFR_X1 \DRAM_mem_reg[16][7]  ( .D(n1644), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[16][7] ) );
  DFFR_X1 \DRAM_mem_reg[16][6]  ( .D(n1643), .CK(CLK), .RN(n76), .Q(
        \DRAM_mem[16][6] ) );
  DFFR_X1 \DRAM_mem_reg[16][5]  ( .D(n1642), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[16][5] ) );
  DFFR_X1 \DRAM_mem_reg[16][4]  ( .D(n1641), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[16][4] ) );
  DFFR_X1 \DRAM_mem_reg[16][3]  ( .D(n1640), .CK(CLK), .RN(n68), .Q(
        \DRAM_mem[16][3] ) );
  DFFR_X1 \DRAM_mem_reg[16][2]  ( .D(n1639), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[16][2] ) );
  DFFR_X1 \DRAM_mem_reg[16][1]  ( .D(n1638), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[16][1] ) );
  DFFR_X1 \DRAM_mem_reg[16][0]  ( .D(n1637), .CK(CLK), .RN(n60), .Q(
        \DRAM_mem[16][0] ) );
  DFFR_X1 \DRAM_mem_reg[17][31]  ( .D(n1636), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[17][31] ) );
  DFFR_X1 \DRAM_mem_reg[17][30]  ( .D(n1635), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[17][30] ) );
  DFFR_X1 \DRAM_mem_reg[17][29]  ( .D(n1634), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[17][29] ) );
  DFFR_X1 \DRAM_mem_reg[17][28]  ( .D(n1633), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[17][28] ) );
  DFFR_X1 \DRAM_mem_reg[17][27]  ( .D(n1632), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[17][27] ) );
  DFFR_X1 \DRAM_mem_reg[17][26]  ( .D(n1631), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[17][26] ) );
  DFFR_X1 \DRAM_mem_reg[17][25]  ( .D(n1630), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[17][25] ) );
  DFFR_X1 \DRAM_mem_reg[17][24]  ( .D(n1629), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[17][24] ) );
  DFFR_X1 \DRAM_mem_reg[17][23]  ( .D(n1628), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[17][23] ) );
  DFFR_X1 \DRAM_mem_reg[17][22]  ( .D(n1627), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[17][22] ) );
  DFFR_X1 \DRAM_mem_reg[17][21]  ( .D(n1626), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[17][21] ) );
  DFFR_X1 \DRAM_mem_reg[17][20]  ( .D(n1625), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[17][20] ) );
  DFFR_X1 \DRAM_mem_reg[17][19]  ( .D(n1624), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[17][19] ) );
  DFFR_X1 \DRAM_mem_reg[17][18]  ( .D(n1623), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[17][18] ) );
  DFFR_X1 \DRAM_mem_reg[17][17]  ( .D(n1622), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[17][17] ) );
  DFFR_X1 \DRAM_mem_reg[17][16]  ( .D(n1621), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[17][16] ) );
  DFFR_X1 \DRAM_mem_reg[17][15]  ( .D(n1620), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[17][15] ) );
  DFFR_X1 \DRAM_mem_reg[17][14]  ( .D(n1619), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[17][14] ) );
  DFFR_X1 \DRAM_mem_reg[17][13]  ( .D(n1618), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[17][13] ) );
  DFFR_X1 \DRAM_mem_reg[17][12]  ( .D(n1617), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[17][12] ) );
  DFFR_X1 \DRAM_mem_reg[17][11]  ( .D(n1616), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[17][11] ) );
  DFFR_X1 \DRAM_mem_reg[17][10]  ( .D(n1615), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[17][10] ) );
  DFFR_X1 \DRAM_mem_reg[17][9]  ( .D(n1614), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[17][9] ) );
  DFFR_X1 \DRAM_mem_reg[17][8]  ( .D(n1613), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[17][8] ) );
  DFFR_X1 \DRAM_mem_reg[17][7]  ( .D(n1612), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[17][7] ) );
  DFFR_X1 \DRAM_mem_reg[17][6]  ( .D(n1611), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[17][6] ) );
  DFFR_X1 \DRAM_mem_reg[17][5]  ( .D(n1610), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[17][5] ) );
  DFFR_X1 \DRAM_mem_reg[17][4]  ( .D(n1609), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[17][4] ) );
  DFFR_X1 \DRAM_mem_reg[17][3]  ( .D(n1608), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[17][3] ) );
  DFFR_X1 \DRAM_mem_reg[17][2]  ( .D(n1607), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[17][2] ) );
  DFFR_X1 \DRAM_mem_reg[17][1]  ( .D(n1606), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[17][1] ) );
  DFFR_X1 \DRAM_mem_reg[17][0]  ( .D(n1605), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[17][0] ) );
  DFFR_X1 \DRAM_mem_reg[18][31]  ( .D(n1604), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[18][31] ) );
  DFFR_X1 \DRAM_mem_reg[18][30]  ( .D(n1603), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[18][30] ) );
  DFFR_X1 \DRAM_mem_reg[18][29]  ( .D(n1602), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[18][29] ) );
  DFFR_X1 \DRAM_mem_reg[18][28]  ( .D(n1601), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[18][28] ) );
  DFFR_X1 \DRAM_mem_reg[18][27]  ( .D(n1600), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[18][27] ) );
  DFFR_X1 \DRAM_mem_reg[18][26]  ( .D(n1599), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[18][26] ) );
  DFFR_X1 \DRAM_mem_reg[18][25]  ( .D(n1598), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[18][25] ) );
  DFFR_X1 \DRAM_mem_reg[18][24]  ( .D(n1597), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[18][24] ) );
  DFFR_X1 \DRAM_mem_reg[18][23]  ( .D(n1596), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[18][23] ) );
  DFFR_X1 \DRAM_mem_reg[18][22]  ( .D(n1595), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[18][22] ) );
  DFFR_X1 \DRAM_mem_reg[18][21]  ( .D(n1594), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[18][21] ) );
  DFFR_X1 \DRAM_mem_reg[18][20]  ( .D(n1593), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[18][20] ) );
  DFFR_X1 \DRAM_mem_reg[18][19]  ( .D(n1592), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[18][19] ) );
  DFFR_X1 \DRAM_mem_reg[18][18]  ( .D(n1591), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[18][18] ) );
  DFFR_X1 \DRAM_mem_reg[18][17]  ( .D(n1590), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[18][17] ) );
  DFFR_X1 \DRAM_mem_reg[18][16]  ( .D(n1589), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[18][16] ) );
  DFFR_X1 \DRAM_mem_reg[18][15]  ( .D(n1588), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[18][15] ) );
  DFFR_X1 \DRAM_mem_reg[18][14]  ( .D(n1587), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[18][14] ) );
  DFFR_X1 \DRAM_mem_reg[18][13]  ( .D(n1586), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[18][13] ) );
  DFFR_X1 \DRAM_mem_reg[18][12]  ( .D(n1585), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[18][12] ) );
  DFFR_X1 \DRAM_mem_reg[18][11]  ( .D(n1584), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[18][11] ) );
  DFFR_X1 \DRAM_mem_reg[18][10]  ( .D(n1583), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[18][10] ) );
  DFFR_X1 \DRAM_mem_reg[18][9]  ( .D(n1582), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[18][9] ) );
  DFFR_X1 \DRAM_mem_reg[18][8]  ( .D(n1581), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[18][8] ) );
  DFFR_X1 \DRAM_mem_reg[18][7]  ( .D(n1580), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[18][7] ) );
  DFFR_X1 \DRAM_mem_reg[18][6]  ( .D(n1579), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[18][6] ) );
  DFFR_X1 \DRAM_mem_reg[18][5]  ( .D(n1578), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[18][5] ) );
  DFFR_X1 \DRAM_mem_reg[18][4]  ( .D(n1577), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[18][4] ) );
  DFFR_X1 \DRAM_mem_reg[18][3]  ( .D(n1576), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[18][3] ) );
  DFFR_X1 \DRAM_mem_reg[18][2]  ( .D(n1575), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[18][2] ) );
  DFFR_X1 \DRAM_mem_reg[18][1]  ( .D(n1574), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[18][1] ) );
  DFFR_X1 \DRAM_mem_reg[18][0]  ( .D(n1573), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[18][0] ) );
  DFFR_X1 \DRAM_mem_reg[19][31]  ( .D(n1572), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[19][31] ) );
  DFFR_X1 \DRAM_mem_reg[19][30]  ( .D(n1571), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[19][30] ) );
  DFFR_X1 \DRAM_mem_reg[19][29]  ( .D(n1570), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[19][29] ) );
  DFFR_X1 \DRAM_mem_reg[19][28]  ( .D(n1569), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[19][28] ) );
  DFFR_X1 \DRAM_mem_reg[19][27]  ( .D(n1568), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[19][27] ) );
  DFFR_X1 \DRAM_mem_reg[19][26]  ( .D(n1567), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[19][26] ) );
  DFFR_X1 \DRAM_mem_reg[19][25]  ( .D(n1566), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[19][25] ) );
  DFFR_X1 \DRAM_mem_reg[19][24]  ( .D(n1565), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[19][24] ) );
  DFFR_X1 \DRAM_mem_reg[19][23]  ( .D(n1564), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[19][23] ) );
  DFFR_X1 \DRAM_mem_reg[19][22]  ( .D(n1563), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[19][22] ) );
  DFFR_X1 \DRAM_mem_reg[19][21]  ( .D(n1562), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[19][21] ) );
  DFFR_X1 \DRAM_mem_reg[19][20]  ( .D(n1561), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[19][20] ) );
  DFFR_X1 \DRAM_mem_reg[19][19]  ( .D(n1560), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[19][19] ) );
  DFFR_X1 \DRAM_mem_reg[19][18]  ( .D(n1559), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[19][18] ) );
  DFFR_X1 \DRAM_mem_reg[19][17]  ( .D(n1558), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[19][17] ) );
  DFFR_X1 \DRAM_mem_reg[19][16]  ( .D(n1557), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[19][16] ) );
  DFFR_X1 \DRAM_mem_reg[19][15]  ( .D(n1556), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[19][15] ) );
  DFFR_X1 \DRAM_mem_reg[19][14]  ( .D(n1555), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[19][14] ) );
  DFFR_X1 \DRAM_mem_reg[19][13]  ( .D(n1554), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[19][13] ) );
  DFFR_X1 \DRAM_mem_reg[19][12]  ( .D(n1553), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[19][12] ) );
  DFFR_X1 \DRAM_mem_reg[19][11]  ( .D(n1552), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[19][11] ) );
  DFFR_X1 \DRAM_mem_reg[19][10]  ( .D(n1551), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[19][10] ) );
  DFFR_X1 \DRAM_mem_reg[19][9]  ( .D(n1550), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[19][9] ) );
  DFFR_X1 \DRAM_mem_reg[19][8]  ( .D(n1549), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[19][8] ) );
  DFFR_X1 \DRAM_mem_reg[19][7]  ( .D(n1548), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[19][7] ) );
  DFFR_X1 \DRAM_mem_reg[19][6]  ( .D(n1547), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[19][6] ) );
  DFFR_X1 \DRAM_mem_reg[19][5]  ( .D(n1546), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[19][5] ) );
  DFFR_X1 \DRAM_mem_reg[19][4]  ( .D(n1545), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[19][4] ) );
  DFFR_X1 \DRAM_mem_reg[19][3]  ( .D(n1544), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[19][3] ) );
  DFFR_X1 \DRAM_mem_reg[19][2]  ( .D(n1543), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[19][2] ) );
  DFFR_X1 \DRAM_mem_reg[19][1]  ( .D(n1542), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[19][1] ) );
  DFFR_X1 \DRAM_mem_reg[19][0]  ( .D(n1541), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[19][0] ) );
  DFFR_X1 \DRAM_mem_reg[20][31]  ( .D(n1540), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[20][31] ) );
  DFFR_X1 \DRAM_mem_reg[20][30]  ( .D(n1539), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[20][30] ) );
  DFFR_X1 \DRAM_mem_reg[20][29]  ( .D(n1538), .CK(CLK), .RN(n7), .Q(
        \DRAM_mem[20][29] ) );
  DFFR_X1 \DRAM_mem_reg[20][28]  ( .D(n1537), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[20][28] ) );
  DFFR_X1 \DRAM_mem_reg[20][27]  ( .D(n1536), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[20][27] ) );
  DFFR_X1 \DRAM_mem_reg[20][26]  ( .D(n1535), .CK(CLK), .RN(n15), .Q(
        \DRAM_mem[20][26] ) );
  DFFR_X1 \DRAM_mem_reg[20][25]  ( .D(n1534), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[20][25] ) );
  DFFR_X1 \DRAM_mem_reg[20][24]  ( .D(n1533), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[20][24] ) );
  DFFR_X1 \DRAM_mem_reg[20][23]  ( .D(n1532), .CK(CLK), .RN(n23), .Q(
        \DRAM_mem[20][23] ) );
  DFFR_X1 \DRAM_mem_reg[20][22]  ( .D(n1531), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[20][22] ) );
  DFFR_X1 \DRAM_mem_reg[20][21]  ( .D(n1530), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[20][21] ) );
  DFFR_X1 \DRAM_mem_reg[20][20]  ( .D(n1529), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[20][20] ) );
  DFFR_X1 \DRAM_mem_reg[20][19]  ( .D(n1528), .CK(CLK), .RN(n39), .Q(
        \DRAM_mem[20][19] ) );
  DFFR_X1 \DRAM_mem_reg[20][18]  ( .D(n1527), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[20][18] ) );
  DFFR_X1 \DRAM_mem_reg[20][17]  ( .D(n1526), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[20][17] ) );
  DFFR_X1 \DRAM_mem_reg[20][16]  ( .D(n1525), .CK(CLK), .RN(n47), .Q(
        \DRAM_mem[20][16] ) );
  DFFR_X1 \DRAM_mem_reg[20][15]  ( .D(n1524), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[20][15] ) );
  DFFR_X1 \DRAM_mem_reg[20][14]  ( .D(n1523), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[20][14] ) );
  DFFR_X1 \DRAM_mem_reg[20][13]  ( .D(n1522), .CK(CLK), .RN(n31), .Q(
        \DRAM_mem[20][13] ) );
  DFFR_X1 \DRAM_mem_reg[20][12]  ( .D(n1521), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[20][12] ) );
  DFFR_X1 \DRAM_mem_reg[20][11]  ( .D(n1520), .CK(CLK), .RN(n55), .Q(
        \DRAM_mem[20][11] ) );
  DFFR_X1 \DRAM_mem_reg[20][10]  ( .D(n1519), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[20][10] ) );
  DFFR_X1 \DRAM_mem_reg[20][9]  ( .D(n1518), .CK(CLK), .RN(n79), .Q(
        \DRAM_mem[20][9] ) );
  DFFR_X1 \DRAM_mem_reg[20][8]  ( .D(n1517), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[20][8] ) );
  DFFR_X1 \DRAM_mem_reg[20][7]  ( .D(n1516), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[20][7] ) );
  DFFR_X1 \DRAM_mem_reg[20][6]  ( .D(n1515), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[20][6] ) );
  DFFR_X1 \DRAM_mem_reg[20][5]  ( .D(n1514), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[20][5] ) );
  DFFR_X1 \DRAM_mem_reg[20][4]  ( .D(n1513), .CK(CLK), .RN(n71), .Q(
        \DRAM_mem[20][4] ) );
  DFFR_X1 \DRAM_mem_reg[20][3]  ( .D(n1512), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[20][3] ) );
  DFFR_X1 \DRAM_mem_reg[20][2]  ( .D(n1511), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[20][2] ) );
  DFFR_X1 \DRAM_mem_reg[20][1]  ( .D(n1510), .CK(CLK), .RN(n63), .Q(
        \DRAM_mem[20][1] ) );
  DFFR_X1 \DRAM_mem_reg[20][0]  ( .D(n1509), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[20][0] ) );
  DFFR_X1 \DRAM_mem_reg[21][31]  ( .D(n1508), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[21][31] ) );
  DFFR_X1 \DRAM_mem_reg[21][30]  ( .D(n1507), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[21][30] ) );
  DFFR_X1 \DRAM_mem_reg[21][29]  ( .D(n1506), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[21][29] ) );
  DFFR_X1 \DRAM_mem_reg[21][28]  ( .D(n1505), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[21][28] ) );
  DFFR_X1 \DRAM_mem_reg[21][27]  ( .D(n1504), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[21][27] ) );
  DFFR_X1 \DRAM_mem_reg[21][26]  ( .D(n1503), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[21][26] ) );
  DFFR_X1 \DRAM_mem_reg[21][25]  ( .D(n1502), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[21][25] ) );
  DFFR_X1 \DRAM_mem_reg[21][24]  ( .D(n1501), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[21][24] ) );
  DFFR_X1 \DRAM_mem_reg[21][23]  ( .D(n1500), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[21][23] ) );
  DFFR_X1 \DRAM_mem_reg[21][22]  ( .D(n1499), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[21][22] ) );
  DFFR_X1 \DRAM_mem_reg[21][21]  ( .D(n1498), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[21][21] ) );
  DFFR_X1 \DRAM_mem_reg[21][20]  ( .D(n1497), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[21][20] ) );
  DFFR_X1 \DRAM_mem_reg[21][19]  ( .D(n1496), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[21][19] ) );
  DFFR_X1 \DRAM_mem_reg[21][18]  ( .D(n1495), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[21][18] ) );
  DFFR_X1 \DRAM_mem_reg[21][17]  ( .D(n1494), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[21][17] ) );
  DFFR_X1 \DRAM_mem_reg[21][16]  ( .D(n1493), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[21][16] ) );
  DFFR_X1 \DRAM_mem_reg[21][15]  ( .D(n1492), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[21][15] ) );
  DFFR_X1 \DRAM_mem_reg[21][14]  ( .D(n1491), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[21][14] ) );
  DFFR_X1 \DRAM_mem_reg[21][13]  ( .D(n1490), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[21][13] ) );
  DFFR_X1 \DRAM_mem_reg[21][12]  ( .D(n1489), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[21][12] ) );
  DFFR_X1 \DRAM_mem_reg[21][11]  ( .D(n1488), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[21][11] ) );
  DFFR_X1 \DRAM_mem_reg[21][10]  ( .D(n1487), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[21][10] ) );
  DFFR_X1 \DRAM_mem_reg[21][9]  ( .D(n1486), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[21][9] ) );
  DFFR_X1 \DRAM_mem_reg[21][8]  ( .D(n1485), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[21][8] ) );
  DFFR_X1 \DRAM_mem_reg[21][7]  ( .D(n1484), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[21][7] ) );
  DFFR_X1 \DRAM_mem_reg[21][6]  ( .D(n1483), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[21][6] ) );
  DFFR_X1 \DRAM_mem_reg[21][5]  ( .D(n1482), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[21][5] ) );
  DFFR_X1 \DRAM_mem_reg[21][4]  ( .D(n1481), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[21][4] ) );
  DFFR_X1 \DRAM_mem_reg[21][3]  ( .D(n1480), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[21][3] ) );
  DFFR_X1 \DRAM_mem_reg[21][2]  ( .D(n1479), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[21][2] ) );
  DFFR_X1 \DRAM_mem_reg[21][1]  ( .D(n1478), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[21][1] ) );
  DFFR_X1 \DRAM_mem_reg[21][0]  ( .D(n1477), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[21][0] ) );
  DFFR_X1 \DRAM_mem_reg[22][31]  ( .D(n1476), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[22][31] ) );
  DFFR_X1 \DRAM_mem_reg[22][30]  ( .D(n1475), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[22][30] ) );
  DFFR_X1 \DRAM_mem_reg[22][29]  ( .D(n1474), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[22][29] ) );
  DFFR_X1 \DRAM_mem_reg[22][28]  ( .D(n1473), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[22][28] ) );
  DFFR_X1 \DRAM_mem_reg[22][27]  ( .D(n1472), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[22][27] ) );
  DFFR_X1 \DRAM_mem_reg[22][26]  ( .D(n1471), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[22][26] ) );
  DFFR_X1 \DRAM_mem_reg[22][25]  ( .D(n1470), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[22][25] ) );
  DFFR_X1 \DRAM_mem_reg[22][24]  ( .D(n1469), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[22][24] ) );
  DFFR_X1 \DRAM_mem_reg[22][23]  ( .D(n1468), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[22][23] ) );
  DFFR_X1 \DRAM_mem_reg[22][22]  ( .D(n1467), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[22][22] ) );
  DFFR_X1 \DRAM_mem_reg[22][21]  ( .D(n1466), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[22][21] ) );
  DFFR_X1 \DRAM_mem_reg[22][20]  ( .D(n1465), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[22][20] ) );
  DFFR_X1 \DRAM_mem_reg[22][19]  ( .D(n1464), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[22][19] ) );
  DFFR_X1 \DRAM_mem_reg[22][18]  ( .D(n1463), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[22][18] ) );
  DFFR_X1 \DRAM_mem_reg[22][17]  ( .D(n1462), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[22][17] ) );
  DFFR_X1 \DRAM_mem_reg[22][16]  ( .D(n1461), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[22][16] ) );
  DFFR_X1 \DRAM_mem_reg[22][15]  ( .D(n1460), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[22][15] ) );
  DFFR_X1 \DRAM_mem_reg[22][14]  ( .D(n1459), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[22][14] ) );
  DFFR_X1 \DRAM_mem_reg[22][13]  ( .D(n1458), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[22][13] ) );
  DFFR_X1 \DRAM_mem_reg[22][12]  ( .D(n1457), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[22][12] ) );
  DFFR_X1 \DRAM_mem_reg[22][11]  ( .D(n1456), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[22][11] ) );
  DFFR_X1 \DRAM_mem_reg[22][10]  ( .D(n1455), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[22][10] ) );
  DFFR_X1 \DRAM_mem_reg[22][9]  ( .D(n1454), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[22][9] ) );
  DFFR_X1 \DRAM_mem_reg[22][8]  ( .D(n1453), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[22][8] ) );
  DFFR_X1 \DRAM_mem_reg[22][7]  ( .D(n1452), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[22][7] ) );
  DFFR_X1 \DRAM_mem_reg[22][6]  ( .D(n1451), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[22][6] ) );
  DFFR_X1 \DRAM_mem_reg[22][5]  ( .D(n1450), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[22][5] ) );
  DFFR_X1 \DRAM_mem_reg[22][4]  ( .D(n1449), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[22][4] ) );
  DFFR_X1 \DRAM_mem_reg[22][3]  ( .D(n1448), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[22][3] ) );
  DFFR_X1 \DRAM_mem_reg[22][2]  ( .D(n1447), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[22][2] ) );
  DFFR_X1 \DRAM_mem_reg[22][1]  ( .D(n1446), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[22][1] ) );
  DFFR_X1 \DRAM_mem_reg[22][0]  ( .D(n1445), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[22][0] ) );
  DFFR_X1 \DRAM_mem_reg[23][31]  ( .D(n1444), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[23][31] ) );
  DFFR_X1 \DRAM_mem_reg[23][30]  ( .D(n1443), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[23][30] ) );
  DFFR_X1 \DRAM_mem_reg[23][29]  ( .D(n1442), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[23][29] ) );
  DFFR_X1 \DRAM_mem_reg[23][28]  ( .D(n1441), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[23][28] ) );
  DFFR_X1 \DRAM_mem_reg[23][27]  ( .D(n1440), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[23][27] ) );
  DFFR_X1 \DRAM_mem_reg[23][26]  ( .D(n1439), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[23][26] ) );
  DFFR_X1 \DRAM_mem_reg[23][25]  ( .D(n1438), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[23][25] ) );
  DFFR_X1 \DRAM_mem_reg[23][24]  ( .D(n1437), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[23][24] ) );
  DFFR_X1 \DRAM_mem_reg[23][23]  ( .D(n1436), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[23][23] ) );
  DFFR_X1 \DRAM_mem_reg[23][22]  ( .D(n1435), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[23][22] ) );
  DFFR_X1 \DRAM_mem_reg[23][21]  ( .D(n1434), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[23][21] ) );
  DFFR_X1 \DRAM_mem_reg[23][20]  ( .D(n1433), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[23][20] ) );
  DFFR_X1 \DRAM_mem_reg[23][19]  ( .D(n1432), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[23][19] ) );
  DFFR_X1 \DRAM_mem_reg[23][18]  ( .D(n1431), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[23][18] ) );
  DFFR_X1 \DRAM_mem_reg[23][17]  ( .D(n1430), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[23][17] ) );
  DFFR_X1 \DRAM_mem_reg[23][16]  ( .D(n1429), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[23][16] ) );
  DFFR_X1 \DRAM_mem_reg[23][15]  ( .D(n1428), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[23][15] ) );
  DFFR_X1 \DRAM_mem_reg[23][14]  ( .D(n1427), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[23][14] ) );
  DFFR_X1 \DRAM_mem_reg[23][13]  ( .D(n1426), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[23][13] ) );
  DFFR_X1 \DRAM_mem_reg[23][12]  ( .D(n1425), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[23][12] ) );
  DFFR_X1 \DRAM_mem_reg[23][11]  ( .D(n1424), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[23][11] ) );
  DFFR_X1 \DRAM_mem_reg[23][10]  ( .D(n1423), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[23][10] ) );
  DFFR_X1 \DRAM_mem_reg[23][9]  ( .D(n1422), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[23][9] ) );
  DFFR_X1 \DRAM_mem_reg[23][8]  ( .D(n1421), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[23][8] ) );
  DFFR_X1 \DRAM_mem_reg[23][7]  ( .D(n1420), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[23][7] ) );
  DFFR_X1 \DRAM_mem_reg[23][6]  ( .D(n1419), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[23][6] ) );
  DFFR_X1 \DRAM_mem_reg[23][5]  ( .D(n1418), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[23][5] ) );
  DFFR_X1 \DRAM_mem_reg[23][4]  ( .D(n1417), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[23][4] ) );
  DFFR_X1 \DRAM_mem_reg[23][3]  ( .D(n1416), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[23][3] ) );
  DFFR_X1 \DRAM_mem_reg[23][2]  ( .D(n1415), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[23][2] ) );
  DFFR_X1 \DRAM_mem_reg[23][1]  ( .D(n1414), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[23][1] ) );
  DFFR_X1 \DRAM_mem_reg[23][0]  ( .D(n1413), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[23][0] ) );
  DFFR_X1 \DRAM_mem_reg[24][31]  ( .D(n1412), .CK(CLK), .RN(n2), .Q(
        \DRAM_mem[24][31] ) );
  DFFR_X1 \DRAM_mem_reg[24][30]  ( .D(n1411), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[24][30] ) );
  DFFR_X1 \DRAM_mem_reg[24][29]  ( .D(n1410), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[24][29] ) );
  DFFR_X1 \DRAM_mem_reg[24][28]  ( .D(n1409), .CK(CLK), .RN(n10), .Q(
        \DRAM_mem[24][28] ) );
  DFFR_X1 \DRAM_mem_reg[24][27]  ( .D(n1408), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[24][27] ) );
  DFFR_X1 \DRAM_mem_reg[24][26]  ( .D(n1407), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[24][26] ) );
  DFFR_X1 \DRAM_mem_reg[24][25]  ( .D(n1406), .CK(CLK), .RN(n18), .Q(
        \DRAM_mem[24][25] ) );
  DFFR_X1 \DRAM_mem_reg[24][24]  ( .D(n1405), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[24][24] ) );
  DFFR_X1 \DRAM_mem_reg[24][23]  ( .D(n1404), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[24][23] ) );
  DFFR_X1 \DRAM_mem_reg[24][22]  ( .D(n1403), .CK(CLK), .RN(n26), .Q(
        \DRAM_mem[24][22] ) );
  DFFR_X1 \DRAM_mem_reg[24][21]  ( .D(n1402), .CK(CLK), .RN(n34), .Q(
        \DRAM_mem[24][21] ) );
  DFFR_X1 \DRAM_mem_reg[24][20]  ( .D(n1401), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[24][20] ) );
  DFFR_X1 \DRAM_mem_reg[24][19]  ( .D(n1400), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[24][19] ) );
  DFFR_X1 \DRAM_mem_reg[24][18]  ( .D(n1399), .CK(CLK), .RN(n42), .Q(
        \DRAM_mem[24][18] ) );
  DFFR_X1 \DRAM_mem_reg[24][17]  ( .D(n1398), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[24][17] ) );
  DFFR_X1 \DRAM_mem_reg[24][16]  ( .D(n1397), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[24][16] ) );
  DFFR_X1 \DRAM_mem_reg[24][15]  ( .D(n1396), .CK(CLK), .RN(n50), .Q(
        \DRAM_mem[24][15] ) );
  DFFR_X1 \DRAM_mem_reg[24][14]  ( .D(n1395), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[24][14] ) );
  DFFR_X1 \DRAM_mem_reg[24][13]  ( .D(n1394), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[24][13] ) );
  DFFR_X1 \DRAM_mem_reg[24][12]  ( .D(n1393), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[24][12] ) );
  DFFR_X1 \DRAM_mem_reg[24][11]  ( .D(n1392), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[24][11] ) );
  DFFR_X1 \DRAM_mem_reg[24][10]  ( .D(n1391), .CK(CLK), .RN(n58), .Q(
        \DRAM_mem[24][10] ) );
  DFFR_X1 \DRAM_mem_reg[24][9]  ( .D(n1390), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[24][9] ) );
  DFFR_X1 \DRAM_mem_reg[24][8]  ( .D(n1389), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[24][8] ) );
  DFFR_X1 \DRAM_mem_reg[24][7]  ( .D(n1388), .CK(CLK), .RN(n82), .Q(
        \DRAM_mem[24][7] ) );
  DFFR_X1 \DRAM_mem_reg[24][6]  ( .D(n1387), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[24][6] ) );
  DFFR_X1 \DRAM_mem_reg[24][5]  ( .D(n1386), .CK(CLK), .RN(n74), .Q(
        \DRAM_mem[24][5] ) );
  DFFR_X1 \DRAM_mem_reg[24][4]  ( .D(n1385), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[24][4] ) );
  DFFR_X1 \DRAM_mem_reg[24][3]  ( .D(n1384), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[24][3] ) );
  DFFR_X1 \DRAM_mem_reg[24][2]  ( .D(n1383), .CK(CLK), .RN(n66), .Q(
        \DRAM_mem[24][2] ) );
  DFFR_X1 \DRAM_mem_reg[24][1]  ( .D(n1382), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[24][1] ) );
  DFFR_X1 \DRAM_mem_reg[24][0]  ( .D(n1381), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[24][0] ) );
  DFFR_X1 \DRAM_mem_reg[25][31]  ( .D(n1380), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[25][31] ) );
  DFFR_X1 \DRAM_mem_reg[25][30]  ( .D(n1379), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[25][30] ) );
  DFFR_X1 \DRAM_mem_reg[25][29]  ( .D(n1378), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[25][29] ) );
  DFFR_X1 \DRAM_mem_reg[25][28]  ( .D(n1377), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[25][28] ) );
  DFFR_X1 \DRAM_mem_reg[25][27]  ( .D(n1376), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[25][27] ) );
  DFFR_X1 \DRAM_mem_reg[25][26]  ( .D(n1375), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[25][26] ) );
  DFFR_X1 \DRAM_mem_reg[25][25]  ( .D(n1374), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[25][25] ) );
  DFFR_X1 \DRAM_mem_reg[25][24]  ( .D(n1373), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[25][24] ) );
  DFFR_X1 \DRAM_mem_reg[25][23]  ( .D(n1372), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[25][23] ) );
  DFFR_X1 \DRAM_mem_reg[25][22]  ( .D(n1371), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[25][22] ) );
  DFFR_X1 \DRAM_mem_reg[25][21]  ( .D(n1370), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[25][21] ) );
  DFFR_X1 \DRAM_mem_reg[25][20]  ( .D(n1369), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[25][20] ) );
  DFFR_X1 \DRAM_mem_reg[25][19]  ( .D(n1368), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[25][19] ) );
  DFFR_X1 \DRAM_mem_reg[25][18]  ( .D(n1367), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[25][18] ) );
  DFFR_X1 \DRAM_mem_reg[25][17]  ( .D(n1366), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[25][17] ) );
  DFFR_X1 \DRAM_mem_reg[25][16]  ( .D(n1365), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[25][16] ) );
  DFFR_X1 \DRAM_mem_reg[25][15]  ( .D(n1364), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[25][15] ) );
  DFFR_X1 \DRAM_mem_reg[25][14]  ( .D(n1363), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[25][14] ) );
  DFFR_X1 \DRAM_mem_reg[25][13]  ( .D(n1362), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[25][13] ) );
  DFFR_X1 \DRAM_mem_reg[25][12]  ( .D(n1361), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[25][12] ) );
  DFFR_X1 \DRAM_mem_reg[25][11]  ( .D(n1360), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[25][11] ) );
  DFFR_X1 \DRAM_mem_reg[25][10]  ( .D(n1359), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[25][10] ) );
  DFFR_X1 \DRAM_mem_reg[25][9]  ( .D(n1358), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[25][9] ) );
  DFFR_X1 \DRAM_mem_reg[25][8]  ( .D(n1357), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[25][8] ) );
  DFFR_X1 \DRAM_mem_reg[25][7]  ( .D(n1356), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[25][7] ) );
  DFFR_X1 \DRAM_mem_reg[25][6]  ( .D(n1355), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[25][6] ) );
  DFFR_X1 \DRAM_mem_reg[25][5]  ( .D(n1354), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[25][5] ) );
  DFFR_X1 \DRAM_mem_reg[25][4]  ( .D(n1353), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[25][4] ) );
  DFFR_X1 \DRAM_mem_reg[25][3]  ( .D(n1352), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[25][3] ) );
  DFFR_X1 \DRAM_mem_reg[25][2]  ( .D(n1351), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[25][2] ) );
  DFFR_X1 \DRAM_mem_reg[25][1]  ( .D(n1350), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[25][1] ) );
  DFFR_X1 \DRAM_mem_reg[25][0]  ( .D(n1349), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[25][0] ) );
  DFFR_X1 \DRAM_mem_reg[26][31]  ( .D(n1348), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[26][31] ) );
  DFFR_X1 \DRAM_mem_reg[26][30]  ( .D(n1347), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[26][30] ) );
  DFFR_X1 \DRAM_mem_reg[26][29]  ( .D(n1346), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[26][29] ) );
  DFFR_X1 \DRAM_mem_reg[26][28]  ( .D(n1345), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[26][28] ) );
  DFFR_X1 \DRAM_mem_reg[26][27]  ( .D(n1344), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[26][27] ) );
  DFFR_X1 \DRAM_mem_reg[26][26]  ( .D(n1343), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[26][26] ) );
  DFFR_X1 \DRAM_mem_reg[26][25]  ( .D(n1342), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[26][25] ) );
  DFFR_X1 \DRAM_mem_reg[26][24]  ( .D(n1341), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[26][24] ) );
  DFFR_X1 \DRAM_mem_reg[26][23]  ( .D(n1340), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[26][23] ) );
  DFFR_X1 \DRAM_mem_reg[26][22]  ( .D(n1339), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[26][22] ) );
  DFFR_X1 \DRAM_mem_reg[26][21]  ( .D(n1338), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[26][21] ) );
  DFFR_X1 \DRAM_mem_reg[26][20]  ( .D(n1337), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[26][20] ) );
  DFFR_X1 \DRAM_mem_reg[26][19]  ( .D(n1336), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[26][19] ) );
  DFFR_X1 \DRAM_mem_reg[26][18]  ( .D(n1335), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[26][18] ) );
  DFFR_X1 \DRAM_mem_reg[26][17]  ( .D(n1334), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[26][17] ) );
  DFFR_X1 \DRAM_mem_reg[26][16]  ( .D(n1333), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[26][16] ) );
  DFFR_X1 \DRAM_mem_reg[26][15]  ( .D(n1332), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[26][15] ) );
  DFFR_X1 \DRAM_mem_reg[26][14]  ( .D(n1331), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[26][14] ) );
  DFFR_X1 \DRAM_mem_reg[26][13]  ( .D(n1330), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[26][13] ) );
  DFFR_X1 \DRAM_mem_reg[26][12]  ( .D(n1329), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[26][12] ) );
  DFFR_X1 \DRAM_mem_reg[26][11]  ( .D(n1328), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[26][11] ) );
  DFFR_X1 \DRAM_mem_reg[26][10]  ( .D(n1327), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[26][10] ) );
  DFFR_X1 \DRAM_mem_reg[26][9]  ( .D(n1326), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[26][9] ) );
  DFFR_X1 \DRAM_mem_reg[26][8]  ( .D(n1325), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[26][8] ) );
  DFFR_X1 \DRAM_mem_reg[26][7]  ( .D(n1324), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[26][7] ) );
  DFFR_X1 \DRAM_mem_reg[26][6]  ( .D(n1323), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[26][6] ) );
  DFFR_X1 \DRAM_mem_reg[26][5]  ( .D(n1322), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[26][5] ) );
  DFFR_X1 \DRAM_mem_reg[26][4]  ( .D(n1321), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[26][4] ) );
  DFFR_X1 \DRAM_mem_reg[26][3]  ( .D(n1320), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[26][3] ) );
  DFFR_X1 \DRAM_mem_reg[26][2]  ( .D(n1319), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[26][2] ) );
  DFFR_X1 \DRAM_mem_reg[26][1]  ( .D(n1318), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[26][1] ) );
  DFFR_X1 \DRAM_mem_reg[26][0]  ( .D(n1317), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[26][0] ) );
  DFFR_X1 \DRAM_mem_reg[27][31]  ( .D(n1316), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[27][31] ) );
  DFFR_X1 \DRAM_mem_reg[27][30]  ( .D(n1315), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[27][30] ) );
  DFFR_X1 \DRAM_mem_reg[27][29]  ( .D(n1314), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[27][29] ) );
  DFFR_X1 \DRAM_mem_reg[27][28]  ( .D(n1313), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[27][28] ) );
  DFFR_X1 \DRAM_mem_reg[27][27]  ( .D(n1312), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[27][27] ) );
  DFFR_X1 \DRAM_mem_reg[27][26]  ( .D(n1311), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[27][26] ) );
  DFFR_X1 \DRAM_mem_reg[27][25]  ( .D(n1310), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[27][25] ) );
  DFFR_X1 \DRAM_mem_reg[27][24]  ( .D(n1309), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[27][24] ) );
  DFFR_X1 \DRAM_mem_reg[27][23]  ( .D(n1308), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[27][23] ) );
  DFFR_X1 \DRAM_mem_reg[27][22]  ( .D(n1307), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[27][22] ) );
  DFFR_X1 \DRAM_mem_reg[27][21]  ( .D(n1306), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[27][21] ) );
  DFFR_X1 \DRAM_mem_reg[27][20]  ( .D(n1305), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[27][20] ) );
  DFFR_X1 \DRAM_mem_reg[27][19]  ( .D(n1304), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[27][19] ) );
  DFFR_X1 \DRAM_mem_reg[27][18]  ( .D(n1303), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[27][18] ) );
  DFFR_X1 \DRAM_mem_reg[27][17]  ( .D(n1302), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[27][17] ) );
  DFFR_X1 \DRAM_mem_reg[27][16]  ( .D(n1301), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[27][16] ) );
  DFFR_X1 \DRAM_mem_reg[27][15]  ( .D(n1300), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[27][15] ) );
  DFFR_X1 \DRAM_mem_reg[27][14]  ( .D(n1299), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[27][14] ) );
  DFFR_X1 \DRAM_mem_reg[27][13]  ( .D(n1298), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[27][13] ) );
  DFFR_X1 \DRAM_mem_reg[27][12]  ( .D(n1297), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[27][12] ) );
  DFFR_X1 \DRAM_mem_reg[27][11]  ( .D(n1296), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[27][11] ) );
  DFFR_X1 \DRAM_mem_reg[27][10]  ( .D(n1295), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[27][10] ) );
  DFFR_X1 \DRAM_mem_reg[27][9]  ( .D(n1294), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[27][9] ) );
  DFFR_X1 \DRAM_mem_reg[27][8]  ( .D(n1293), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[27][8] ) );
  DFFR_X1 \DRAM_mem_reg[27][7]  ( .D(n1292), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[27][7] ) );
  DFFR_X1 \DRAM_mem_reg[27][6]  ( .D(n1291), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[27][6] ) );
  DFFR_X1 \DRAM_mem_reg[27][5]  ( .D(n1290), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[27][5] ) );
  DFFR_X1 \DRAM_mem_reg[27][4]  ( .D(n1289), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[27][4] ) );
  DFFR_X1 \DRAM_mem_reg[27][3]  ( .D(n1288), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[27][3] ) );
  DFFR_X1 \DRAM_mem_reg[27][2]  ( .D(n1287), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[27][2] ) );
  DFFR_X1 \DRAM_mem_reg[27][1]  ( .D(n1286), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[27][1] ) );
  DFFR_X1 \DRAM_mem_reg[27][0]  ( .D(n1285), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[27][0] ) );
  DFFR_X1 \DRAM_mem_reg[28][31]  ( .D(n1284), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[28][31] ) );
  DFFR_X1 \DRAM_mem_reg[28][30]  ( .D(n1283), .CK(CLK), .RN(n5), .Q(
        \DRAM_mem[28][30] ) );
  DFFR_X1 \DRAM_mem_reg[28][29]  ( .D(n1282), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[28][29] ) );
  DFFR_X1 \DRAM_mem_reg[28][28]  ( .D(n1281), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[28][28] ) );
  DFFR_X1 \DRAM_mem_reg[28][27]  ( .D(n1280), .CK(CLK), .RN(n13), .Q(
        \DRAM_mem[28][27] ) );
  DFFR_X1 \DRAM_mem_reg[28][26]  ( .D(n1279), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[28][26] ) );
  DFFR_X1 \DRAM_mem_reg[28][25]  ( .D(n1278), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[28][25] ) );
  DFFR_X1 \DRAM_mem_reg[28][24]  ( .D(n1277), .CK(CLK), .RN(n21), .Q(
        \DRAM_mem[28][24] ) );
  DFFR_X1 \DRAM_mem_reg[28][23]  ( .D(n1276), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[28][23] ) );
  DFFR_X1 \DRAM_mem_reg[28][22]  ( .D(n1275), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[28][22] ) );
  DFFR_X1 \DRAM_mem_reg[28][21]  ( .D(n1274), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[28][21] ) );
  DFFR_X1 \DRAM_mem_reg[28][20]  ( .D(n1273), .CK(CLK), .RN(n37), .Q(
        \DRAM_mem[28][20] ) );
  DFFR_X1 \DRAM_mem_reg[28][19]  ( .D(n1272), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[28][19] ) );
  DFFR_X1 \DRAM_mem_reg[28][18]  ( .D(n1271), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[28][18] ) );
  DFFR_X1 \DRAM_mem_reg[28][17]  ( .D(n1270), .CK(CLK), .RN(n45), .Q(
        \DRAM_mem[28][17] ) );
  DFFR_X1 \DRAM_mem_reg[28][16]  ( .D(n1269), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[28][16] ) );
  DFFR_X1 \DRAM_mem_reg[28][15]  ( .D(n1268), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[28][15] ) );
  DFFR_X1 \DRAM_mem_reg[28][14]  ( .D(n1267), .CK(CLK), .RN(n53), .Q(
        \DRAM_mem[28][14] ) );
  DFFR_X1 \DRAM_mem_reg[28][13]  ( .D(n1266), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[28][13] ) );
  DFFR_X1 \DRAM_mem_reg[28][12]  ( .D(n1265), .CK(CLK), .RN(n29), .Q(
        \DRAM_mem[28][12] ) );
  DFFR_X1 \DRAM_mem_reg[28][11]  ( .D(n1264), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[28][11] ) );
  DFFR_X1 \DRAM_mem_reg[28][10]  ( .D(n1263), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[28][10] ) );
  DFFR_X1 \DRAM_mem_reg[28][9]  ( .D(n1262), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[28][9] ) );
  DFFR_X1 \DRAM_mem_reg[28][8]  ( .D(n1261), .CK(CLK), .RN(n85), .Q(
        \DRAM_mem[28][8] ) );
  DFFR_X1 \DRAM_mem_reg[28][7]  ( .D(n1260), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[28][7] ) );
  DFFR_X1 \DRAM_mem_reg[28][6]  ( .D(n1259), .CK(CLK), .RN(n77), .Q(
        \DRAM_mem[28][6] ) );
  DFFR_X1 \DRAM_mem_reg[28][5]  ( .D(n1258), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[28][5] ) );
  DFFR_X1 \DRAM_mem_reg[28][4]  ( .D(n1257), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[28][4] ) );
  DFFR_X1 \DRAM_mem_reg[28][3]  ( .D(n1256), .CK(CLK), .RN(n69), .Q(
        \DRAM_mem[28][3] ) );
  DFFR_X1 \DRAM_mem_reg[28][2]  ( .D(n1255), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[28][2] ) );
  DFFR_X1 \DRAM_mem_reg[28][1]  ( .D(n1254), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[28][1] ) );
  DFFR_X1 \DRAM_mem_reg[28][0]  ( .D(n1253), .CK(CLK), .RN(n61), .Q(
        \DRAM_mem[28][0] ) );
  DFFR_X1 \DRAM_mem_reg[29][31]  ( .D(n1252), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[29][31] ) );
  DFFR_X1 \DRAM_mem_reg[29][30]  ( .D(n1251), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[29][30] ) );
  DFFR_X1 \DRAM_mem_reg[29][29]  ( .D(n1250), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[29][29] ) );
  DFFR_X1 \DRAM_mem_reg[29][28]  ( .D(n1249), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[29][28] ) );
  DFFR_X1 \DRAM_mem_reg[29][27]  ( .D(n1248), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[29][27] ) );
  DFFR_X1 \DRAM_mem_reg[29][26]  ( .D(n1247), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[29][26] ) );
  DFFR_X1 \DRAM_mem_reg[29][25]  ( .D(n1246), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[29][25] ) );
  DFFR_X1 \DRAM_mem_reg[29][24]  ( .D(n1245), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[29][24] ) );
  DFFR_X1 \DRAM_mem_reg[29][23]  ( .D(n1244), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[29][23] ) );
  DFFR_X1 \DRAM_mem_reg[29][22]  ( .D(n1243), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[29][22] ) );
  DFFR_X1 \DRAM_mem_reg[29][21]  ( .D(n1242), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[29][21] ) );
  DFFR_X1 \DRAM_mem_reg[29][20]  ( .D(n1241), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[29][20] ) );
  DFFR_X1 \DRAM_mem_reg[29][19]  ( .D(n1240), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[29][19] ) );
  DFFR_X1 \DRAM_mem_reg[29][18]  ( .D(n1239), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[29][18] ) );
  DFFR_X1 \DRAM_mem_reg[29][17]  ( .D(n1238), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[29][17] ) );
  DFFR_X1 \DRAM_mem_reg[29][16]  ( .D(n1237), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[29][16] ) );
  DFFR_X1 \DRAM_mem_reg[29][15]  ( .D(n1236), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[29][15] ) );
  DFFR_X1 \DRAM_mem_reg[29][14]  ( .D(n1235), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[29][14] ) );
  DFFR_X1 \DRAM_mem_reg[29][13]  ( .D(n1234), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[29][13] ) );
  DFFR_X1 \DRAM_mem_reg[29][12]  ( .D(n1233), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[29][12] ) );
  DFFR_X1 \DRAM_mem_reg[29][11]  ( .D(n1232), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[29][11] ) );
  DFFR_X1 \DRAM_mem_reg[29][10]  ( .D(n1231), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[29][10] ) );
  DFFR_X1 \DRAM_mem_reg[29][9]  ( .D(n1230), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[29][9] ) );
  DFFR_X1 \DRAM_mem_reg[29][8]  ( .D(n1229), .CK(CLK), .RN(n86), .Q(
        \DRAM_mem[29][8] ) );
  DFFR_X1 \DRAM_mem_reg[29][7]  ( .D(n1228), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[29][7] ) );
  DFFR_X1 \DRAM_mem_reg[29][6]  ( .D(n1227), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[29][6] ) );
  DFFR_X1 \DRAM_mem_reg[29][5]  ( .D(n1226), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[29][5] ) );
  DFFR_X1 \DRAM_mem_reg[29][4]  ( .D(n1225), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[29][4] ) );
  DFFR_X1 \DRAM_mem_reg[29][3]  ( .D(n1224), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[29][3] ) );
  DFFR_X1 \DRAM_mem_reg[29][2]  ( .D(n1223), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[29][2] ) );
  DFFR_X1 \DRAM_mem_reg[29][1]  ( .D(n1222), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[29][1] ) );
  DFFR_X1 \DRAM_mem_reg[29][0]  ( .D(n1221), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[29][0] ) );
  DFFR_X1 \DRAM_mem_reg[30][31]  ( .D(n1220), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[30][31] ) );
  DFFR_X1 \DRAM_mem_reg[30][30]  ( .D(n1219), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[30][30] ) );
  DFFR_X1 \DRAM_mem_reg[30][29]  ( .D(n1218), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[30][29] ) );
  DFFR_X1 \DRAM_mem_reg[30][28]  ( .D(n1217), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[30][28] ) );
  DFFR_X1 \DRAM_mem_reg[30][27]  ( .D(n1216), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[30][27] ) );
  DFFR_X1 \DRAM_mem_reg[30][26]  ( .D(n1215), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[30][26] ) );
  DFFR_X1 \DRAM_mem_reg[30][25]  ( .D(n1214), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[30][25] ) );
  DFFR_X1 \DRAM_mem_reg[30][24]  ( .D(n1213), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[30][24] ) );
  DFFR_X1 \DRAM_mem_reg[30][23]  ( .D(n1212), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[30][23] ) );
  DFFR_X1 \DRAM_mem_reg[30][22]  ( .D(n1211), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[30][22] ) );
  DFFR_X1 \DRAM_mem_reg[30][21]  ( .D(n1210), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[30][21] ) );
  DFFR_X1 \DRAM_mem_reg[30][20]  ( .D(n1209), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[30][20] ) );
  DFFR_X1 \DRAM_mem_reg[30][19]  ( .D(n1208), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[30][19] ) );
  DFFR_X1 \DRAM_mem_reg[30][18]  ( .D(n1207), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[30][18] ) );
  DFFR_X1 \DRAM_mem_reg[30][17]  ( .D(n1206), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[30][17] ) );
  DFFR_X1 \DRAM_mem_reg[30][16]  ( .D(n1205), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[30][16] ) );
  DFFR_X1 \DRAM_mem_reg[30][15]  ( .D(n1204), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[30][15] ) );
  DFFR_X1 \DRAM_mem_reg[30][14]  ( .D(n1203), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[30][14] ) );
  DFFR_X1 \DRAM_mem_reg[30][13]  ( .D(n1202), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[30][13] ) );
  DFFR_X1 \DRAM_mem_reg[30][12]  ( .D(n1201), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[30][12] ) );
  DFFR_X1 \DRAM_mem_reg[30][11]  ( .D(n1200), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[30][11] ) );
  DFFR_X1 \DRAM_mem_reg[30][10]  ( .D(n1199), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[30][10] ) );
  DFFR_X1 \DRAM_mem_reg[30][9]  ( .D(n1198), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[30][9] ) );
  DFFR_X1 \DRAM_mem_reg[30][8]  ( .D(n1197), .CK(CLK), .RN(n86), .Q(
        \DRAM_mem[30][8] ) );
  DFFR_X1 \DRAM_mem_reg[30][7]  ( .D(n1196), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[30][7] ) );
  DFFR_X1 \DRAM_mem_reg[30][6]  ( .D(n1195), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[30][6] ) );
  DFFR_X1 \DRAM_mem_reg[30][5]  ( .D(n1194), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[30][5] ) );
  DFFR_X1 \DRAM_mem_reg[30][4]  ( .D(n1193), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[30][4] ) );
  DFFR_X1 \DRAM_mem_reg[30][3]  ( .D(n1192), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[30][3] ) );
  DFFR_X1 \DRAM_mem_reg[30][2]  ( .D(n1191), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[30][2] ) );
  DFFR_X1 \DRAM_mem_reg[30][1]  ( .D(n1190), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[30][1] ) );
  DFFR_X1 \DRAM_mem_reg[30][0]  ( .D(n1189), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[30][0] ) );
  DFFR_X1 \DRAM_mem_reg[31][31]  ( .D(n1188), .CK(CLK), .RN(n3), .Q(
        \DRAM_mem[31][31] ) );
  DFFR_X1 \DRAM_mem_reg[31][30]  ( .D(n1187), .CK(CLK), .RN(n6), .Q(
        \DRAM_mem[31][30] ) );
  DFFR_X1 \DRAM_mem_reg[31][29]  ( .D(n1186), .CK(CLK), .RN(n8), .Q(
        \DRAM_mem[31][29] ) );
  DFFR_X1 \DRAM_mem_reg[31][28]  ( .D(n1185), .CK(CLK), .RN(n11), .Q(
        \DRAM_mem[31][28] ) );
  DFFR_X1 \DRAM_mem_reg[31][27]  ( .D(n1184), .CK(CLK), .RN(n14), .Q(
        \DRAM_mem[31][27] ) );
  DFFR_X1 \DRAM_mem_reg[31][26]  ( .D(n1183), .CK(CLK), .RN(n16), .Q(
        \DRAM_mem[31][26] ) );
  DFFR_X1 \DRAM_mem_reg[31][25]  ( .D(n1182), .CK(CLK), .RN(n19), .Q(
        \DRAM_mem[31][25] ) );
  DFFR_X1 \DRAM_mem_reg[31][24]  ( .D(n1181), .CK(CLK), .RN(n22), .Q(
        \DRAM_mem[31][24] ) );
  DFFR_X1 \DRAM_mem_reg[31][23]  ( .D(n1180), .CK(CLK), .RN(n24), .Q(
        \DRAM_mem[31][23] ) );
  DFFR_X1 \DRAM_mem_reg[31][22]  ( .D(n1179), .CK(CLK), .RN(n27), .Q(
        \DRAM_mem[31][22] ) );
  DFFR_X1 \DRAM_mem_reg[31][21]  ( .D(n1178), .CK(CLK), .RN(n35), .Q(
        \DRAM_mem[31][21] ) );
  DFFR_X1 \DRAM_mem_reg[31][20]  ( .D(n1177), .CK(CLK), .RN(n38), .Q(
        \DRAM_mem[31][20] ) );
  DFFR_X1 \DRAM_mem_reg[31][19]  ( .D(n1176), .CK(CLK), .RN(n40), .Q(
        \DRAM_mem[31][19] ) );
  DFFR_X1 \DRAM_mem_reg[31][18]  ( .D(n1175), .CK(CLK), .RN(n43), .Q(
        \DRAM_mem[31][18] ) );
  DFFR_X1 \DRAM_mem_reg[31][17]  ( .D(n1174), .CK(CLK), .RN(n46), .Q(
        \DRAM_mem[31][17] ) );
  DFFR_X1 \DRAM_mem_reg[31][16]  ( .D(n1173), .CK(CLK), .RN(n48), .Q(
        \DRAM_mem[31][16] ) );
  DFFR_X1 \DRAM_mem_reg[31][15]  ( .D(n1172), .CK(CLK), .RN(n51), .Q(
        \DRAM_mem[31][15] ) );
  DFFR_X1 \DRAM_mem_reg[31][14]  ( .D(n1171), .CK(CLK), .RN(n54), .Q(
        \DRAM_mem[31][14] ) );
  DFFR_X1 \DRAM_mem_reg[31][13]  ( .D(n1170), .CK(CLK), .RN(n32), .Q(
        \DRAM_mem[31][13] ) );
  DFFR_X1 \DRAM_mem_reg[31][12]  ( .D(n1169), .CK(CLK), .RN(n30), .Q(
        \DRAM_mem[31][12] ) );
  DFFR_X1 \DRAM_mem_reg[31][11]  ( .D(n1168), .CK(CLK), .RN(n56), .Q(
        \DRAM_mem[31][11] ) );
  DFFR_X1 \DRAM_mem_reg[31][10]  ( .D(n1167), .CK(CLK), .RN(n59), .Q(
        \DRAM_mem[31][10] ) );
  DFFR_X1 \DRAM_mem_reg[31][9]  ( .D(n1166), .CK(CLK), .RN(n80), .Q(
        \DRAM_mem[31][9] ) );
  DFFR_X1 \DRAM_mem_reg[31][8]  ( .D(n1165), .CK(CLK), .RN(n86), .Q(
        \DRAM_mem[31][8] ) );
  DFFR_X1 \DRAM_mem_reg[31][7]  ( .D(n1164), .CK(CLK), .RN(n83), .Q(
        \DRAM_mem[31][7] ) );
  DFFR_X1 \DRAM_mem_reg[31][6]  ( .D(n1163), .CK(CLK), .RN(n78), .Q(
        \DRAM_mem[31][6] ) );
  DFFR_X1 \DRAM_mem_reg[31][5]  ( .D(n1162), .CK(CLK), .RN(n75), .Q(
        \DRAM_mem[31][5] ) );
  DFFR_X1 \DRAM_mem_reg[31][4]  ( .D(n1161), .CK(CLK), .RN(n72), .Q(
        \DRAM_mem[31][4] ) );
  DFFR_X1 \DRAM_mem_reg[31][3]  ( .D(n1160), .CK(CLK), .RN(n70), .Q(
        \DRAM_mem[31][3] ) );
  DFFR_X1 \DRAM_mem_reg[31][2]  ( .D(n1159), .CK(CLK), .RN(n67), .Q(
        \DRAM_mem[31][2] ) );
  DFFR_X1 \DRAM_mem_reg[31][1]  ( .D(n1158), .CK(CLK), .RN(n64), .Q(
        \DRAM_mem[31][1] ) );
  DFFR_X1 \DRAM_mem_reg[31][0]  ( .D(n1157), .CK(CLK), .RN(n62), .Q(
        \DRAM_mem[31][0] ) );
  DLH_X1 \Dout_reg[31]  ( .G(N598), .D(N597), .Q(Dout[31]) );
  DLH_X1 \Dout_reg[30]  ( .G(N598), .D(N596), .Q(Dout[30]) );
  DLH_X1 \Dout_reg[29]  ( .G(N598), .D(N595), .Q(Dout[29]) );
  DLH_X1 \Dout_reg[28]  ( .G(N598), .D(N594), .Q(Dout[28]) );
  DLH_X1 \Dout_reg[27]  ( .G(N598), .D(N593), .Q(Dout[27]) );
  DLH_X1 \Dout_reg[26]  ( .G(N598), .D(N592), .Q(Dout[26]) );
  DLH_X1 \Dout_reg[25]  ( .G(N598), .D(N591), .Q(Dout[25]) );
  DLH_X1 \Dout_reg[24]  ( .G(N598), .D(N590), .Q(Dout[24]) );
  DLH_X1 \Dout_reg[23]  ( .G(N598), .D(N589), .Q(Dout[23]) );
  DLH_X1 \Dout_reg[22]  ( .G(N598), .D(N588), .Q(Dout[22]) );
  DLH_X1 \Dout_reg[21]  ( .G(N598), .D(N587), .Q(Dout[21]) );
  DLH_X1 \Dout_reg[20]  ( .G(N598), .D(N586), .Q(Dout[20]) );
  DLH_X1 \Dout_reg[19]  ( .G(N598), .D(N585), .Q(Dout[19]) );
  DLH_X1 \Dout_reg[18]  ( .G(N598), .D(N584), .Q(Dout[18]) );
  DLH_X1 \Dout_reg[17]  ( .G(N598), .D(N583), .Q(Dout[17]) );
  DLH_X1 \Dout_reg[16]  ( .G(N598), .D(N582), .Q(Dout[16]) );
  DLH_X1 \Dout_reg[15]  ( .G(N598), .D(N581), .Q(Dout[15]) );
  DLH_X1 \Dout_reg[14]  ( .G(N598), .D(N580), .Q(Dout[14]) );
  DLH_X1 \Dout_reg[13]  ( .G(N598), .D(N579), .Q(Dout[13]) );
  DLH_X1 \Dout_reg[12]  ( .G(N598), .D(N578), .Q(Dout[12]) );
  DLH_X1 \Dout_reg[11]  ( .G(N598), .D(N577), .Q(Dout[11]) );
  DLH_X1 \Dout_reg[10]  ( .G(N598), .D(N576), .Q(Dout[10]) );
  DLH_X1 \Dout_reg[9]  ( .G(N598), .D(N575), .Q(Dout[9]) );
  DLH_X1 \Dout_reg[8]  ( .G(N598), .D(N574), .Q(Dout[8]) );
  DLH_X1 \Dout_reg[7]  ( .G(N598), .D(N573), .Q(Dout[7]) );
  DLH_X1 \Dout_reg[6]  ( .G(N598), .D(N572), .Q(Dout[6]) );
  DLH_X1 \Dout_reg[5]  ( .G(N598), .D(N571), .Q(Dout[5]) );
  DLH_X1 \Dout_reg[4]  ( .G(N598), .D(N570), .Q(Dout[4]) );
  DLH_X1 \Dout_reg[3]  ( .G(N598), .D(N569), .Q(Dout[3]) );
  DLH_X1 \Dout_reg[2]  ( .G(N598), .D(N568), .Q(Dout[2]) );
  DLH_X1 \Dout_reg[1]  ( .G(N598), .D(N567), .Q(Dout[1]) );
  DLH_X1 \Dout_reg[0]  ( .G(N598), .D(N566), .Q(Dout[0]) );
  AND2_X2 U2 ( .A1(n2203), .A2(n2197), .ZN(n2202) );
  AND2_X2 U3 ( .A1(n2214), .A2(n2201), .ZN(n2216) );
  AND2_X2 U4 ( .A1(n2223), .A2(n2199), .ZN(n2224) );
  AND2_X2 U5 ( .A1(n2232), .A2(n2196), .ZN(n2231) );
  AND2_X2 U6 ( .A1(n2201), .A2(n2197), .ZN(n2200) );
  AND2_X2 U7 ( .A1(n2214), .A2(n2203), .ZN(n2217) );
  AND2_X2 U8 ( .A1(n2223), .A2(n2196), .ZN(n2222) );
  AND2_X2 U9 ( .A1(n2232), .A2(n2199), .ZN(n2233) );
  AND2_X2 U10 ( .A1(n2199), .A2(n2197), .ZN(n2198) );
  AND2_X2 U11 ( .A1(n2214), .A2(n2196), .ZN(n2213) );
  AND2_X2 U12 ( .A1(n2223), .A2(n2203), .ZN(n2226) );
  AND2_X2 U13 ( .A1(n2232), .A2(n2201), .ZN(n2235) );
  AND2_X2 U14 ( .A1(n2196), .A2(n2197), .ZN(n1140) );
  AND2_X2 U15 ( .A1(n2214), .A2(n2199), .ZN(n2215) );
  AND2_X2 U16 ( .A1(n2223), .A2(n2201), .ZN(n2225) );
  AND2_X2 U17 ( .A1(n2232), .A2(n2203), .ZN(n2237) );
  AND2_X2 U18 ( .A1(n2211), .A2(n2197), .ZN(n2210) );
  AND2_X2 U19 ( .A1(n2214), .A2(n2209), .ZN(n2220) );
  AND2_X2 U20 ( .A1(n2223), .A2(n2207), .ZN(n2228) );
  AND2_X2 U21 ( .A1(n2232), .A2(n2205), .ZN(n2238) );
  AND2_X2 U22 ( .A1(n2209), .A2(n2197), .ZN(n2208) );
  AND2_X2 U23 ( .A1(n2214), .A2(n2211), .ZN(n2221) );
  AND2_X2 U24 ( .A1(n2223), .A2(n2205), .ZN(n2227) );
  AND2_X2 U25 ( .A1(n2232), .A2(n2207), .ZN(n2239) );
  AND2_X2 U26 ( .A1(n2207), .A2(n2197), .ZN(n2206) );
  AND2_X2 U27 ( .A1(n2214), .A2(n2205), .ZN(n2218) );
  AND2_X2 U28 ( .A1(n2223), .A2(n2211), .ZN(n2230) );
  AND2_X2 U29 ( .A1(n2232), .A2(n2209), .ZN(n2240) );
  AOI21_X2 U30 ( .B1(n2263), .B2(N484), .A(n2295), .ZN(n2279) );
  AND2_X2 U31 ( .A1(n2205), .A2(n2197), .ZN(n2204) );
  AND2_X2 U32 ( .A1(n2214), .A2(n2207), .ZN(n2219) );
  AND2_X2 U33 ( .A1(n2223), .A2(n2209), .ZN(n2229) );
  AND2_X2 U34 ( .A1(n2232), .A2(n2211), .ZN(n2241) );
  BUF_X1 U35 ( .A(n178), .Z(n173) );
  BUF_X1 U36 ( .A(n178), .Z(n172) );
  BUF_X1 U37 ( .A(n178), .Z(n174) );
  BUF_X1 U38 ( .A(n178), .Z(n171) );
  BUF_X1 U39 ( .A(n178), .Z(n176) );
  BUF_X1 U40 ( .A(n178), .Z(n175) );
  BUF_X1 U41 ( .A(n2309), .Z(n91) );
  BUF_X1 U42 ( .A(n2309), .Z(n90) );
  BUF_X1 U43 ( .A(n2309), .Z(n89) );
  BUF_X1 U44 ( .A(n2309), .Z(n87) );
  BUF_X1 U45 ( .A(n2309), .Z(n88) );
  BUF_X1 U46 ( .A(n2309), .Z(n92) );
  BUF_X1 U47 ( .A(n2309), .Z(n93) );
  BUF_X1 U48 ( .A(n2309), .Z(n94) );
  BUF_X1 U49 ( .A(n2309), .Z(n95) );
  BUF_X1 U50 ( .A(n2309), .Z(n96) );
  BUF_X1 U51 ( .A(n2309), .Z(n97) );
  BUF_X1 U52 ( .A(n2309), .Z(n98) );
  BUF_X1 U53 ( .A(n2309), .Z(n99) );
  BUF_X1 U54 ( .A(n2309), .Z(n100) );
  BUF_X1 U55 ( .A(n2309), .Z(n101) );
  BUF_X1 U56 ( .A(n178), .Z(n177) );
  INV_X1 U57 ( .A(Addr[3]), .ZN(n132) );
  INV_X1 U58 ( .A(Addr[4]), .ZN(n178) );
  CLKBUF_X1 U59 ( .A(n101), .Z(n1) );
  CLKBUF_X1 U60 ( .A(n101), .Z(n2) );
  CLKBUF_X1 U61 ( .A(n100), .Z(n3) );
  CLKBUF_X1 U62 ( .A(n100), .Z(n4) );
  CLKBUF_X1 U63 ( .A(n100), .Z(n5) );
  CLKBUF_X1 U64 ( .A(n100), .Z(n6) );
  CLKBUF_X1 U65 ( .A(n100), .Z(n7) );
  CLKBUF_X1 U66 ( .A(n100), .Z(n8) );
  CLKBUF_X1 U67 ( .A(n99), .Z(n9) );
  CLKBUF_X1 U68 ( .A(n99), .Z(n10) );
  CLKBUF_X1 U69 ( .A(n99), .Z(n11) );
  CLKBUF_X1 U70 ( .A(n99), .Z(n12) );
  CLKBUF_X1 U71 ( .A(n99), .Z(n13) );
  CLKBUF_X1 U72 ( .A(n99), .Z(n14) );
  CLKBUF_X1 U73 ( .A(n98), .Z(n15) );
  CLKBUF_X1 U74 ( .A(n98), .Z(n16) );
  CLKBUF_X1 U75 ( .A(n98), .Z(n17) );
  CLKBUF_X1 U76 ( .A(n98), .Z(n18) );
  CLKBUF_X1 U77 ( .A(n98), .Z(n19) );
  CLKBUF_X1 U78 ( .A(n98), .Z(n20) );
  CLKBUF_X1 U79 ( .A(n97), .Z(n21) );
  CLKBUF_X1 U80 ( .A(n97), .Z(n22) );
  CLKBUF_X1 U81 ( .A(n97), .Z(n23) );
  CLKBUF_X1 U82 ( .A(n97), .Z(n24) );
  CLKBUF_X1 U83 ( .A(n97), .Z(n25) );
  CLKBUF_X1 U84 ( .A(n97), .Z(n26) );
  CLKBUF_X1 U85 ( .A(n96), .Z(n27) );
  CLKBUF_X1 U86 ( .A(n96), .Z(n28) );
  CLKBUF_X1 U87 ( .A(n96), .Z(n29) );
  CLKBUF_X1 U88 ( .A(n96), .Z(n30) );
  CLKBUF_X1 U89 ( .A(n96), .Z(n31) );
  CLKBUF_X1 U90 ( .A(n96), .Z(n32) );
  CLKBUF_X1 U91 ( .A(n95), .Z(n33) );
  CLKBUF_X1 U92 ( .A(n95), .Z(n34) );
  CLKBUF_X1 U93 ( .A(n95), .Z(n35) );
  CLKBUF_X1 U94 ( .A(n95), .Z(n36) );
  CLKBUF_X1 U95 ( .A(n95), .Z(n37) );
  CLKBUF_X1 U96 ( .A(n95), .Z(n38) );
  CLKBUF_X1 U97 ( .A(n94), .Z(n39) );
  CLKBUF_X1 U98 ( .A(n94), .Z(n40) );
  CLKBUF_X1 U99 ( .A(n94), .Z(n41) );
  CLKBUF_X1 U100 ( .A(n94), .Z(n42) );
  CLKBUF_X1 U101 ( .A(n94), .Z(n43) );
  CLKBUF_X1 U102 ( .A(n94), .Z(n44) );
  CLKBUF_X1 U103 ( .A(n93), .Z(n45) );
  CLKBUF_X1 U104 ( .A(n93), .Z(n46) );
  CLKBUF_X1 U105 ( .A(n93), .Z(n47) );
  CLKBUF_X1 U106 ( .A(n93), .Z(n48) );
  CLKBUF_X1 U107 ( .A(n93), .Z(n49) );
  CLKBUF_X1 U108 ( .A(n93), .Z(n50) );
  CLKBUF_X1 U109 ( .A(n92), .Z(n51) );
  CLKBUF_X1 U110 ( .A(n92), .Z(n52) );
  CLKBUF_X1 U111 ( .A(n92), .Z(n53) );
  CLKBUF_X1 U112 ( .A(n92), .Z(n54) );
  CLKBUF_X1 U113 ( .A(n92), .Z(n55) );
  CLKBUF_X1 U114 ( .A(n92), .Z(n56) );
  CLKBUF_X1 U115 ( .A(n91), .Z(n57) );
  CLKBUF_X1 U116 ( .A(n91), .Z(n58) );
  CLKBUF_X1 U117 ( .A(n91), .Z(n59) );
  CLKBUF_X1 U118 ( .A(n91), .Z(n60) );
  CLKBUF_X1 U119 ( .A(n91), .Z(n61) );
  CLKBUF_X1 U120 ( .A(n91), .Z(n62) );
  CLKBUF_X1 U121 ( .A(n90), .Z(n63) );
  CLKBUF_X1 U122 ( .A(n90), .Z(n64) );
  CLKBUF_X1 U123 ( .A(n90), .Z(n65) );
  CLKBUF_X1 U124 ( .A(n90), .Z(n66) );
  CLKBUF_X1 U125 ( .A(n90), .Z(n67) );
  CLKBUF_X1 U126 ( .A(n90), .Z(n68) );
  CLKBUF_X1 U127 ( .A(n89), .Z(n69) );
  CLKBUF_X1 U128 ( .A(n89), .Z(n70) );
  CLKBUF_X1 U129 ( .A(n89), .Z(n71) );
  CLKBUF_X1 U130 ( .A(n89), .Z(n72) );
  CLKBUF_X1 U131 ( .A(n89), .Z(n73) );
  CLKBUF_X1 U132 ( .A(n89), .Z(n74) );
  CLKBUF_X1 U133 ( .A(n88), .Z(n75) );
  CLKBUF_X1 U134 ( .A(n88), .Z(n76) );
  CLKBUF_X1 U135 ( .A(n88), .Z(n77) );
  CLKBUF_X1 U136 ( .A(n88), .Z(n78) );
  CLKBUF_X1 U137 ( .A(n88), .Z(n79) );
  CLKBUF_X1 U138 ( .A(n88), .Z(n80) );
  CLKBUF_X1 U139 ( .A(n87), .Z(n81) );
  CLKBUF_X1 U140 ( .A(n87), .Z(n82) );
  CLKBUF_X1 U141 ( .A(n87), .Z(n83) );
  CLKBUF_X1 U142 ( .A(n87), .Z(n84) );
  CLKBUF_X1 U143 ( .A(n87), .Z(n85) );
  CLKBUF_X1 U144 ( .A(n87), .Z(n86) );
  CLKBUF_X1 U145 ( .A(Addr[2]), .Z(n102) );
  CLKBUF_X1 U146 ( .A(Addr[2]), .Z(n103) );
  CLKBUF_X1 U147 ( .A(Addr[2]), .Z(n104) );
  CLKBUF_X1 U148 ( .A(Addr[2]), .Z(n105) );
  CLKBUF_X1 U149 ( .A(Addr[2]), .Z(n106) );
  CLKBUF_X1 U150 ( .A(Addr[2]), .Z(n107) );
  CLKBUF_X1 U151 ( .A(Addr[2]), .Z(n108) );
  CLKBUF_X1 U152 ( .A(Addr[2]), .Z(n109) );
  CLKBUF_X1 U153 ( .A(Addr[2]), .Z(n110) );
  CLKBUF_X1 U154 ( .A(Addr[2]), .Z(n111) );
  CLKBUF_X1 U155 ( .A(Addr[2]), .Z(n112) );
  CLKBUF_X1 U156 ( .A(Addr[2]), .Z(n113) );
  INV_X1 U157 ( .A(n132), .ZN(n114) );
  INV_X1 U158 ( .A(n132), .ZN(n115) );
  INV_X1 U159 ( .A(n132), .ZN(n116) );
  INV_X1 U160 ( .A(n132), .ZN(n117) );
  INV_X1 U161 ( .A(n132), .ZN(n118) );
  INV_X1 U162 ( .A(n132), .ZN(n119) );
  INV_X1 U163 ( .A(n132), .ZN(n120) );
  INV_X1 U164 ( .A(n132), .ZN(n121) );
  INV_X1 U165 ( .A(n132), .ZN(n122) );
  INV_X1 U166 ( .A(n132), .ZN(n123) );
  INV_X1 U167 ( .A(n132), .ZN(n124) );
  INV_X1 U168 ( .A(n132), .ZN(n125) );
  INV_X1 U169 ( .A(n132), .ZN(n126) );
  INV_X1 U170 ( .A(n132), .ZN(n127) );
  INV_X1 U171 ( .A(n132), .ZN(n128) );
  INV_X1 U172 ( .A(n132), .ZN(n129) );
  INV_X1 U173 ( .A(n132), .ZN(n130) );
  INV_X1 U174 ( .A(n132), .ZN(n131) );
  INV_X1 U175 ( .A(n176), .ZN(n133) );
  INV_X1 U176 ( .A(n176), .ZN(n134) );
  INV_X1 U177 ( .A(n176), .ZN(n135) );
  INV_X1 U178 ( .A(n176), .ZN(n136) );
  INV_X1 U179 ( .A(n176), .ZN(n137) );
  INV_X1 U180 ( .A(n176), .ZN(n138) );
  INV_X1 U181 ( .A(n176), .ZN(n139) );
  INV_X1 U182 ( .A(n175), .ZN(n140) );
  INV_X1 U183 ( .A(n175), .ZN(n141) );
  INV_X1 U184 ( .A(n175), .ZN(n142) );
  INV_X1 U185 ( .A(n175), .ZN(n143) );
  INV_X1 U186 ( .A(n175), .ZN(n144) );
  INV_X1 U187 ( .A(n175), .ZN(n145) );
  INV_X1 U188 ( .A(n175), .ZN(n146) );
  INV_X1 U189 ( .A(n174), .ZN(n147) );
  INV_X1 U190 ( .A(n174), .ZN(n148) );
  INV_X1 U191 ( .A(n174), .ZN(n149) );
  INV_X1 U192 ( .A(n174), .ZN(n150) );
  INV_X1 U193 ( .A(n174), .ZN(n151) );
  INV_X1 U194 ( .A(n174), .ZN(n152) );
  INV_X1 U195 ( .A(n174), .ZN(n153) );
  INV_X1 U196 ( .A(n173), .ZN(n154) );
  INV_X1 U197 ( .A(n173), .ZN(n155) );
  INV_X1 U198 ( .A(n173), .ZN(n156) );
  INV_X1 U199 ( .A(n173), .ZN(n157) );
  INV_X1 U200 ( .A(n173), .ZN(n158) );
  INV_X1 U201 ( .A(n173), .ZN(n159) );
  INV_X1 U202 ( .A(n173), .ZN(n160) );
  INV_X1 U203 ( .A(n172), .ZN(n161) );
  INV_X1 U204 ( .A(n172), .ZN(n162) );
  INV_X1 U205 ( .A(n172), .ZN(n163) );
  INV_X1 U206 ( .A(n172), .ZN(n164) );
  INV_X1 U207 ( .A(n172), .ZN(n165) );
  INV_X1 U208 ( .A(n172), .ZN(n166) );
  INV_X1 U209 ( .A(n172), .ZN(n167) );
  INV_X1 U210 ( .A(n171), .ZN(n168) );
  INV_X1 U211 ( .A(n171), .ZN(n169) );
  INV_X1 U212 ( .A(n171), .ZN(n170) );
  MUX2_X1 U213 ( .A(\DRAM_mem[15][0] ), .B(\DRAM_mem[31][0] ), .S(Addr[4]), 
        .Z(n179) );
  MUX2_X1 U214 ( .A(\DRAM_mem[7][0] ), .B(\DRAM_mem[23][0] ), .S(n154), .Z(
        n180) );
  MUX2_X1 U215 ( .A(n180), .B(n179), .S(n114), .Z(n181) );
  MUX2_X1 U216 ( .A(\DRAM_mem[11][0] ), .B(\DRAM_mem[27][0] ), .S(Addr[4]), 
        .Z(n182) );
  MUX2_X1 U217 ( .A(\DRAM_mem[3][0] ), .B(\DRAM_mem[19][0] ), .S(Addr[4]), .Z(
        n183) );
  MUX2_X1 U218 ( .A(n183), .B(n182), .S(n114), .Z(n184) );
  MUX2_X1 U219 ( .A(n184), .B(n181), .S(n102), .Z(n185) );
  MUX2_X1 U220 ( .A(\DRAM_mem[14][0] ), .B(\DRAM_mem[30][0] ), .S(Addr[4]), 
        .Z(n186) );
  MUX2_X1 U221 ( .A(\DRAM_mem[6][0] ), .B(\DRAM_mem[22][0] ), .S(Addr[4]), .Z(
        n187) );
  MUX2_X1 U222 ( .A(n187), .B(n186), .S(n114), .Z(n188) );
  MUX2_X1 U223 ( .A(\DRAM_mem[10][0] ), .B(\DRAM_mem[26][0] ), .S(Addr[4]), 
        .Z(n189) );
  MUX2_X1 U224 ( .A(\DRAM_mem[2][0] ), .B(\DRAM_mem[18][0] ), .S(Addr[4]), .Z(
        n190) );
  MUX2_X1 U225 ( .A(n190), .B(n189), .S(n114), .Z(n191) );
  MUX2_X1 U226 ( .A(n191), .B(n188), .S(n102), .Z(n192) );
  MUX2_X1 U227 ( .A(n192), .B(n185), .S(Addr[0]), .Z(n193) );
  MUX2_X1 U228 ( .A(\DRAM_mem[13][0] ), .B(\DRAM_mem[29][0] ), .S(Addr[4]), 
        .Z(n194) );
  MUX2_X1 U229 ( .A(\DRAM_mem[5][0] ), .B(\DRAM_mem[21][0] ), .S(Addr[4]), .Z(
        n195) );
  MUX2_X1 U230 ( .A(n195), .B(n194), .S(n114), .Z(n196) );
  MUX2_X1 U231 ( .A(\DRAM_mem[9][0] ), .B(\DRAM_mem[25][0] ), .S(Addr[4]), .Z(
        n197) );
  MUX2_X1 U232 ( .A(\DRAM_mem[1][0] ), .B(\DRAM_mem[17][0] ), .S(Addr[4]), .Z(
        n198) );
  MUX2_X1 U233 ( .A(n198), .B(n197), .S(n114), .Z(n199) );
  MUX2_X1 U234 ( .A(n199), .B(n196), .S(n102), .Z(n200) );
  MUX2_X1 U235 ( .A(\DRAM_mem[12][0] ), .B(\DRAM_mem[28][0] ), .S(n133), .Z(
        n201) );
  MUX2_X1 U236 ( .A(\DRAM_mem[4][0] ), .B(\DRAM_mem[20][0] ), .S(n133), .Z(
        n202) );
  MUX2_X1 U237 ( .A(n202), .B(n201), .S(n114), .Z(n203) );
  MUX2_X1 U238 ( .A(\DRAM_mem[8][0] ), .B(\DRAM_mem[24][0] ), .S(n133), .Z(
        n204) );
  MUX2_X1 U239 ( .A(\DRAM_mem[0][0] ), .B(\DRAM_mem[16][0] ), .S(n133), .Z(
        n205) );
  MUX2_X1 U240 ( .A(n205), .B(n204), .S(n114), .Z(n206) );
  MUX2_X1 U241 ( .A(n206), .B(n203), .S(n102), .Z(n207) );
  MUX2_X1 U242 ( .A(n207), .B(n200), .S(Addr[0]), .Z(n208) );
  MUX2_X1 U243 ( .A(n208), .B(n193), .S(Addr[1]), .Z(N499) );
  MUX2_X1 U244 ( .A(\DRAM_mem[15][1] ), .B(\DRAM_mem[31][1] ), .S(n133), .Z(
        n209) );
  MUX2_X1 U245 ( .A(\DRAM_mem[7][1] ), .B(\DRAM_mem[23][1] ), .S(n133), .Z(
        n210) );
  MUX2_X1 U246 ( .A(n210), .B(n209), .S(n114), .Z(n211) );
  MUX2_X1 U247 ( .A(\DRAM_mem[11][1] ), .B(\DRAM_mem[27][1] ), .S(n133), .Z(
        n212) );
  MUX2_X1 U248 ( .A(\DRAM_mem[3][1] ), .B(\DRAM_mem[19][1] ), .S(n133), .Z(
        n213) );
  MUX2_X1 U249 ( .A(n213), .B(n212), .S(n114), .Z(n214) );
  MUX2_X1 U250 ( .A(n214), .B(n211), .S(n102), .Z(n215) );
  MUX2_X1 U251 ( .A(\DRAM_mem[14][1] ), .B(\DRAM_mem[30][1] ), .S(n133), .Z(
        n216) );
  MUX2_X1 U252 ( .A(\DRAM_mem[6][1] ), .B(\DRAM_mem[22][1] ), .S(n133), .Z(
        n217) );
  MUX2_X1 U253 ( .A(n217), .B(n216), .S(n114), .Z(n218) );
  MUX2_X1 U254 ( .A(\DRAM_mem[10][1] ), .B(\DRAM_mem[26][1] ), .S(n133), .Z(
        n219) );
  MUX2_X1 U255 ( .A(\DRAM_mem[2][1] ), .B(\DRAM_mem[18][1] ), .S(n133), .Z(
        n220) );
  MUX2_X1 U256 ( .A(n220), .B(n219), .S(n114), .Z(n221) );
  MUX2_X1 U257 ( .A(n221), .B(n218), .S(n102), .Z(n222) );
  MUX2_X1 U258 ( .A(n222), .B(n215), .S(Addr[0]), .Z(n223) );
  MUX2_X1 U259 ( .A(\DRAM_mem[13][1] ), .B(\DRAM_mem[29][1] ), .S(n134), .Z(
        n224) );
  MUX2_X1 U260 ( .A(\DRAM_mem[5][1] ), .B(\DRAM_mem[21][1] ), .S(n134), .Z(
        n225) );
  MUX2_X1 U261 ( .A(n225), .B(n224), .S(n115), .Z(n226) );
  MUX2_X1 U262 ( .A(\DRAM_mem[9][1] ), .B(\DRAM_mem[25][1] ), .S(n134), .Z(
        n227) );
  MUX2_X1 U263 ( .A(\DRAM_mem[1][1] ), .B(\DRAM_mem[17][1] ), .S(n134), .Z(
        n228) );
  MUX2_X1 U264 ( .A(n228), .B(n227), .S(n115), .Z(n229) );
  MUX2_X1 U265 ( .A(n229), .B(n226), .S(n102), .Z(n230) );
  MUX2_X1 U266 ( .A(\DRAM_mem[12][1] ), .B(\DRAM_mem[28][1] ), .S(n134), .Z(
        n231) );
  MUX2_X1 U267 ( .A(\DRAM_mem[4][1] ), .B(\DRAM_mem[20][1] ), .S(n134), .Z(
        n232) );
  MUX2_X1 U268 ( .A(n232), .B(n231), .S(n115), .Z(n233) );
  MUX2_X1 U269 ( .A(\DRAM_mem[8][1] ), .B(\DRAM_mem[24][1] ), .S(n134), .Z(
        n234) );
  MUX2_X1 U270 ( .A(\DRAM_mem[0][1] ), .B(\DRAM_mem[16][1] ), .S(n134), .Z(
        n235) );
  MUX2_X1 U271 ( .A(n235), .B(n234), .S(n115), .Z(n236) );
  MUX2_X1 U272 ( .A(n236), .B(n233), .S(n102), .Z(n237) );
  MUX2_X1 U273 ( .A(n237), .B(n230), .S(Addr[0]), .Z(n238) );
  MUX2_X1 U274 ( .A(n238), .B(n223), .S(Addr[1]), .Z(N498) );
  MUX2_X1 U275 ( .A(\DRAM_mem[15][2] ), .B(\DRAM_mem[31][2] ), .S(n134), .Z(
        n239) );
  MUX2_X1 U276 ( .A(\DRAM_mem[7][2] ), .B(\DRAM_mem[23][2] ), .S(n134), .Z(
        n240) );
  MUX2_X1 U277 ( .A(n240), .B(n239), .S(n115), .Z(n241) );
  MUX2_X1 U278 ( .A(\DRAM_mem[11][2] ), .B(\DRAM_mem[27][2] ), .S(n134), .Z(
        n242) );
  MUX2_X1 U279 ( .A(\DRAM_mem[3][2] ), .B(\DRAM_mem[19][2] ), .S(n134), .Z(
        n243) );
  MUX2_X1 U280 ( .A(n243), .B(n242), .S(n115), .Z(n244) );
  MUX2_X1 U281 ( .A(n244), .B(n241), .S(n102), .Z(n245) );
  MUX2_X1 U282 ( .A(\DRAM_mem[14][2] ), .B(\DRAM_mem[30][2] ), .S(n135), .Z(
        n246) );
  MUX2_X1 U283 ( .A(\DRAM_mem[6][2] ), .B(\DRAM_mem[22][2] ), .S(n135), .Z(
        n247) );
  MUX2_X1 U284 ( .A(n247), .B(n246), .S(n115), .Z(n248) );
  MUX2_X1 U285 ( .A(\DRAM_mem[10][2] ), .B(\DRAM_mem[26][2] ), .S(n135), .Z(
        n249) );
  MUX2_X1 U286 ( .A(\DRAM_mem[2][2] ), .B(\DRAM_mem[18][2] ), .S(n135), .Z(
        n250) );
  MUX2_X1 U287 ( .A(n250), .B(n249), .S(n115), .Z(n251) );
  MUX2_X1 U288 ( .A(n251), .B(n248), .S(n102), .Z(n252) );
  MUX2_X1 U289 ( .A(n252), .B(n245), .S(Addr[0]), .Z(n253) );
  MUX2_X1 U290 ( .A(\DRAM_mem[13][2] ), .B(\DRAM_mem[29][2] ), .S(n135), .Z(
        n254) );
  MUX2_X1 U291 ( .A(\DRAM_mem[5][2] ), .B(\DRAM_mem[21][2] ), .S(n135), .Z(
        n255) );
  MUX2_X1 U292 ( .A(n255), .B(n254), .S(n115), .Z(n256) );
  MUX2_X1 U293 ( .A(\DRAM_mem[9][2] ), .B(\DRAM_mem[25][2] ), .S(n135), .Z(
        n257) );
  MUX2_X1 U294 ( .A(\DRAM_mem[1][2] ), .B(\DRAM_mem[17][2] ), .S(n135), .Z(
        n258) );
  MUX2_X1 U295 ( .A(n258), .B(n257), .S(n115), .Z(n259) );
  MUX2_X1 U296 ( .A(n259), .B(n256), .S(n102), .Z(n260) );
  MUX2_X1 U297 ( .A(\DRAM_mem[12][2] ), .B(\DRAM_mem[28][2] ), .S(n135), .Z(
        n261) );
  MUX2_X1 U298 ( .A(\DRAM_mem[4][2] ), .B(\DRAM_mem[20][2] ), .S(n135), .Z(
        n262) );
  MUX2_X1 U299 ( .A(n262), .B(n261), .S(n115), .Z(n263) );
  MUX2_X1 U300 ( .A(\DRAM_mem[8][2] ), .B(\DRAM_mem[24][2] ), .S(n135), .Z(
        n264) );
  MUX2_X1 U301 ( .A(\DRAM_mem[0][2] ), .B(\DRAM_mem[16][2] ), .S(n135), .Z(
        n265) );
  MUX2_X1 U302 ( .A(n265), .B(n264), .S(n115), .Z(n266) );
  MUX2_X1 U303 ( .A(n266), .B(n263), .S(n102), .Z(n267) );
  MUX2_X1 U304 ( .A(n267), .B(n260), .S(Addr[0]), .Z(n268) );
  MUX2_X1 U305 ( .A(n268), .B(n253), .S(Addr[1]), .Z(N497) );
  MUX2_X1 U306 ( .A(\DRAM_mem[15][3] ), .B(\DRAM_mem[31][3] ), .S(n136), .Z(
        n269) );
  MUX2_X1 U307 ( .A(\DRAM_mem[7][3] ), .B(\DRAM_mem[23][3] ), .S(n136), .Z(
        n270) );
  MUX2_X1 U308 ( .A(n270), .B(n269), .S(n116), .Z(n271) );
  MUX2_X1 U309 ( .A(\DRAM_mem[11][3] ), .B(\DRAM_mem[27][3] ), .S(n136), .Z(
        n272) );
  MUX2_X1 U310 ( .A(\DRAM_mem[3][3] ), .B(\DRAM_mem[19][3] ), .S(n136), .Z(
        n273) );
  MUX2_X1 U311 ( .A(n273), .B(n272), .S(n116), .Z(n274) );
  MUX2_X1 U312 ( .A(n274), .B(n271), .S(n103), .Z(n275) );
  MUX2_X1 U313 ( .A(\DRAM_mem[14][3] ), .B(\DRAM_mem[30][3] ), .S(n136), .Z(
        n276) );
  MUX2_X1 U314 ( .A(\DRAM_mem[6][3] ), .B(\DRAM_mem[22][3] ), .S(n136), .Z(
        n277) );
  MUX2_X1 U315 ( .A(n277), .B(n276), .S(n116), .Z(n278) );
  MUX2_X1 U316 ( .A(\DRAM_mem[10][3] ), .B(\DRAM_mem[26][3] ), .S(n136), .Z(
        n279) );
  MUX2_X1 U317 ( .A(\DRAM_mem[2][3] ), .B(\DRAM_mem[18][3] ), .S(n136), .Z(
        n280) );
  MUX2_X1 U318 ( .A(n280), .B(n279), .S(n116), .Z(n281) );
  MUX2_X1 U319 ( .A(n281), .B(n278), .S(n103), .Z(n282) );
  MUX2_X1 U320 ( .A(n282), .B(n275), .S(Addr[0]), .Z(n283) );
  MUX2_X1 U321 ( .A(\DRAM_mem[13][3] ), .B(\DRAM_mem[29][3] ), .S(n136), .Z(
        n284) );
  MUX2_X1 U322 ( .A(\DRAM_mem[5][3] ), .B(\DRAM_mem[21][3] ), .S(n136), .Z(
        n285) );
  MUX2_X1 U323 ( .A(n285), .B(n284), .S(n116), .Z(n286) );
  MUX2_X1 U324 ( .A(\DRAM_mem[9][3] ), .B(\DRAM_mem[25][3] ), .S(n136), .Z(
        n287) );
  MUX2_X1 U325 ( .A(\DRAM_mem[1][3] ), .B(\DRAM_mem[17][3] ), .S(n136), .Z(
        n288) );
  MUX2_X1 U326 ( .A(n288), .B(n287), .S(n116), .Z(n289) );
  MUX2_X1 U327 ( .A(n289), .B(n286), .S(n103), .Z(n290) );
  MUX2_X1 U328 ( .A(\DRAM_mem[12][3] ), .B(\DRAM_mem[28][3] ), .S(n137), .Z(
        n291) );
  MUX2_X1 U329 ( .A(\DRAM_mem[4][3] ), .B(\DRAM_mem[20][3] ), .S(n137), .Z(
        n292) );
  MUX2_X1 U330 ( .A(n292), .B(n291), .S(n116), .Z(n293) );
  MUX2_X1 U331 ( .A(\DRAM_mem[8][3] ), .B(\DRAM_mem[24][3] ), .S(n137), .Z(
        n294) );
  MUX2_X1 U332 ( .A(\DRAM_mem[0][3] ), .B(\DRAM_mem[16][3] ), .S(n137), .Z(
        n295) );
  MUX2_X1 U333 ( .A(n295), .B(n294), .S(n116), .Z(n296) );
  MUX2_X1 U334 ( .A(n296), .B(n293), .S(n103), .Z(n297) );
  MUX2_X1 U335 ( .A(n297), .B(n290), .S(Addr[0]), .Z(n298) );
  MUX2_X1 U336 ( .A(n298), .B(n283), .S(Addr[1]), .Z(N496) );
  MUX2_X1 U337 ( .A(\DRAM_mem[15][4] ), .B(\DRAM_mem[31][4] ), .S(n137), .Z(
        n299) );
  MUX2_X1 U338 ( .A(\DRAM_mem[7][4] ), .B(\DRAM_mem[23][4] ), .S(n137), .Z(
        n300) );
  MUX2_X1 U339 ( .A(n300), .B(n299), .S(n116), .Z(n301) );
  MUX2_X1 U340 ( .A(\DRAM_mem[11][4] ), .B(\DRAM_mem[27][4] ), .S(n137), .Z(
        n302) );
  MUX2_X1 U341 ( .A(\DRAM_mem[3][4] ), .B(\DRAM_mem[19][4] ), .S(n137), .Z(
        n303) );
  MUX2_X1 U342 ( .A(n303), .B(n302), .S(n116), .Z(n304) );
  MUX2_X1 U343 ( .A(n304), .B(n301), .S(n103), .Z(n305) );
  MUX2_X1 U344 ( .A(\DRAM_mem[14][4] ), .B(\DRAM_mem[30][4] ), .S(n137), .Z(
        n306) );
  MUX2_X1 U345 ( .A(\DRAM_mem[6][4] ), .B(\DRAM_mem[22][4] ), .S(n137), .Z(
        n307) );
  MUX2_X1 U346 ( .A(n307), .B(n306), .S(n116), .Z(n308) );
  MUX2_X1 U347 ( .A(\DRAM_mem[10][4] ), .B(\DRAM_mem[26][4] ), .S(n137), .Z(
        n309) );
  MUX2_X1 U348 ( .A(\DRAM_mem[2][4] ), .B(\DRAM_mem[18][4] ), .S(n137), .Z(
        n310) );
  MUX2_X1 U349 ( .A(n310), .B(n309), .S(n116), .Z(n311) );
  MUX2_X1 U350 ( .A(n311), .B(n308), .S(n103), .Z(n312) );
  MUX2_X1 U351 ( .A(n312), .B(n305), .S(Addr[0]), .Z(n313) );
  MUX2_X1 U352 ( .A(\DRAM_mem[13][4] ), .B(\DRAM_mem[29][4] ), .S(n138), .Z(
        n314) );
  MUX2_X1 U353 ( .A(\DRAM_mem[5][4] ), .B(\DRAM_mem[21][4] ), .S(n138), .Z(
        n315) );
  MUX2_X1 U354 ( .A(n315), .B(n314), .S(n117), .Z(n316) );
  MUX2_X1 U355 ( .A(\DRAM_mem[9][4] ), .B(\DRAM_mem[25][4] ), .S(n138), .Z(
        n317) );
  MUX2_X1 U356 ( .A(\DRAM_mem[1][4] ), .B(\DRAM_mem[17][4] ), .S(n138), .Z(
        n318) );
  MUX2_X1 U357 ( .A(n318), .B(n317), .S(n117), .Z(n319) );
  MUX2_X1 U358 ( .A(n319), .B(n316), .S(n103), .Z(n320) );
  MUX2_X1 U359 ( .A(\DRAM_mem[12][4] ), .B(\DRAM_mem[28][4] ), .S(n138), .Z(
        n321) );
  MUX2_X1 U360 ( .A(\DRAM_mem[4][4] ), .B(\DRAM_mem[20][4] ), .S(n138), .Z(
        n322) );
  MUX2_X1 U361 ( .A(n322), .B(n321), .S(n117), .Z(n323) );
  MUX2_X1 U362 ( .A(\DRAM_mem[8][4] ), .B(\DRAM_mem[24][4] ), .S(n138), .Z(
        n324) );
  MUX2_X1 U363 ( .A(\DRAM_mem[0][4] ), .B(\DRAM_mem[16][4] ), .S(n138), .Z(
        n325) );
  MUX2_X1 U364 ( .A(n325), .B(n324), .S(n117), .Z(n326) );
  MUX2_X1 U365 ( .A(n326), .B(n323), .S(n103), .Z(n327) );
  MUX2_X1 U366 ( .A(n327), .B(n320), .S(Addr[0]), .Z(n328) );
  MUX2_X1 U367 ( .A(n328), .B(n313), .S(Addr[1]), .Z(N495) );
  MUX2_X1 U368 ( .A(\DRAM_mem[15][5] ), .B(\DRAM_mem[31][5] ), .S(n138), .Z(
        n329) );
  MUX2_X1 U369 ( .A(\DRAM_mem[7][5] ), .B(\DRAM_mem[23][5] ), .S(n138), .Z(
        n330) );
  MUX2_X1 U370 ( .A(n330), .B(n329), .S(n117), .Z(n331) );
  MUX2_X1 U371 ( .A(\DRAM_mem[11][5] ), .B(\DRAM_mem[27][5] ), .S(n138), .Z(
        n332) );
  MUX2_X1 U372 ( .A(\DRAM_mem[3][5] ), .B(\DRAM_mem[19][5] ), .S(n138), .Z(
        n333) );
  MUX2_X1 U373 ( .A(n333), .B(n332), .S(n117), .Z(n334) );
  MUX2_X1 U374 ( .A(n334), .B(n331), .S(n103), .Z(n335) );
  MUX2_X1 U375 ( .A(\DRAM_mem[14][5] ), .B(\DRAM_mem[30][5] ), .S(n139), .Z(
        n336) );
  MUX2_X1 U376 ( .A(\DRAM_mem[6][5] ), .B(\DRAM_mem[22][5] ), .S(n139), .Z(
        n337) );
  MUX2_X1 U377 ( .A(n337), .B(n336), .S(n117), .Z(n338) );
  MUX2_X1 U378 ( .A(\DRAM_mem[10][5] ), .B(\DRAM_mem[26][5] ), .S(n139), .Z(
        n339) );
  MUX2_X1 U379 ( .A(\DRAM_mem[2][5] ), .B(\DRAM_mem[18][5] ), .S(n139), .Z(
        n340) );
  MUX2_X1 U380 ( .A(n340), .B(n339), .S(n117), .Z(n341) );
  MUX2_X1 U381 ( .A(n341), .B(n338), .S(n103), .Z(n342) );
  MUX2_X1 U382 ( .A(n342), .B(n335), .S(Addr[0]), .Z(n343) );
  MUX2_X1 U383 ( .A(\DRAM_mem[13][5] ), .B(\DRAM_mem[29][5] ), .S(n139), .Z(
        n344) );
  MUX2_X1 U384 ( .A(\DRAM_mem[5][5] ), .B(\DRAM_mem[21][5] ), .S(n139), .Z(
        n345) );
  MUX2_X1 U385 ( .A(n345), .B(n344), .S(n117), .Z(n346) );
  MUX2_X1 U386 ( .A(\DRAM_mem[9][5] ), .B(\DRAM_mem[25][5] ), .S(n139), .Z(
        n347) );
  MUX2_X1 U387 ( .A(\DRAM_mem[1][5] ), .B(\DRAM_mem[17][5] ), .S(n139), .Z(
        n348) );
  MUX2_X1 U388 ( .A(n348), .B(n347), .S(n117), .Z(n349) );
  MUX2_X1 U389 ( .A(n349), .B(n346), .S(n103), .Z(n350) );
  MUX2_X1 U390 ( .A(\DRAM_mem[12][5] ), .B(\DRAM_mem[28][5] ), .S(n139), .Z(
        n351) );
  MUX2_X1 U391 ( .A(\DRAM_mem[4][5] ), .B(\DRAM_mem[20][5] ), .S(n139), .Z(
        n352) );
  MUX2_X1 U392 ( .A(n352), .B(n351), .S(n117), .Z(n353) );
  MUX2_X1 U393 ( .A(\DRAM_mem[8][5] ), .B(\DRAM_mem[24][5] ), .S(n139), .Z(
        n354) );
  MUX2_X1 U394 ( .A(\DRAM_mem[0][5] ), .B(\DRAM_mem[16][5] ), .S(n139), .Z(
        n355) );
  MUX2_X1 U395 ( .A(n355), .B(n354), .S(n117), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n353), .S(n103), .Z(n357) );
  MUX2_X1 U397 ( .A(n357), .B(n350), .S(Addr[0]), .Z(n358) );
  MUX2_X1 U398 ( .A(n358), .B(n343), .S(Addr[1]), .Z(N494) );
  MUX2_X1 U399 ( .A(\DRAM_mem[15][6] ), .B(\DRAM_mem[31][6] ), .S(n140), .Z(
        n359) );
  MUX2_X1 U400 ( .A(\DRAM_mem[7][6] ), .B(\DRAM_mem[23][6] ), .S(n140), .Z(
        n360) );
  MUX2_X1 U401 ( .A(n360), .B(n359), .S(n118), .Z(n361) );
  MUX2_X1 U402 ( .A(\DRAM_mem[11][6] ), .B(\DRAM_mem[27][6] ), .S(n140), .Z(
        n362) );
  MUX2_X1 U403 ( .A(\DRAM_mem[3][6] ), .B(\DRAM_mem[19][6] ), .S(n140), .Z(
        n363) );
  MUX2_X1 U404 ( .A(n363), .B(n362), .S(n118), .Z(n364) );
  MUX2_X1 U405 ( .A(n364), .B(n361), .S(n104), .Z(n365) );
  MUX2_X1 U406 ( .A(\DRAM_mem[14][6] ), .B(\DRAM_mem[30][6] ), .S(n140), .Z(
        n366) );
  MUX2_X1 U407 ( .A(\DRAM_mem[6][6] ), .B(\DRAM_mem[22][6] ), .S(n140), .Z(
        n367) );
  MUX2_X1 U408 ( .A(n367), .B(n366), .S(n118), .Z(n368) );
  MUX2_X1 U409 ( .A(\DRAM_mem[10][6] ), .B(\DRAM_mem[26][6] ), .S(n140), .Z(
        n369) );
  MUX2_X1 U410 ( .A(\DRAM_mem[2][6] ), .B(\DRAM_mem[18][6] ), .S(n140), .Z(
        n370) );
  MUX2_X1 U411 ( .A(n370), .B(n369), .S(n118), .Z(n371) );
  MUX2_X1 U412 ( .A(n371), .B(n368), .S(n104), .Z(n372) );
  MUX2_X1 U413 ( .A(n372), .B(n365), .S(Addr[0]), .Z(n373) );
  MUX2_X1 U414 ( .A(\DRAM_mem[13][6] ), .B(\DRAM_mem[29][6] ), .S(n140), .Z(
        n374) );
  MUX2_X1 U415 ( .A(\DRAM_mem[5][6] ), .B(\DRAM_mem[21][6] ), .S(n140), .Z(
        n375) );
  MUX2_X1 U416 ( .A(n375), .B(n374), .S(n118), .Z(n376) );
  MUX2_X1 U417 ( .A(\DRAM_mem[9][6] ), .B(\DRAM_mem[25][6] ), .S(n140), .Z(
        n377) );
  MUX2_X1 U418 ( .A(\DRAM_mem[1][6] ), .B(\DRAM_mem[17][6] ), .S(n140), .Z(
        n378) );
  MUX2_X1 U419 ( .A(n378), .B(n377), .S(n118), .Z(n379) );
  MUX2_X1 U420 ( .A(n379), .B(n376), .S(n104), .Z(n380) );
  MUX2_X1 U421 ( .A(\DRAM_mem[12][6] ), .B(\DRAM_mem[28][6] ), .S(n141), .Z(
        n381) );
  MUX2_X1 U422 ( .A(\DRAM_mem[4][6] ), .B(\DRAM_mem[20][6] ), .S(n141), .Z(
        n382) );
  MUX2_X1 U423 ( .A(n382), .B(n381), .S(n118), .Z(n383) );
  MUX2_X1 U424 ( .A(\DRAM_mem[8][6] ), .B(\DRAM_mem[24][6] ), .S(n141), .Z(
        n384) );
  MUX2_X1 U425 ( .A(\DRAM_mem[0][6] ), .B(\DRAM_mem[16][6] ), .S(n141), .Z(
        n385) );
  MUX2_X1 U426 ( .A(n385), .B(n384), .S(n118), .Z(n386) );
  MUX2_X1 U427 ( .A(n386), .B(n383), .S(n104), .Z(n387) );
  MUX2_X1 U428 ( .A(n387), .B(n380), .S(Addr[0]), .Z(n388) );
  MUX2_X1 U429 ( .A(n388), .B(n373), .S(Addr[1]), .Z(N493) );
  MUX2_X1 U430 ( .A(\DRAM_mem[15][7] ), .B(\DRAM_mem[31][7] ), .S(n141), .Z(
        n389) );
  MUX2_X1 U431 ( .A(\DRAM_mem[7][7] ), .B(\DRAM_mem[23][7] ), .S(n141), .Z(
        n390) );
  MUX2_X1 U432 ( .A(n390), .B(n389), .S(n118), .Z(n391) );
  MUX2_X1 U433 ( .A(\DRAM_mem[11][7] ), .B(\DRAM_mem[27][7] ), .S(n141), .Z(
        n392) );
  MUX2_X1 U434 ( .A(\DRAM_mem[3][7] ), .B(\DRAM_mem[19][7] ), .S(n141), .Z(
        n393) );
  MUX2_X1 U435 ( .A(n393), .B(n392), .S(n118), .Z(n394) );
  MUX2_X1 U436 ( .A(n394), .B(n391), .S(n104), .Z(n395) );
  MUX2_X1 U437 ( .A(\DRAM_mem[14][7] ), .B(\DRAM_mem[30][7] ), .S(n141), .Z(
        n396) );
  MUX2_X1 U438 ( .A(\DRAM_mem[6][7] ), .B(\DRAM_mem[22][7] ), .S(n141), .Z(
        n397) );
  MUX2_X1 U439 ( .A(n397), .B(n396), .S(n118), .Z(n398) );
  MUX2_X1 U440 ( .A(\DRAM_mem[10][7] ), .B(\DRAM_mem[26][7] ), .S(n141), .Z(
        n399) );
  MUX2_X1 U441 ( .A(\DRAM_mem[2][7] ), .B(\DRAM_mem[18][7] ), .S(n141), .Z(
        n400) );
  MUX2_X1 U442 ( .A(n400), .B(n399), .S(n118), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n398), .S(n104), .Z(n402) );
  MUX2_X1 U444 ( .A(n402), .B(n395), .S(Addr[0]), .Z(n403) );
  MUX2_X1 U445 ( .A(\DRAM_mem[13][7] ), .B(\DRAM_mem[29][7] ), .S(n142), .Z(
        n404) );
  MUX2_X1 U446 ( .A(\DRAM_mem[5][7] ), .B(\DRAM_mem[21][7] ), .S(n142), .Z(
        n405) );
  MUX2_X1 U447 ( .A(n405), .B(n404), .S(n119), .Z(n406) );
  MUX2_X1 U448 ( .A(\DRAM_mem[9][7] ), .B(\DRAM_mem[25][7] ), .S(n142), .Z(
        n407) );
  MUX2_X1 U449 ( .A(\DRAM_mem[1][7] ), .B(\DRAM_mem[17][7] ), .S(n142), .Z(
        n408) );
  MUX2_X1 U450 ( .A(n408), .B(n407), .S(n119), .Z(n409) );
  MUX2_X1 U451 ( .A(n409), .B(n406), .S(n104), .Z(n410) );
  MUX2_X1 U452 ( .A(\DRAM_mem[12][7] ), .B(\DRAM_mem[28][7] ), .S(n142), .Z(
        n411) );
  MUX2_X1 U453 ( .A(\DRAM_mem[4][7] ), .B(\DRAM_mem[20][7] ), .S(n142), .Z(
        n412) );
  MUX2_X1 U454 ( .A(n412), .B(n411), .S(n119), .Z(n413) );
  MUX2_X1 U455 ( .A(\DRAM_mem[8][7] ), .B(\DRAM_mem[24][7] ), .S(n142), .Z(
        n414) );
  MUX2_X1 U456 ( .A(\DRAM_mem[0][7] ), .B(\DRAM_mem[16][7] ), .S(n142), .Z(
        n415) );
  MUX2_X1 U457 ( .A(n415), .B(n414), .S(n119), .Z(n416) );
  MUX2_X1 U458 ( .A(n416), .B(n413), .S(n104), .Z(n417) );
  MUX2_X1 U459 ( .A(n417), .B(n410), .S(Addr[0]), .Z(n418) );
  MUX2_X1 U460 ( .A(n418), .B(n403), .S(Addr[1]), .Z(N492) );
  MUX2_X1 U461 ( .A(\DRAM_mem[15][8] ), .B(\DRAM_mem[31][8] ), .S(n142), .Z(
        n419) );
  MUX2_X1 U462 ( .A(\DRAM_mem[7][8] ), .B(\DRAM_mem[23][8] ), .S(n142), .Z(
        n420) );
  MUX2_X1 U463 ( .A(n420), .B(n419), .S(n119), .Z(n421) );
  MUX2_X1 U464 ( .A(\DRAM_mem[11][8] ), .B(\DRAM_mem[27][8] ), .S(n142), .Z(
        n422) );
  MUX2_X1 U465 ( .A(\DRAM_mem[3][8] ), .B(\DRAM_mem[19][8] ), .S(n142), .Z(
        n423) );
  MUX2_X1 U466 ( .A(n423), .B(n422), .S(n119), .Z(n424) );
  MUX2_X1 U467 ( .A(n424), .B(n421), .S(n104), .Z(n425) );
  MUX2_X1 U468 ( .A(\DRAM_mem[14][8] ), .B(\DRAM_mem[30][8] ), .S(n143), .Z(
        n426) );
  MUX2_X1 U469 ( .A(\DRAM_mem[6][8] ), .B(\DRAM_mem[22][8] ), .S(n143), .Z(
        n427) );
  MUX2_X1 U470 ( .A(n427), .B(n426), .S(n119), .Z(n428) );
  MUX2_X1 U471 ( .A(\DRAM_mem[10][8] ), .B(\DRAM_mem[26][8] ), .S(n143), .Z(
        n429) );
  MUX2_X1 U472 ( .A(\DRAM_mem[2][8] ), .B(\DRAM_mem[18][8] ), .S(n143), .Z(
        n430) );
  MUX2_X1 U473 ( .A(n430), .B(n429), .S(n119), .Z(n431) );
  MUX2_X1 U474 ( .A(n431), .B(n428), .S(n104), .Z(n432) );
  MUX2_X1 U475 ( .A(n432), .B(n425), .S(Addr[0]), .Z(n433) );
  MUX2_X1 U476 ( .A(\DRAM_mem[13][8] ), .B(\DRAM_mem[29][8] ), .S(n143), .Z(
        n434) );
  MUX2_X1 U477 ( .A(\DRAM_mem[5][8] ), .B(\DRAM_mem[21][8] ), .S(n143), .Z(
        n435) );
  MUX2_X1 U478 ( .A(n435), .B(n434), .S(n119), .Z(n436) );
  MUX2_X1 U479 ( .A(\DRAM_mem[9][8] ), .B(\DRAM_mem[25][8] ), .S(n143), .Z(
        n437) );
  MUX2_X1 U480 ( .A(\DRAM_mem[1][8] ), .B(\DRAM_mem[17][8] ), .S(n143), .Z(
        n438) );
  MUX2_X1 U481 ( .A(n438), .B(n437), .S(n119), .Z(n439) );
  MUX2_X1 U482 ( .A(n439), .B(n436), .S(n104), .Z(n440) );
  MUX2_X1 U483 ( .A(\DRAM_mem[12][8] ), .B(\DRAM_mem[28][8] ), .S(n143), .Z(
        n441) );
  MUX2_X1 U484 ( .A(\DRAM_mem[4][8] ), .B(\DRAM_mem[20][8] ), .S(n143), .Z(
        n442) );
  MUX2_X1 U485 ( .A(n442), .B(n441), .S(n119), .Z(n443) );
  MUX2_X1 U486 ( .A(\DRAM_mem[8][8] ), .B(\DRAM_mem[24][8] ), .S(n143), .Z(
        n444) );
  MUX2_X1 U487 ( .A(\DRAM_mem[0][8] ), .B(\DRAM_mem[16][8] ), .S(n143), .Z(
        n445) );
  MUX2_X1 U488 ( .A(n445), .B(n444), .S(n119), .Z(n446) );
  MUX2_X1 U489 ( .A(n446), .B(n443), .S(n104), .Z(n447) );
  MUX2_X1 U490 ( .A(n447), .B(n440), .S(Addr[0]), .Z(n448) );
  MUX2_X1 U491 ( .A(n448), .B(n433), .S(Addr[1]), .Z(N491) );
  MUX2_X1 U492 ( .A(\DRAM_mem[15][9] ), .B(\DRAM_mem[31][9] ), .S(n144), .Z(
        n449) );
  MUX2_X1 U493 ( .A(\DRAM_mem[7][9] ), .B(\DRAM_mem[23][9] ), .S(n144), .Z(
        n450) );
  MUX2_X1 U494 ( .A(n450), .B(n449), .S(n120), .Z(n451) );
  MUX2_X1 U495 ( .A(\DRAM_mem[11][9] ), .B(\DRAM_mem[27][9] ), .S(n144), .Z(
        n452) );
  MUX2_X1 U496 ( .A(\DRAM_mem[3][9] ), .B(\DRAM_mem[19][9] ), .S(n144), .Z(
        n453) );
  MUX2_X1 U497 ( .A(n453), .B(n452), .S(n120), .Z(n454) );
  MUX2_X1 U498 ( .A(n454), .B(n451), .S(n105), .Z(n455) );
  MUX2_X1 U499 ( .A(\DRAM_mem[14][9] ), .B(\DRAM_mem[30][9] ), .S(n144), .Z(
        n456) );
  MUX2_X1 U500 ( .A(\DRAM_mem[6][9] ), .B(\DRAM_mem[22][9] ), .S(n144), .Z(
        n457) );
  MUX2_X1 U501 ( .A(n457), .B(n456), .S(n120), .Z(n458) );
  MUX2_X1 U502 ( .A(\DRAM_mem[10][9] ), .B(\DRAM_mem[26][9] ), .S(n144), .Z(
        n459) );
  MUX2_X1 U503 ( .A(\DRAM_mem[2][9] ), .B(\DRAM_mem[18][9] ), .S(n144), .Z(
        n460) );
  MUX2_X1 U504 ( .A(n460), .B(n459), .S(n120), .Z(n461) );
  MUX2_X1 U505 ( .A(n461), .B(n458), .S(n105), .Z(n462) );
  MUX2_X1 U506 ( .A(n462), .B(n455), .S(Addr[0]), .Z(n463) );
  MUX2_X1 U507 ( .A(\DRAM_mem[13][9] ), .B(\DRAM_mem[29][9] ), .S(n144), .Z(
        n464) );
  MUX2_X1 U508 ( .A(\DRAM_mem[5][9] ), .B(\DRAM_mem[21][9] ), .S(n144), .Z(
        n465) );
  MUX2_X1 U509 ( .A(n465), .B(n464), .S(n120), .Z(n466) );
  MUX2_X1 U510 ( .A(\DRAM_mem[9][9] ), .B(\DRAM_mem[25][9] ), .S(n144), .Z(
        n467) );
  MUX2_X1 U511 ( .A(\DRAM_mem[1][9] ), .B(\DRAM_mem[17][9] ), .S(n144), .Z(
        n468) );
  MUX2_X1 U512 ( .A(n468), .B(n467), .S(n120), .Z(n469) );
  MUX2_X1 U513 ( .A(n469), .B(n466), .S(n105), .Z(n470) );
  MUX2_X1 U514 ( .A(\DRAM_mem[12][9] ), .B(\DRAM_mem[28][9] ), .S(n145), .Z(
        n471) );
  MUX2_X1 U515 ( .A(\DRAM_mem[4][9] ), .B(\DRAM_mem[20][9] ), .S(n145), .Z(
        n472) );
  MUX2_X1 U516 ( .A(n472), .B(n471), .S(n120), .Z(n473) );
  MUX2_X1 U517 ( .A(\DRAM_mem[8][9] ), .B(\DRAM_mem[24][9] ), .S(n145), .Z(
        n474) );
  MUX2_X1 U518 ( .A(\DRAM_mem[0][9] ), .B(\DRAM_mem[16][9] ), .S(n145), .Z(
        n475) );
  MUX2_X1 U519 ( .A(n475), .B(n474), .S(n120), .Z(n476) );
  MUX2_X1 U520 ( .A(n476), .B(n473), .S(n105), .Z(n477) );
  MUX2_X1 U521 ( .A(n477), .B(n470), .S(Addr[0]), .Z(n478) );
  MUX2_X1 U522 ( .A(n478), .B(n463), .S(Addr[1]), .Z(N490) );
  MUX2_X1 U523 ( .A(\DRAM_mem[15][10] ), .B(\DRAM_mem[31][10] ), .S(n145), .Z(
        n479) );
  MUX2_X1 U524 ( .A(\DRAM_mem[7][10] ), .B(\DRAM_mem[23][10] ), .S(n145), .Z(
        n480) );
  MUX2_X1 U525 ( .A(n480), .B(n479), .S(n120), .Z(n481) );
  MUX2_X1 U526 ( .A(\DRAM_mem[11][10] ), .B(\DRAM_mem[27][10] ), .S(n145), .Z(
        n482) );
  MUX2_X1 U527 ( .A(\DRAM_mem[3][10] ), .B(\DRAM_mem[19][10] ), .S(n145), .Z(
        n483) );
  MUX2_X1 U528 ( .A(n483), .B(n482), .S(n120), .Z(n484) );
  MUX2_X1 U529 ( .A(n484), .B(n481), .S(n105), .Z(n485) );
  MUX2_X1 U530 ( .A(\DRAM_mem[14][10] ), .B(\DRAM_mem[30][10] ), .S(n145), .Z(
        n486) );
  MUX2_X1 U531 ( .A(\DRAM_mem[6][10] ), .B(\DRAM_mem[22][10] ), .S(n145), .Z(
        n487) );
  MUX2_X1 U532 ( .A(n487), .B(n486), .S(n120), .Z(n488) );
  MUX2_X1 U533 ( .A(\DRAM_mem[10][10] ), .B(\DRAM_mem[26][10] ), .S(n145), .Z(
        n489) );
  MUX2_X1 U534 ( .A(\DRAM_mem[2][10] ), .B(\DRAM_mem[18][10] ), .S(n145), .Z(
        n490) );
  MUX2_X1 U535 ( .A(n490), .B(n489), .S(n120), .Z(n491) );
  MUX2_X1 U536 ( .A(n491), .B(n488), .S(n105), .Z(n492) );
  MUX2_X1 U537 ( .A(n492), .B(n485), .S(Addr[0]), .Z(n493) );
  MUX2_X1 U538 ( .A(\DRAM_mem[13][10] ), .B(\DRAM_mem[29][10] ), .S(n146), .Z(
        n494) );
  MUX2_X1 U539 ( .A(\DRAM_mem[5][10] ), .B(\DRAM_mem[21][10] ), .S(n146), .Z(
        n495) );
  MUX2_X1 U540 ( .A(n495), .B(n494), .S(n121), .Z(n496) );
  MUX2_X1 U541 ( .A(\DRAM_mem[9][10] ), .B(\DRAM_mem[25][10] ), .S(n146), .Z(
        n497) );
  MUX2_X1 U542 ( .A(\DRAM_mem[1][10] ), .B(\DRAM_mem[17][10] ), .S(n146), .Z(
        n498) );
  MUX2_X1 U543 ( .A(n498), .B(n497), .S(n121), .Z(n499) );
  MUX2_X1 U544 ( .A(n499), .B(n496), .S(n105), .Z(n500) );
  MUX2_X1 U545 ( .A(\DRAM_mem[12][10] ), .B(\DRAM_mem[28][10] ), .S(n146), .Z(
        n501) );
  MUX2_X1 U546 ( .A(\DRAM_mem[4][10] ), .B(\DRAM_mem[20][10] ), .S(n146), .Z(
        n502) );
  MUX2_X1 U547 ( .A(n502), .B(n501), .S(n121), .Z(n503) );
  MUX2_X1 U548 ( .A(\DRAM_mem[8][10] ), .B(\DRAM_mem[24][10] ), .S(n146), .Z(
        n504) );
  MUX2_X1 U549 ( .A(\DRAM_mem[0][10] ), .B(\DRAM_mem[16][10] ), .S(n146), .Z(
        n505) );
  MUX2_X1 U550 ( .A(n505), .B(n504), .S(n121), .Z(n506) );
  MUX2_X1 U551 ( .A(n506), .B(n503), .S(n105), .Z(n507) );
  MUX2_X1 U552 ( .A(n507), .B(n500), .S(Addr[0]), .Z(n508) );
  MUX2_X1 U553 ( .A(n508), .B(n493), .S(Addr[1]), .Z(N489) );
  MUX2_X1 U554 ( .A(\DRAM_mem[15][11] ), .B(\DRAM_mem[31][11] ), .S(n146), .Z(
        n509) );
  MUX2_X1 U555 ( .A(\DRAM_mem[7][11] ), .B(\DRAM_mem[23][11] ), .S(n146), .Z(
        n510) );
  MUX2_X1 U556 ( .A(n510), .B(n509), .S(n121), .Z(n511) );
  MUX2_X1 U557 ( .A(\DRAM_mem[11][11] ), .B(\DRAM_mem[27][11] ), .S(n146), .Z(
        n512) );
  MUX2_X1 U558 ( .A(\DRAM_mem[3][11] ), .B(\DRAM_mem[19][11] ), .S(n146), .Z(
        n513) );
  MUX2_X1 U559 ( .A(n513), .B(n512), .S(n121), .Z(n514) );
  MUX2_X1 U560 ( .A(n514), .B(n511), .S(n105), .Z(n515) );
  MUX2_X1 U561 ( .A(\DRAM_mem[14][11] ), .B(\DRAM_mem[30][11] ), .S(n147), .Z(
        n516) );
  MUX2_X1 U562 ( .A(\DRAM_mem[6][11] ), .B(\DRAM_mem[22][11] ), .S(n147), .Z(
        n517) );
  MUX2_X1 U563 ( .A(n517), .B(n516), .S(n121), .Z(n518) );
  MUX2_X1 U564 ( .A(\DRAM_mem[10][11] ), .B(\DRAM_mem[26][11] ), .S(n147), .Z(
        n519) );
  MUX2_X1 U565 ( .A(\DRAM_mem[2][11] ), .B(\DRAM_mem[18][11] ), .S(n147), .Z(
        n520) );
  MUX2_X1 U566 ( .A(n520), .B(n519), .S(n121), .Z(n521) );
  MUX2_X1 U567 ( .A(n521), .B(n518), .S(n105), .Z(n522) );
  MUX2_X1 U568 ( .A(n522), .B(n515), .S(Addr[0]), .Z(n523) );
  MUX2_X1 U569 ( .A(\DRAM_mem[13][11] ), .B(\DRAM_mem[29][11] ), .S(n147), .Z(
        n524) );
  MUX2_X1 U570 ( .A(\DRAM_mem[5][11] ), .B(\DRAM_mem[21][11] ), .S(n147), .Z(
        n525) );
  MUX2_X1 U571 ( .A(n525), .B(n524), .S(n121), .Z(n526) );
  MUX2_X1 U572 ( .A(\DRAM_mem[9][11] ), .B(\DRAM_mem[25][11] ), .S(n147), .Z(
        n527) );
  MUX2_X1 U573 ( .A(\DRAM_mem[1][11] ), .B(\DRAM_mem[17][11] ), .S(n147), .Z(
        n528) );
  MUX2_X1 U574 ( .A(n528), .B(n527), .S(n121), .Z(n529) );
  MUX2_X1 U575 ( .A(n529), .B(n526), .S(n105), .Z(n530) );
  MUX2_X1 U576 ( .A(\DRAM_mem[12][11] ), .B(\DRAM_mem[28][11] ), .S(n147), .Z(
        n531) );
  MUX2_X1 U577 ( .A(\DRAM_mem[4][11] ), .B(\DRAM_mem[20][11] ), .S(n147), .Z(
        n532) );
  MUX2_X1 U578 ( .A(n532), .B(n531), .S(n121), .Z(n533) );
  MUX2_X1 U579 ( .A(\DRAM_mem[8][11] ), .B(\DRAM_mem[24][11] ), .S(n147), .Z(
        n534) );
  MUX2_X1 U580 ( .A(\DRAM_mem[0][11] ), .B(\DRAM_mem[16][11] ), .S(n147), .Z(
        n535) );
  MUX2_X1 U581 ( .A(n535), .B(n534), .S(n121), .Z(n536) );
  MUX2_X1 U582 ( .A(n536), .B(n533), .S(n105), .Z(n537) );
  MUX2_X1 U583 ( .A(n537), .B(n530), .S(Addr[0]), .Z(n538) );
  MUX2_X1 U584 ( .A(n538), .B(n523), .S(Addr[1]), .Z(N488) );
  MUX2_X1 U585 ( .A(\DRAM_mem[15][12] ), .B(\DRAM_mem[31][12] ), .S(n148), .Z(
        n539) );
  MUX2_X1 U586 ( .A(\DRAM_mem[7][12] ), .B(\DRAM_mem[23][12] ), .S(n148), .Z(
        n540) );
  MUX2_X1 U587 ( .A(n540), .B(n539), .S(n122), .Z(n541) );
  MUX2_X1 U588 ( .A(\DRAM_mem[11][12] ), .B(\DRAM_mem[27][12] ), .S(n148), .Z(
        n542) );
  MUX2_X1 U589 ( .A(\DRAM_mem[3][12] ), .B(\DRAM_mem[19][12] ), .S(n148), .Z(
        n543) );
  MUX2_X1 U590 ( .A(n543), .B(n542), .S(n122), .Z(n544) );
  MUX2_X1 U591 ( .A(n544), .B(n541), .S(n106), .Z(n545) );
  MUX2_X1 U592 ( .A(\DRAM_mem[14][12] ), .B(\DRAM_mem[30][12] ), .S(n148), .Z(
        n546) );
  MUX2_X1 U593 ( .A(\DRAM_mem[6][12] ), .B(\DRAM_mem[22][12] ), .S(n148), .Z(
        n547) );
  MUX2_X1 U594 ( .A(n547), .B(n546), .S(n122), .Z(n548) );
  MUX2_X1 U595 ( .A(\DRAM_mem[10][12] ), .B(\DRAM_mem[26][12] ), .S(n148), .Z(
        n549) );
  MUX2_X1 U596 ( .A(\DRAM_mem[2][12] ), .B(\DRAM_mem[18][12] ), .S(n148), .Z(
        n550) );
  MUX2_X1 U597 ( .A(n550), .B(n549), .S(n122), .Z(n551) );
  MUX2_X1 U598 ( .A(n551), .B(n548), .S(n106), .Z(n552) );
  MUX2_X1 U599 ( .A(n552), .B(n545), .S(Addr[0]), .Z(n553) );
  MUX2_X1 U600 ( .A(\DRAM_mem[13][12] ), .B(\DRAM_mem[29][12] ), .S(n148), .Z(
        n554) );
  MUX2_X1 U601 ( .A(\DRAM_mem[5][12] ), .B(\DRAM_mem[21][12] ), .S(n148), .Z(
        n555) );
  MUX2_X1 U602 ( .A(n555), .B(n554), .S(n122), .Z(n556) );
  MUX2_X1 U603 ( .A(\DRAM_mem[9][12] ), .B(\DRAM_mem[25][12] ), .S(n148), .Z(
        n557) );
  MUX2_X1 U604 ( .A(\DRAM_mem[1][12] ), .B(\DRAM_mem[17][12] ), .S(n148), .Z(
        n558) );
  MUX2_X1 U605 ( .A(n558), .B(n557), .S(n122), .Z(n559) );
  MUX2_X1 U606 ( .A(n559), .B(n556), .S(n106), .Z(n560) );
  MUX2_X1 U607 ( .A(\DRAM_mem[12][12] ), .B(\DRAM_mem[28][12] ), .S(n149), .Z(
        n561) );
  MUX2_X1 U608 ( .A(\DRAM_mem[4][12] ), .B(\DRAM_mem[20][12] ), .S(n149), .Z(
        n562) );
  MUX2_X1 U609 ( .A(n562), .B(n561), .S(n122), .Z(n563) );
  MUX2_X1 U610 ( .A(\DRAM_mem[8][12] ), .B(\DRAM_mem[24][12] ), .S(n149), .Z(
        n564) );
  MUX2_X1 U611 ( .A(\DRAM_mem[0][12] ), .B(\DRAM_mem[16][12] ), .S(n149), .Z(
        n565) );
  MUX2_X1 U612 ( .A(n565), .B(n564), .S(n122), .Z(n566) );
  MUX2_X1 U613 ( .A(n566), .B(n563), .S(n106), .Z(n567) );
  MUX2_X1 U614 ( .A(n567), .B(n560), .S(Addr[0]), .Z(n568) );
  MUX2_X1 U615 ( .A(n568), .B(n553), .S(Addr[1]), .Z(N487) );
  MUX2_X1 U616 ( .A(\DRAM_mem[15][13] ), .B(\DRAM_mem[31][13] ), .S(n149), .Z(
        n569) );
  MUX2_X1 U617 ( .A(\DRAM_mem[7][13] ), .B(\DRAM_mem[23][13] ), .S(n149), .Z(
        n570) );
  MUX2_X1 U618 ( .A(n570), .B(n569), .S(n122), .Z(n571) );
  MUX2_X1 U619 ( .A(\DRAM_mem[11][13] ), .B(\DRAM_mem[27][13] ), .S(n149), .Z(
        n572) );
  MUX2_X1 U620 ( .A(\DRAM_mem[3][13] ), .B(\DRAM_mem[19][13] ), .S(n149), .Z(
        n573) );
  MUX2_X1 U621 ( .A(n573), .B(n572), .S(n122), .Z(n574) );
  MUX2_X1 U622 ( .A(n574), .B(n571), .S(n106), .Z(n575) );
  MUX2_X1 U623 ( .A(\DRAM_mem[14][13] ), .B(\DRAM_mem[30][13] ), .S(n149), .Z(
        n576) );
  MUX2_X1 U624 ( .A(\DRAM_mem[6][13] ), .B(\DRAM_mem[22][13] ), .S(n149), .Z(
        n577) );
  MUX2_X1 U625 ( .A(n577), .B(n576), .S(n122), .Z(n578) );
  MUX2_X1 U626 ( .A(\DRAM_mem[10][13] ), .B(\DRAM_mem[26][13] ), .S(n149), .Z(
        n579) );
  MUX2_X1 U627 ( .A(\DRAM_mem[2][13] ), .B(\DRAM_mem[18][13] ), .S(n149), .Z(
        n580) );
  MUX2_X1 U628 ( .A(n580), .B(n579), .S(n122), .Z(n581) );
  MUX2_X1 U629 ( .A(n581), .B(n578), .S(n106), .Z(n582) );
  MUX2_X1 U630 ( .A(n582), .B(n575), .S(Addr[0]), .Z(n583) );
  MUX2_X1 U631 ( .A(\DRAM_mem[13][13] ), .B(\DRAM_mem[29][13] ), .S(n150), .Z(
        n584) );
  MUX2_X1 U632 ( .A(\DRAM_mem[5][13] ), .B(\DRAM_mem[21][13] ), .S(n150), .Z(
        n585) );
  MUX2_X1 U633 ( .A(n585), .B(n584), .S(n123), .Z(n586) );
  MUX2_X1 U634 ( .A(\DRAM_mem[9][13] ), .B(\DRAM_mem[25][13] ), .S(n150), .Z(
        n587) );
  MUX2_X1 U635 ( .A(\DRAM_mem[1][13] ), .B(\DRAM_mem[17][13] ), .S(n150), .Z(
        n588) );
  MUX2_X1 U636 ( .A(n588), .B(n587), .S(n123), .Z(n589) );
  MUX2_X1 U637 ( .A(n589), .B(n586), .S(n106), .Z(n590) );
  MUX2_X1 U638 ( .A(\DRAM_mem[12][13] ), .B(\DRAM_mem[28][13] ), .S(n150), .Z(
        n591) );
  MUX2_X1 U639 ( .A(\DRAM_mem[4][13] ), .B(\DRAM_mem[20][13] ), .S(n150), .Z(
        n592) );
  MUX2_X1 U640 ( .A(n592), .B(n591), .S(n123), .Z(n593) );
  MUX2_X1 U641 ( .A(\DRAM_mem[8][13] ), .B(\DRAM_mem[24][13] ), .S(n150), .Z(
        n594) );
  MUX2_X1 U642 ( .A(\DRAM_mem[0][13] ), .B(\DRAM_mem[16][13] ), .S(n150), .Z(
        n595) );
  MUX2_X1 U643 ( .A(n595), .B(n594), .S(n123), .Z(n596) );
  MUX2_X1 U644 ( .A(n596), .B(n593), .S(n106), .Z(n597) );
  MUX2_X1 U645 ( .A(n597), .B(n590), .S(Addr[0]), .Z(n598) );
  MUX2_X1 U646 ( .A(n598), .B(n583), .S(Addr[1]), .Z(N486) );
  MUX2_X1 U647 ( .A(\DRAM_mem[15][14] ), .B(\DRAM_mem[31][14] ), .S(n150), .Z(
        n599) );
  MUX2_X1 U648 ( .A(\DRAM_mem[7][14] ), .B(\DRAM_mem[23][14] ), .S(n150), .Z(
        n600) );
  MUX2_X1 U649 ( .A(n600), .B(n599), .S(n123), .Z(n601) );
  MUX2_X1 U650 ( .A(\DRAM_mem[11][14] ), .B(\DRAM_mem[27][14] ), .S(n150), .Z(
        n602) );
  MUX2_X1 U651 ( .A(\DRAM_mem[3][14] ), .B(\DRAM_mem[19][14] ), .S(n150), .Z(
        n603) );
  MUX2_X1 U652 ( .A(n603), .B(n602), .S(n123), .Z(n604) );
  MUX2_X1 U653 ( .A(n604), .B(n601), .S(n106), .Z(n605) );
  MUX2_X1 U654 ( .A(\DRAM_mem[14][14] ), .B(\DRAM_mem[30][14] ), .S(n151), .Z(
        n606) );
  MUX2_X1 U655 ( .A(\DRAM_mem[6][14] ), .B(\DRAM_mem[22][14] ), .S(n151), .Z(
        n607) );
  MUX2_X1 U656 ( .A(n607), .B(n606), .S(n123), .Z(n608) );
  MUX2_X1 U657 ( .A(\DRAM_mem[10][14] ), .B(\DRAM_mem[26][14] ), .S(n151), .Z(
        n609) );
  MUX2_X1 U658 ( .A(\DRAM_mem[2][14] ), .B(\DRAM_mem[18][14] ), .S(n151), .Z(
        n610) );
  MUX2_X1 U659 ( .A(n610), .B(n609), .S(n123), .Z(n611) );
  MUX2_X1 U660 ( .A(n611), .B(n608), .S(n106), .Z(n612) );
  MUX2_X1 U661 ( .A(n612), .B(n605), .S(Addr[0]), .Z(n613) );
  MUX2_X1 U662 ( .A(\DRAM_mem[13][14] ), .B(\DRAM_mem[29][14] ), .S(n151), .Z(
        n614) );
  MUX2_X1 U663 ( .A(\DRAM_mem[5][14] ), .B(\DRAM_mem[21][14] ), .S(n151), .Z(
        n615) );
  MUX2_X1 U664 ( .A(n615), .B(n614), .S(n123), .Z(n616) );
  MUX2_X1 U665 ( .A(\DRAM_mem[9][14] ), .B(\DRAM_mem[25][14] ), .S(n151), .Z(
        n617) );
  MUX2_X1 U666 ( .A(\DRAM_mem[1][14] ), .B(\DRAM_mem[17][14] ), .S(n151), .Z(
        n618) );
  MUX2_X1 U667 ( .A(n618), .B(n617), .S(n123), .Z(n619) );
  MUX2_X1 U668 ( .A(n619), .B(n616), .S(n106), .Z(n620) );
  MUX2_X1 U669 ( .A(\DRAM_mem[12][14] ), .B(\DRAM_mem[28][14] ), .S(n151), .Z(
        n621) );
  MUX2_X1 U670 ( .A(\DRAM_mem[4][14] ), .B(\DRAM_mem[20][14] ), .S(n151), .Z(
        n622) );
  MUX2_X1 U671 ( .A(n622), .B(n621), .S(n123), .Z(n623) );
  MUX2_X1 U672 ( .A(\DRAM_mem[8][14] ), .B(\DRAM_mem[24][14] ), .S(n151), .Z(
        n624) );
  MUX2_X1 U673 ( .A(\DRAM_mem[0][14] ), .B(\DRAM_mem[16][14] ), .S(n151), .Z(
        n625) );
  MUX2_X1 U674 ( .A(n625), .B(n624), .S(n123), .Z(n626) );
  MUX2_X1 U675 ( .A(n626), .B(n623), .S(n106), .Z(n627) );
  MUX2_X1 U676 ( .A(n627), .B(n620), .S(Addr[0]), .Z(n628) );
  MUX2_X1 U677 ( .A(n628), .B(n613), .S(Addr[1]), .Z(N485) );
  MUX2_X1 U678 ( .A(\DRAM_mem[15][15] ), .B(\DRAM_mem[31][15] ), .S(n152), .Z(
        n629) );
  MUX2_X1 U679 ( .A(\DRAM_mem[7][15] ), .B(\DRAM_mem[23][15] ), .S(n152), .Z(
        n630) );
  MUX2_X1 U680 ( .A(n630), .B(n629), .S(n124), .Z(n631) );
  MUX2_X1 U681 ( .A(\DRAM_mem[11][15] ), .B(\DRAM_mem[27][15] ), .S(n152), .Z(
        n632) );
  MUX2_X1 U682 ( .A(\DRAM_mem[3][15] ), .B(\DRAM_mem[19][15] ), .S(n152), .Z(
        n633) );
  MUX2_X1 U683 ( .A(n633), .B(n632), .S(n124), .Z(n634) );
  MUX2_X1 U684 ( .A(n634), .B(n631), .S(n107), .Z(n635) );
  MUX2_X1 U685 ( .A(\DRAM_mem[14][15] ), .B(\DRAM_mem[30][15] ), .S(n152), .Z(
        n636) );
  MUX2_X1 U686 ( .A(\DRAM_mem[6][15] ), .B(\DRAM_mem[22][15] ), .S(n152), .Z(
        n637) );
  MUX2_X1 U687 ( .A(n637), .B(n636), .S(n124), .Z(n638) );
  MUX2_X1 U688 ( .A(\DRAM_mem[10][15] ), .B(\DRAM_mem[26][15] ), .S(n152), .Z(
        n639) );
  MUX2_X1 U689 ( .A(\DRAM_mem[2][15] ), .B(\DRAM_mem[18][15] ), .S(n152), .Z(
        n640) );
  MUX2_X1 U690 ( .A(n640), .B(n639), .S(n124), .Z(n641) );
  MUX2_X1 U691 ( .A(n641), .B(n638), .S(n107), .Z(n642) );
  MUX2_X1 U692 ( .A(n642), .B(n635), .S(Addr[0]), .Z(n643) );
  MUX2_X1 U693 ( .A(\DRAM_mem[13][15] ), .B(\DRAM_mem[29][15] ), .S(n152), .Z(
        n644) );
  MUX2_X1 U694 ( .A(\DRAM_mem[5][15] ), .B(\DRAM_mem[21][15] ), .S(n152), .Z(
        n645) );
  MUX2_X1 U695 ( .A(n645), .B(n644), .S(n124), .Z(n646) );
  MUX2_X1 U696 ( .A(\DRAM_mem[9][15] ), .B(\DRAM_mem[25][15] ), .S(n152), .Z(
        n647) );
  MUX2_X1 U697 ( .A(\DRAM_mem[1][15] ), .B(\DRAM_mem[17][15] ), .S(n152), .Z(
        n648) );
  MUX2_X1 U698 ( .A(n648), .B(n647), .S(n124), .Z(n649) );
  MUX2_X1 U699 ( .A(n649), .B(n646), .S(n107), .Z(n650) );
  MUX2_X1 U700 ( .A(\DRAM_mem[12][15] ), .B(\DRAM_mem[28][15] ), .S(n153), .Z(
        n651) );
  MUX2_X1 U701 ( .A(\DRAM_mem[4][15] ), .B(\DRAM_mem[20][15] ), .S(n153), .Z(
        n652) );
  MUX2_X1 U702 ( .A(n652), .B(n651), .S(n124), .Z(n653) );
  MUX2_X1 U703 ( .A(\DRAM_mem[8][15] ), .B(\DRAM_mem[24][15] ), .S(n153), .Z(
        n654) );
  MUX2_X1 U704 ( .A(\DRAM_mem[0][15] ), .B(\DRAM_mem[16][15] ), .S(n153), .Z(
        n655) );
  MUX2_X1 U705 ( .A(n655), .B(n654), .S(n124), .Z(n656) );
  MUX2_X1 U706 ( .A(n656), .B(n653), .S(n107), .Z(n657) );
  MUX2_X1 U707 ( .A(n657), .B(n650), .S(Addr[0]), .Z(n658) );
  MUX2_X1 U708 ( .A(n658), .B(n643), .S(Addr[1]), .Z(N484) );
  MUX2_X1 U709 ( .A(\DRAM_mem[15][16] ), .B(\DRAM_mem[31][16] ), .S(n153), .Z(
        n659) );
  MUX2_X1 U710 ( .A(\DRAM_mem[7][16] ), .B(\DRAM_mem[23][16] ), .S(n153), .Z(
        n660) );
  MUX2_X1 U711 ( .A(n660), .B(n659), .S(n124), .Z(n661) );
  MUX2_X1 U712 ( .A(\DRAM_mem[11][16] ), .B(\DRAM_mem[27][16] ), .S(n153), .Z(
        n662) );
  MUX2_X1 U713 ( .A(\DRAM_mem[3][16] ), .B(\DRAM_mem[19][16] ), .S(n153), .Z(
        n663) );
  MUX2_X1 U714 ( .A(n663), .B(n662), .S(n124), .Z(n664) );
  MUX2_X1 U715 ( .A(n664), .B(n661), .S(n107), .Z(n665) );
  MUX2_X1 U716 ( .A(\DRAM_mem[14][16] ), .B(\DRAM_mem[30][16] ), .S(n153), .Z(
        n666) );
  MUX2_X1 U717 ( .A(\DRAM_mem[6][16] ), .B(\DRAM_mem[22][16] ), .S(n153), .Z(
        n667) );
  MUX2_X1 U718 ( .A(n667), .B(n666), .S(n124), .Z(n668) );
  MUX2_X1 U719 ( .A(\DRAM_mem[10][16] ), .B(\DRAM_mem[26][16] ), .S(n153), .Z(
        n669) );
  MUX2_X1 U720 ( .A(\DRAM_mem[2][16] ), .B(\DRAM_mem[18][16] ), .S(n153), .Z(
        n670) );
  MUX2_X1 U721 ( .A(n670), .B(n669), .S(n124), .Z(n671) );
  MUX2_X1 U722 ( .A(n671), .B(n668), .S(n107), .Z(n672) );
  MUX2_X1 U723 ( .A(n672), .B(n665), .S(Addr[0]), .Z(n673) );
  MUX2_X1 U724 ( .A(\DRAM_mem[13][16] ), .B(\DRAM_mem[29][16] ), .S(n154), .Z(
        n674) );
  MUX2_X1 U725 ( .A(\DRAM_mem[5][16] ), .B(\DRAM_mem[21][16] ), .S(n154), .Z(
        n675) );
  MUX2_X1 U726 ( .A(n675), .B(n674), .S(n125), .Z(n676) );
  MUX2_X1 U727 ( .A(\DRAM_mem[9][16] ), .B(\DRAM_mem[25][16] ), .S(n154), .Z(
        n677) );
  MUX2_X1 U728 ( .A(\DRAM_mem[1][16] ), .B(\DRAM_mem[17][16] ), .S(n154), .Z(
        n678) );
  MUX2_X1 U729 ( .A(n678), .B(n677), .S(n125), .Z(n679) );
  MUX2_X1 U730 ( .A(n679), .B(n676), .S(n107), .Z(n680) );
  MUX2_X1 U731 ( .A(\DRAM_mem[12][16] ), .B(\DRAM_mem[28][16] ), .S(n154), .Z(
        n681) );
  MUX2_X1 U732 ( .A(\DRAM_mem[4][16] ), .B(\DRAM_mem[20][16] ), .S(n154), .Z(
        n682) );
  MUX2_X1 U733 ( .A(n682), .B(n681), .S(n125), .Z(n683) );
  MUX2_X1 U734 ( .A(\DRAM_mem[8][16] ), .B(\DRAM_mem[24][16] ), .S(n154), .Z(
        n684) );
  MUX2_X1 U735 ( .A(\DRAM_mem[0][16] ), .B(\DRAM_mem[16][16] ), .S(n154), .Z(
        n685) );
  MUX2_X1 U736 ( .A(n685), .B(n684), .S(n125), .Z(n686) );
  MUX2_X1 U737 ( .A(n686), .B(n683), .S(n107), .Z(n687) );
  MUX2_X1 U738 ( .A(n687), .B(n680), .S(Addr[0]), .Z(n688) );
  MUX2_X1 U739 ( .A(n688), .B(n673), .S(Addr[1]), .Z(N401) );
  MUX2_X1 U740 ( .A(\DRAM_mem[15][17] ), .B(\DRAM_mem[31][17] ), .S(n154), .Z(
        n689) );
  MUX2_X1 U741 ( .A(\DRAM_mem[7][17] ), .B(\DRAM_mem[23][17] ), .S(n154), .Z(
        n690) );
  MUX2_X1 U742 ( .A(n690), .B(n689), .S(n125), .Z(n691) );
  MUX2_X1 U743 ( .A(\DRAM_mem[11][17] ), .B(\DRAM_mem[27][17] ), .S(n154), .Z(
        n692) );
  MUX2_X1 U744 ( .A(\DRAM_mem[3][17] ), .B(\DRAM_mem[19][17] ), .S(n154), .Z(
        n693) );
  MUX2_X1 U745 ( .A(n693), .B(n692), .S(n125), .Z(n694) );
  MUX2_X1 U746 ( .A(n694), .B(n691), .S(n107), .Z(n695) );
  MUX2_X1 U747 ( .A(\DRAM_mem[14][17] ), .B(\DRAM_mem[30][17] ), .S(n155), .Z(
        n696) );
  MUX2_X1 U748 ( .A(\DRAM_mem[6][17] ), .B(\DRAM_mem[22][17] ), .S(n155), .Z(
        n697) );
  MUX2_X1 U749 ( .A(n697), .B(n696), .S(n125), .Z(n698) );
  MUX2_X1 U750 ( .A(\DRAM_mem[10][17] ), .B(\DRAM_mem[26][17] ), .S(n155), .Z(
        n699) );
  MUX2_X1 U751 ( .A(\DRAM_mem[2][17] ), .B(\DRAM_mem[18][17] ), .S(n155), .Z(
        n700) );
  MUX2_X1 U752 ( .A(n700), .B(n699), .S(n125), .Z(n701) );
  MUX2_X1 U753 ( .A(n701), .B(n698), .S(n107), .Z(n702) );
  MUX2_X1 U754 ( .A(n702), .B(n695), .S(Addr[0]), .Z(n703) );
  MUX2_X1 U755 ( .A(\DRAM_mem[13][17] ), .B(\DRAM_mem[29][17] ), .S(n155), .Z(
        n704) );
  MUX2_X1 U756 ( .A(\DRAM_mem[5][17] ), .B(\DRAM_mem[21][17] ), .S(n155), .Z(
        n705) );
  MUX2_X1 U757 ( .A(n705), .B(n704), .S(n125), .Z(n706) );
  MUX2_X1 U758 ( .A(\DRAM_mem[9][17] ), .B(\DRAM_mem[25][17] ), .S(n155), .Z(
        n707) );
  MUX2_X1 U759 ( .A(\DRAM_mem[1][17] ), .B(\DRAM_mem[17][17] ), .S(n155), .Z(
        n708) );
  MUX2_X1 U760 ( .A(n708), .B(n707), .S(n125), .Z(n709) );
  MUX2_X1 U761 ( .A(n709), .B(n706), .S(n107), .Z(n710) );
  MUX2_X1 U762 ( .A(\DRAM_mem[12][17] ), .B(\DRAM_mem[28][17] ), .S(n155), .Z(
        n711) );
  MUX2_X1 U763 ( .A(\DRAM_mem[4][17] ), .B(\DRAM_mem[20][17] ), .S(n155), .Z(
        n712) );
  MUX2_X1 U764 ( .A(n712), .B(n711), .S(n125), .Z(n713) );
  MUX2_X1 U765 ( .A(\DRAM_mem[8][17] ), .B(\DRAM_mem[24][17] ), .S(n155), .Z(
        n714) );
  MUX2_X1 U766 ( .A(\DRAM_mem[0][17] ), .B(\DRAM_mem[16][17] ), .S(n155), .Z(
        n715) );
  MUX2_X1 U767 ( .A(n715), .B(n714), .S(n125), .Z(n716) );
  MUX2_X1 U768 ( .A(n716), .B(n713), .S(n107), .Z(n717) );
  MUX2_X1 U769 ( .A(n717), .B(n710), .S(Addr[0]), .Z(n718) );
  MUX2_X1 U770 ( .A(n718), .B(n703), .S(Addr[1]), .Z(N400) );
  MUX2_X1 U771 ( .A(\DRAM_mem[15][18] ), .B(\DRAM_mem[31][18] ), .S(n156), .Z(
        n719) );
  MUX2_X1 U772 ( .A(\DRAM_mem[7][18] ), .B(\DRAM_mem[23][18] ), .S(n156), .Z(
        n720) );
  MUX2_X1 U773 ( .A(n720), .B(n719), .S(n126), .Z(n721) );
  MUX2_X1 U774 ( .A(\DRAM_mem[11][18] ), .B(\DRAM_mem[27][18] ), .S(n156), .Z(
        n722) );
  MUX2_X1 U775 ( .A(\DRAM_mem[3][18] ), .B(\DRAM_mem[19][18] ), .S(n156), .Z(
        n723) );
  MUX2_X1 U776 ( .A(n723), .B(n722), .S(n126), .Z(n724) );
  MUX2_X1 U777 ( .A(n724), .B(n721), .S(n108), .Z(n725) );
  MUX2_X1 U778 ( .A(\DRAM_mem[14][18] ), .B(\DRAM_mem[30][18] ), .S(n156), .Z(
        n726) );
  MUX2_X1 U779 ( .A(\DRAM_mem[6][18] ), .B(\DRAM_mem[22][18] ), .S(n156), .Z(
        n727) );
  MUX2_X1 U780 ( .A(n727), .B(n726), .S(n126), .Z(n728) );
  MUX2_X1 U781 ( .A(\DRAM_mem[10][18] ), .B(\DRAM_mem[26][18] ), .S(n156), .Z(
        n729) );
  MUX2_X1 U782 ( .A(\DRAM_mem[2][18] ), .B(\DRAM_mem[18][18] ), .S(n156), .Z(
        n730) );
  MUX2_X1 U783 ( .A(n730), .B(n729), .S(n126), .Z(n731) );
  MUX2_X1 U784 ( .A(n731), .B(n728), .S(n108), .Z(n732) );
  MUX2_X1 U785 ( .A(n732), .B(n725), .S(Addr[0]), .Z(n733) );
  MUX2_X1 U786 ( .A(\DRAM_mem[13][18] ), .B(\DRAM_mem[29][18] ), .S(n156), .Z(
        n734) );
  MUX2_X1 U787 ( .A(\DRAM_mem[5][18] ), .B(\DRAM_mem[21][18] ), .S(n156), .Z(
        n735) );
  MUX2_X1 U788 ( .A(n735), .B(n734), .S(n126), .Z(n736) );
  MUX2_X1 U789 ( .A(\DRAM_mem[9][18] ), .B(\DRAM_mem[25][18] ), .S(n156), .Z(
        n737) );
  MUX2_X1 U790 ( .A(\DRAM_mem[1][18] ), .B(\DRAM_mem[17][18] ), .S(n156), .Z(
        n738) );
  MUX2_X1 U791 ( .A(n738), .B(n737), .S(n126), .Z(n739) );
  MUX2_X1 U792 ( .A(n739), .B(n736), .S(n108), .Z(n740) );
  MUX2_X1 U793 ( .A(\DRAM_mem[12][18] ), .B(\DRAM_mem[28][18] ), .S(n157), .Z(
        n741) );
  MUX2_X1 U794 ( .A(\DRAM_mem[4][18] ), .B(\DRAM_mem[20][18] ), .S(n157), .Z(
        n742) );
  MUX2_X1 U795 ( .A(n742), .B(n741), .S(n126), .Z(n743) );
  MUX2_X1 U796 ( .A(\DRAM_mem[8][18] ), .B(\DRAM_mem[24][18] ), .S(n157), .Z(
        n744) );
  MUX2_X1 U797 ( .A(\DRAM_mem[0][18] ), .B(\DRAM_mem[16][18] ), .S(n157), .Z(
        n745) );
  MUX2_X1 U798 ( .A(n745), .B(n744), .S(n126), .Z(n746) );
  MUX2_X1 U799 ( .A(n746), .B(n743), .S(n108), .Z(n747) );
  MUX2_X1 U800 ( .A(n747), .B(n740), .S(Addr[0]), .Z(n748) );
  MUX2_X1 U801 ( .A(n748), .B(n733), .S(Addr[1]), .Z(N399) );
  MUX2_X1 U802 ( .A(\DRAM_mem[15][19] ), .B(\DRAM_mem[31][19] ), .S(n157), .Z(
        n749) );
  MUX2_X1 U803 ( .A(\DRAM_mem[7][19] ), .B(\DRAM_mem[23][19] ), .S(n157), .Z(
        n750) );
  MUX2_X1 U804 ( .A(n750), .B(n749), .S(n126), .Z(n751) );
  MUX2_X1 U805 ( .A(\DRAM_mem[11][19] ), .B(\DRAM_mem[27][19] ), .S(n157), .Z(
        n752) );
  MUX2_X1 U806 ( .A(\DRAM_mem[3][19] ), .B(\DRAM_mem[19][19] ), .S(n157), .Z(
        n753) );
  MUX2_X1 U807 ( .A(n753), .B(n752), .S(n126), .Z(n754) );
  MUX2_X1 U808 ( .A(n754), .B(n751), .S(n108), .Z(n755) );
  MUX2_X1 U809 ( .A(\DRAM_mem[14][19] ), .B(\DRAM_mem[30][19] ), .S(n157), .Z(
        n756) );
  MUX2_X1 U810 ( .A(\DRAM_mem[6][19] ), .B(\DRAM_mem[22][19] ), .S(n157), .Z(
        n757) );
  MUX2_X1 U811 ( .A(n757), .B(n756), .S(n126), .Z(n758) );
  MUX2_X1 U812 ( .A(\DRAM_mem[10][19] ), .B(\DRAM_mem[26][19] ), .S(n157), .Z(
        n759) );
  MUX2_X1 U813 ( .A(\DRAM_mem[2][19] ), .B(\DRAM_mem[18][19] ), .S(n157), .Z(
        n760) );
  MUX2_X1 U814 ( .A(n760), .B(n759), .S(n126), .Z(n761) );
  MUX2_X1 U815 ( .A(n761), .B(n758), .S(n108), .Z(n762) );
  MUX2_X1 U816 ( .A(n762), .B(n755), .S(Addr[0]), .Z(n763) );
  MUX2_X1 U817 ( .A(\DRAM_mem[13][19] ), .B(\DRAM_mem[29][19] ), .S(n158), .Z(
        n764) );
  MUX2_X1 U818 ( .A(\DRAM_mem[5][19] ), .B(\DRAM_mem[21][19] ), .S(n158), .Z(
        n765) );
  MUX2_X1 U819 ( .A(n765), .B(n764), .S(n127), .Z(n766) );
  MUX2_X1 U820 ( .A(\DRAM_mem[9][19] ), .B(\DRAM_mem[25][19] ), .S(n158), .Z(
        n767) );
  MUX2_X1 U821 ( .A(\DRAM_mem[1][19] ), .B(\DRAM_mem[17][19] ), .S(n158), .Z(
        n768) );
  MUX2_X1 U822 ( .A(n768), .B(n767), .S(n127), .Z(n769) );
  MUX2_X1 U823 ( .A(n769), .B(n766), .S(n108), .Z(n770) );
  MUX2_X1 U824 ( .A(\DRAM_mem[12][19] ), .B(\DRAM_mem[28][19] ), .S(n158), .Z(
        n771) );
  MUX2_X1 U825 ( .A(\DRAM_mem[4][19] ), .B(\DRAM_mem[20][19] ), .S(n158), .Z(
        n772) );
  MUX2_X1 U826 ( .A(n772), .B(n771), .S(n127), .Z(n773) );
  MUX2_X1 U827 ( .A(\DRAM_mem[8][19] ), .B(\DRAM_mem[24][19] ), .S(n158), .Z(
        n774) );
  MUX2_X1 U828 ( .A(\DRAM_mem[0][19] ), .B(\DRAM_mem[16][19] ), .S(n158), .Z(
        n775) );
  MUX2_X1 U829 ( .A(n775), .B(n774), .S(n127), .Z(n776) );
  MUX2_X1 U830 ( .A(n776), .B(n773), .S(n108), .Z(n777) );
  MUX2_X1 U831 ( .A(n777), .B(n770), .S(Addr[0]), .Z(n778) );
  MUX2_X1 U832 ( .A(n778), .B(n763), .S(Addr[1]), .Z(N398) );
  MUX2_X1 U833 ( .A(\DRAM_mem[15][20] ), .B(\DRAM_mem[31][20] ), .S(n158), .Z(
        n779) );
  MUX2_X1 U834 ( .A(\DRAM_mem[7][20] ), .B(\DRAM_mem[23][20] ), .S(n158), .Z(
        n780) );
  MUX2_X1 U835 ( .A(n780), .B(n779), .S(n127), .Z(n781) );
  MUX2_X1 U836 ( .A(\DRAM_mem[11][20] ), .B(\DRAM_mem[27][20] ), .S(n158), .Z(
        n782) );
  MUX2_X1 U837 ( .A(\DRAM_mem[3][20] ), .B(\DRAM_mem[19][20] ), .S(n158), .Z(
        n783) );
  MUX2_X1 U838 ( .A(n783), .B(n782), .S(n127), .Z(n784) );
  MUX2_X1 U839 ( .A(n784), .B(n781), .S(n108), .Z(n785) );
  MUX2_X1 U840 ( .A(\DRAM_mem[14][20] ), .B(\DRAM_mem[30][20] ), .S(n159), .Z(
        n786) );
  MUX2_X1 U841 ( .A(\DRAM_mem[6][20] ), .B(\DRAM_mem[22][20] ), .S(n159), .Z(
        n787) );
  MUX2_X1 U842 ( .A(n787), .B(n786), .S(n127), .Z(n788) );
  MUX2_X1 U843 ( .A(\DRAM_mem[10][20] ), .B(\DRAM_mem[26][20] ), .S(n159), .Z(
        n789) );
  MUX2_X1 U844 ( .A(\DRAM_mem[2][20] ), .B(\DRAM_mem[18][20] ), .S(n159), .Z(
        n790) );
  MUX2_X1 U845 ( .A(n790), .B(n789), .S(n127), .Z(n791) );
  MUX2_X1 U846 ( .A(n791), .B(n788), .S(n108), .Z(n792) );
  MUX2_X1 U847 ( .A(n792), .B(n785), .S(Addr[0]), .Z(n793) );
  MUX2_X1 U848 ( .A(\DRAM_mem[13][20] ), .B(\DRAM_mem[29][20] ), .S(n159), .Z(
        n794) );
  MUX2_X1 U849 ( .A(\DRAM_mem[5][20] ), .B(\DRAM_mem[21][20] ), .S(n159), .Z(
        n795) );
  MUX2_X1 U850 ( .A(n795), .B(n794), .S(n127), .Z(n796) );
  MUX2_X1 U851 ( .A(\DRAM_mem[9][20] ), .B(\DRAM_mem[25][20] ), .S(n159), .Z(
        n797) );
  MUX2_X1 U852 ( .A(\DRAM_mem[1][20] ), .B(\DRAM_mem[17][20] ), .S(n159), .Z(
        n798) );
  MUX2_X1 U853 ( .A(n798), .B(n797), .S(n127), .Z(n799) );
  MUX2_X1 U854 ( .A(n799), .B(n796), .S(n108), .Z(n800) );
  MUX2_X1 U855 ( .A(\DRAM_mem[12][20] ), .B(\DRAM_mem[28][20] ), .S(n159), .Z(
        n801) );
  MUX2_X1 U856 ( .A(\DRAM_mem[4][20] ), .B(\DRAM_mem[20][20] ), .S(n159), .Z(
        n802) );
  MUX2_X1 U857 ( .A(n802), .B(n801), .S(n127), .Z(n803) );
  MUX2_X1 U858 ( .A(\DRAM_mem[8][20] ), .B(\DRAM_mem[24][20] ), .S(n159), .Z(
        n804) );
  MUX2_X1 U859 ( .A(\DRAM_mem[0][20] ), .B(\DRAM_mem[16][20] ), .S(n159), .Z(
        n805) );
  MUX2_X1 U860 ( .A(n805), .B(n804), .S(n127), .Z(n806) );
  MUX2_X1 U861 ( .A(n806), .B(n803), .S(n108), .Z(n807) );
  MUX2_X1 U862 ( .A(n807), .B(n800), .S(Addr[0]), .Z(n808) );
  MUX2_X1 U863 ( .A(n808), .B(n793), .S(Addr[1]), .Z(N397) );
  MUX2_X1 U864 ( .A(\DRAM_mem[15][21] ), .B(\DRAM_mem[31][21] ), .S(n160), .Z(
        n809) );
  MUX2_X1 U865 ( .A(\DRAM_mem[7][21] ), .B(\DRAM_mem[23][21] ), .S(n160), .Z(
        n810) );
  MUX2_X1 U866 ( .A(n810), .B(n809), .S(n128), .Z(n811) );
  MUX2_X1 U867 ( .A(\DRAM_mem[11][21] ), .B(\DRAM_mem[27][21] ), .S(n160), .Z(
        n812) );
  MUX2_X1 U868 ( .A(\DRAM_mem[3][21] ), .B(\DRAM_mem[19][21] ), .S(n160), .Z(
        n813) );
  MUX2_X1 U869 ( .A(n813), .B(n812), .S(n128), .Z(n814) );
  MUX2_X1 U870 ( .A(n814), .B(n811), .S(n109), .Z(n815) );
  MUX2_X1 U871 ( .A(\DRAM_mem[14][21] ), .B(\DRAM_mem[30][21] ), .S(n160), .Z(
        n816) );
  MUX2_X1 U872 ( .A(\DRAM_mem[6][21] ), .B(\DRAM_mem[22][21] ), .S(n160), .Z(
        n817) );
  MUX2_X1 U873 ( .A(n817), .B(n816), .S(n128), .Z(n818) );
  MUX2_X1 U874 ( .A(\DRAM_mem[10][21] ), .B(\DRAM_mem[26][21] ), .S(n160), .Z(
        n819) );
  MUX2_X1 U875 ( .A(\DRAM_mem[2][21] ), .B(\DRAM_mem[18][21] ), .S(n160), .Z(
        n820) );
  MUX2_X1 U876 ( .A(n820), .B(n819), .S(n128), .Z(n821) );
  MUX2_X1 U877 ( .A(n821), .B(n818), .S(n109), .Z(n822) );
  MUX2_X1 U878 ( .A(n822), .B(n815), .S(Addr[0]), .Z(n823) );
  MUX2_X1 U879 ( .A(\DRAM_mem[13][21] ), .B(\DRAM_mem[29][21] ), .S(n160), .Z(
        n824) );
  MUX2_X1 U880 ( .A(\DRAM_mem[5][21] ), .B(\DRAM_mem[21][21] ), .S(n160), .Z(
        n825) );
  MUX2_X1 U881 ( .A(n825), .B(n824), .S(n128), .Z(n826) );
  MUX2_X1 U882 ( .A(\DRAM_mem[9][21] ), .B(\DRAM_mem[25][21] ), .S(n160), .Z(
        n827) );
  MUX2_X1 U883 ( .A(\DRAM_mem[1][21] ), .B(\DRAM_mem[17][21] ), .S(n160), .Z(
        n828) );
  MUX2_X1 U884 ( .A(n828), .B(n827), .S(n128), .Z(n829) );
  MUX2_X1 U885 ( .A(n829), .B(n826), .S(n109), .Z(n830) );
  MUX2_X1 U886 ( .A(\DRAM_mem[12][21] ), .B(\DRAM_mem[28][21] ), .S(n161), .Z(
        n831) );
  MUX2_X1 U887 ( .A(\DRAM_mem[4][21] ), .B(\DRAM_mem[20][21] ), .S(n161), .Z(
        n832) );
  MUX2_X1 U888 ( .A(n832), .B(n831), .S(n128), .Z(n833) );
  MUX2_X1 U889 ( .A(\DRAM_mem[8][21] ), .B(\DRAM_mem[24][21] ), .S(n161), .Z(
        n834) );
  MUX2_X1 U890 ( .A(\DRAM_mem[0][21] ), .B(\DRAM_mem[16][21] ), .S(n161), .Z(
        n835) );
  MUX2_X1 U891 ( .A(n835), .B(n834), .S(n128), .Z(n836) );
  MUX2_X1 U892 ( .A(n836), .B(n833), .S(n109), .Z(n837) );
  MUX2_X1 U893 ( .A(n837), .B(n830), .S(Addr[0]), .Z(n838) );
  MUX2_X1 U894 ( .A(n838), .B(n823), .S(Addr[1]), .Z(N396) );
  MUX2_X1 U895 ( .A(\DRAM_mem[15][22] ), .B(\DRAM_mem[31][22] ), .S(n161), .Z(
        n839) );
  MUX2_X1 U896 ( .A(\DRAM_mem[7][22] ), .B(\DRAM_mem[23][22] ), .S(n161), .Z(
        n840) );
  MUX2_X1 U897 ( .A(n840), .B(n839), .S(n128), .Z(n841) );
  MUX2_X1 U898 ( .A(\DRAM_mem[11][22] ), .B(\DRAM_mem[27][22] ), .S(n161), .Z(
        n842) );
  MUX2_X1 U899 ( .A(\DRAM_mem[3][22] ), .B(\DRAM_mem[19][22] ), .S(n161), .Z(
        n843) );
  MUX2_X1 U900 ( .A(n843), .B(n842), .S(n128), .Z(n844) );
  MUX2_X1 U901 ( .A(n844), .B(n841), .S(n109), .Z(n845) );
  MUX2_X1 U902 ( .A(\DRAM_mem[14][22] ), .B(\DRAM_mem[30][22] ), .S(n161), .Z(
        n846) );
  MUX2_X1 U903 ( .A(\DRAM_mem[6][22] ), .B(\DRAM_mem[22][22] ), .S(n161), .Z(
        n847) );
  MUX2_X1 U904 ( .A(n847), .B(n846), .S(n128), .Z(n848) );
  MUX2_X1 U905 ( .A(\DRAM_mem[10][22] ), .B(\DRAM_mem[26][22] ), .S(n161), .Z(
        n849) );
  MUX2_X1 U906 ( .A(\DRAM_mem[2][22] ), .B(\DRAM_mem[18][22] ), .S(n161), .Z(
        n850) );
  MUX2_X1 U907 ( .A(n850), .B(n849), .S(n128), .Z(n851) );
  MUX2_X1 U908 ( .A(n851), .B(n848), .S(n109), .Z(n852) );
  MUX2_X1 U909 ( .A(n852), .B(n845), .S(Addr[0]), .Z(n853) );
  MUX2_X1 U910 ( .A(\DRAM_mem[13][22] ), .B(\DRAM_mem[29][22] ), .S(n162), .Z(
        n854) );
  MUX2_X1 U911 ( .A(\DRAM_mem[5][22] ), .B(\DRAM_mem[21][22] ), .S(n162), .Z(
        n855) );
  MUX2_X1 U912 ( .A(n855), .B(n854), .S(n129), .Z(n856) );
  MUX2_X1 U913 ( .A(\DRAM_mem[9][22] ), .B(\DRAM_mem[25][22] ), .S(n162), .Z(
        n857) );
  MUX2_X1 U914 ( .A(\DRAM_mem[1][22] ), .B(\DRAM_mem[17][22] ), .S(n162), .Z(
        n858) );
  MUX2_X1 U915 ( .A(n858), .B(n857), .S(n129), .Z(n859) );
  MUX2_X1 U916 ( .A(n859), .B(n856), .S(n109), .Z(n860) );
  MUX2_X1 U917 ( .A(\DRAM_mem[12][22] ), .B(\DRAM_mem[28][22] ), .S(n162), .Z(
        n861) );
  MUX2_X1 U918 ( .A(\DRAM_mem[4][22] ), .B(\DRAM_mem[20][22] ), .S(n162), .Z(
        n862) );
  MUX2_X1 U919 ( .A(n862), .B(n861), .S(n129), .Z(n863) );
  MUX2_X1 U920 ( .A(\DRAM_mem[8][22] ), .B(\DRAM_mem[24][22] ), .S(n162), .Z(
        n864) );
  MUX2_X1 U921 ( .A(\DRAM_mem[0][22] ), .B(\DRAM_mem[16][22] ), .S(n162), .Z(
        n865) );
  MUX2_X1 U922 ( .A(n865), .B(n864), .S(n129), .Z(n866) );
  MUX2_X1 U923 ( .A(n866), .B(n863), .S(n109), .Z(n867) );
  MUX2_X1 U924 ( .A(n867), .B(n860), .S(Addr[0]), .Z(n868) );
  MUX2_X1 U925 ( .A(n868), .B(n853), .S(Addr[1]), .Z(N395) );
  MUX2_X1 U926 ( .A(\DRAM_mem[15][23] ), .B(\DRAM_mem[31][23] ), .S(n162), .Z(
        n869) );
  MUX2_X1 U927 ( .A(\DRAM_mem[7][23] ), .B(\DRAM_mem[23][23] ), .S(n162), .Z(
        n870) );
  MUX2_X1 U928 ( .A(n870), .B(n869), .S(n129), .Z(n871) );
  MUX2_X1 U929 ( .A(\DRAM_mem[11][23] ), .B(\DRAM_mem[27][23] ), .S(n162), .Z(
        n872) );
  MUX2_X1 U930 ( .A(\DRAM_mem[3][23] ), .B(\DRAM_mem[19][23] ), .S(n162), .Z(
        n873) );
  MUX2_X1 U931 ( .A(n873), .B(n872), .S(n129), .Z(n874) );
  MUX2_X1 U932 ( .A(n874), .B(n871), .S(n109), .Z(n875) );
  MUX2_X1 U933 ( .A(\DRAM_mem[14][23] ), .B(\DRAM_mem[30][23] ), .S(n163), .Z(
        n876) );
  MUX2_X1 U934 ( .A(\DRAM_mem[6][23] ), .B(\DRAM_mem[22][23] ), .S(n163), .Z(
        n877) );
  MUX2_X1 U935 ( .A(n877), .B(n876), .S(n129), .Z(n878) );
  MUX2_X1 U936 ( .A(\DRAM_mem[10][23] ), .B(\DRAM_mem[26][23] ), .S(n163), .Z(
        n879) );
  MUX2_X1 U937 ( .A(\DRAM_mem[2][23] ), .B(\DRAM_mem[18][23] ), .S(n163), .Z(
        n880) );
  MUX2_X1 U938 ( .A(n880), .B(n879), .S(n129), .Z(n881) );
  MUX2_X1 U939 ( .A(n881), .B(n878), .S(n109), .Z(n882) );
  MUX2_X1 U940 ( .A(n882), .B(n875), .S(Addr[0]), .Z(n883) );
  MUX2_X1 U941 ( .A(\DRAM_mem[13][23] ), .B(\DRAM_mem[29][23] ), .S(n163), .Z(
        n884) );
  MUX2_X1 U942 ( .A(\DRAM_mem[5][23] ), .B(\DRAM_mem[21][23] ), .S(n163), .Z(
        n885) );
  MUX2_X1 U943 ( .A(n885), .B(n884), .S(n129), .Z(n886) );
  MUX2_X1 U944 ( .A(\DRAM_mem[9][23] ), .B(\DRAM_mem[25][23] ), .S(n163), .Z(
        n887) );
  MUX2_X1 U945 ( .A(\DRAM_mem[1][23] ), .B(\DRAM_mem[17][23] ), .S(n163), .Z(
        n888) );
  MUX2_X1 U946 ( .A(n888), .B(n887), .S(n129), .Z(n889) );
  MUX2_X1 U947 ( .A(n889), .B(n886), .S(n109), .Z(n890) );
  MUX2_X1 U948 ( .A(\DRAM_mem[12][23] ), .B(\DRAM_mem[28][23] ), .S(n163), .Z(
        n891) );
  MUX2_X1 U949 ( .A(\DRAM_mem[4][23] ), .B(\DRAM_mem[20][23] ), .S(n163), .Z(
        n892) );
  MUX2_X1 U950 ( .A(n892), .B(n891), .S(n129), .Z(n893) );
  MUX2_X1 U951 ( .A(\DRAM_mem[8][23] ), .B(\DRAM_mem[24][23] ), .S(n163), .Z(
        n894) );
  MUX2_X1 U952 ( .A(\DRAM_mem[0][23] ), .B(\DRAM_mem[16][23] ), .S(n163), .Z(
        n895) );
  MUX2_X1 U953 ( .A(n895), .B(n894), .S(n129), .Z(n896) );
  MUX2_X1 U954 ( .A(n896), .B(n893), .S(n109), .Z(n897) );
  MUX2_X1 U955 ( .A(n897), .B(n890), .S(Addr[0]), .Z(n898) );
  MUX2_X1 U956 ( .A(n898), .B(n883), .S(Addr[1]), .Z(N394) );
  MUX2_X1 U957 ( .A(\DRAM_mem[15][24] ), .B(\DRAM_mem[31][24] ), .S(n164), .Z(
        n899) );
  MUX2_X1 U958 ( .A(\DRAM_mem[7][24] ), .B(\DRAM_mem[23][24] ), .S(n164), .Z(
        n900) );
  MUX2_X1 U959 ( .A(n900), .B(n899), .S(n130), .Z(n901) );
  MUX2_X1 U960 ( .A(\DRAM_mem[11][24] ), .B(\DRAM_mem[27][24] ), .S(n164), .Z(
        n902) );
  MUX2_X1 U961 ( .A(\DRAM_mem[3][24] ), .B(\DRAM_mem[19][24] ), .S(n164), .Z(
        n903) );
  MUX2_X1 U962 ( .A(n903), .B(n902), .S(n130), .Z(n904) );
  MUX2_X1 U963 ( .A(n904), .B(n901), .S(n110), .Z(n905) );
  MUX2_X1 U964 ( .A(\DRAM_mem[14][24] ), .B(\DRAM_mem[30][24] ), .S(n164), .Z(
        n906) );
  MUX2_X1 U965 ( .A(\DRAM_mem[6][24] ), .B(\DRAM_mem[22][24] ), .S(n164), .Z(
        n907) );
  MUX2_X1 U966 ( .A(n907), .B(n906), .S(n130), .Z(n908) );
  MUX2_X1 U967 ( .A(\DRAM_mem[10][24] ), .B(\DRAM_mem[26][24] ), .S(n164), .Z(
        n909) );
  MUX2_X1 U968 ( .A(\DRAM_mem[2][24] ), .B(\DRAM_mem[18][24] ), .S(n164), .Z(
        n910) );
  MUX2_X1 U969 ( .A(n910), .B(n909), .S(n130), .Z(n911) );
  MUX2_X1 U970 ( .A(n911), .B(n908), .S(n110), .Z(n912) );
  MUX2_X1 U971 ( .A(n912), .B(n905), .S(Addr[0]), .Z(n913) );
  MUX2_X1 U972 ( .A(\DRAM_mem[13][24] ), .B(\DRAM_mem[29][24] ), .S(n164), .Z(
        n914) );
  MUX2_X1 U973 ( .A(\DRAM_mem[5][24] ), .B(\DRAM_mem[21][24] ), .S(n164), .Z(
        n915) );
  MUX2_X1 U974 ( .A(n915), .B(n914), .S(n130), .Z(n916) );
  MUX2_X1 U975 ( .A(\DRAM_mem[9][24] ), .B(\DRAM_mem[25][24] ), .S(n164), .Z(
        n917) );
  MUX2_X1 U976 ( .A(\DRAM_mem[1][24] ), .B(\DRAM_mem[17][24] ), .S(n164), .Z(
        n918) );
  MUX2_X1 U977 ( .A(n918), .B(n917), .S(n130), .Z(n919) );
  MUX2_X1 U978 ( .A(n919), .B(n916), .S(n110), .Z(n920) );
  MUX2_X1 U979 ( .A(\DRAM_mem[12][24] ), .B(\DRAM_mem[28][24] ), .S(n165), .Z(
        n921) );
  MUX2_X1 U980 ( .A(\DRAM_mem[4][24] ), .B(\DRAM_mem[20][24] ), .S(n165), .Z(
        n922) );
  MUX2_X1 U981 ( .A(n922), .B(n921), .S(n130), .Z(n923) );
  MUX2_X1 U982 ( .A(\DRAM_mem[8][24] ), .B(\DRAM_mem[24][24] ), .S(n165), .Z(
        n924) );
  MUX2_X1 U983 ( .A(\DRAM_mem[0][24] ), .B(\DRAM_mem[16][24] ), .S(n165), .Z(
        n925) );
  MUX2_X1 U984 ( .A(n925), .B(n924), .S(n130), .Z(n926) );
  MUX2_X1 U985 ( .A(n926), .B(n923), .S(n110), .Z(n927) );
  MUX2_X1 U986 ( .A(n927), .B(n920), .S(Addr[0]), .Z(n928) );
  MUX2_X1 U987 ( .A(n928), .B(n913), .S(Addr[1]), .Z(N393) );
  MUX2_X1 U988 ( .A(\DRAM_mem[15][25] ), .B(\DRAM_mem[31][25] ), .S(n165), .Z(
        n929) );
  MUX2_X1 U989 ( .A(\DRAM_mem[7][25] ), .B(\DRAM_mem[23][25] ), .S(n165), .Z(
        n930) );
  MUX2_X1 U990 ( .A(n930), .B(n929), .S(n130), .Z(n931) );
  MUX2_X1 U991 ( .A(\DRAM_mem[11][25] ), .B(\DRAM_mem[27][25] ), .S(n165), .Z(
        n932) );
  MUX2_X1 U992 ( .A(\DRAM_mem[3][25] ), .B(\DRAM_mem[19][25] ), .S(n165), .Z(
        n933) );
  MUX2_X1 U993 ( .A(n933), .B(n932), .S(n130), .Z(n934) );
  MUX2_X1 U994 ( .A(n934), .B(n931), .S(n110), .Z(n935) );
  MUX2_X1 U995 ( .A(\DRAM_mem[14][25] ), .B(\DRAM_mem[30][25] ), .S(n165), .Z(
        n936) );
  MUX2_X1 U996 ( .A(\DRAM_mem[6][25] ), .B(\DRAM_mem[22][25] ), .S(n165), .Z(
        n937) );
  MUX2_X1 U997 ( .A(n937), .B(n936), .S(n130), .Z(n938) );
  MUX2_X1 U998 ( .A(\DRAM_mem[10][25] ), .B(\DRAM_mem[26][25] ), .S(n165), .Z(
        n939) );
  MUX2_X1 U999 ( .A(\DRAM_mem[2][25] ), .B(\DRAM_mem[18][25] ), .S(n165), .Z(
        n940) );
  MUX2_X1 U1000 ( .A(n940), .B(n939), .S(n130), .Z(n941) );
  MUX2_X1 U1001 ( .A(n941), .B(n938), .S(n110), .Z(n942) );
  MUX2_X1 U1002 ( .A(n942), .B(n935), .S(Addr[0]), .Z(n943) );
  MUX2_X1 U1003 ( .A(\DRAM_mem[13][25] ), .B(\DRAM_mem[29][25] ), .S(n166), 
        .Z(n944) );
  MUX2_X1 U1004 ( .A(\DRAM_mem[5][25] ), .B(\DRAM_mem[21][25] ), .S(n166), .Z(
        n945) );
  MUX2_X1 U1005 ( .A(n945), .B(n944), .S(n131), .Z(n946) );
  MUX2_X1 U1006 ( .A(\DRAM_mem[9][25] ), .B(\DRAM_mem[25][25] ), .S(n166), .Z(
        n947) );
  MUX2_X1 U1007 ( .A(\DRAM_mem[1][25] ), .B(\DRAM_mem[17][25] ), .S(n166), .Z(
        n948) );
  MUX2_X1 U1008 ( .A(n948), .B(n947), .S(n131), .Z(n949) );
  MUX2_X1 U1009 ( .A(n949), .B(n946), .S(n110), .Z(n950) );
  MUX2_X1 U1010 ( .A(\DRAM_mem[12][25] ), .B(\DRAM_mem[28][25] ), .S(n166), 
        .Z(n951) );
  MUX2_X1 U1011 ( .A(\DRAM_mem[4][25] ), .B(\DRAM_mem[20][25] ), .S(n166), .Z(
        n952) );
  MUX2_X1 U1012 ( .A(n952), .B(n951), .S(n131), .Z(n953) );
  MUX2_X1 U1013 ( .A(\DRAM_mem[8][25] ), .B(\DRAM_mem[24][25] ), .S(n166), .Z(
        n954) );
  MUX2_X1 U1014 ( .A(\DRAM_mem[0][25] ), .B(\DRAM_mem[16][25] ), .S(n166), .Z(
        n955) );
  MUX2_X1 U1015 ( .A(n955), .B(n954), .S(n131), .Z(n956) );
  MUX2_X1 U1016 ( .A(n956), .B(n953), .S(n110), .Z(n957) );
  MUX2_X1 U1017 ( .A(n957), .B(n950), .S(Addr[0]), .Z(n958) );
  MUX2_X1 U1018 ( .A(n958), .B(n943), .S(Addr[1]), .Z(N392) );
  MUX2_X1 U1019 ( .A(\DRAM_mem[15][26] ), .B(\DRAM_mem[31][26] ), .S(n166), 
        .Z(n959) );
  MUX2_X1 U1020 ( .A(\DRAM_mem[7][26] ), .B(\DRAM_mem[23][26] ), .S(n166), .Z(
        n960) );
  MUX2_X1 U1021 ( .A(n960), .B(n959), .S(n131), .Z(n961) );
  MUX2_X1 U1022 ( .A(\DRAM_mem[11][26] ), .B(\DRAM_mem[27][26] ), .S(n166), 
        .Z(n962) );
  MUX2_X1 U1023 ( .A(\DRAM_mem[3][26] ), .B(\DRAM_mem[19][26] ), .S(n166), .Z(
        n963) );
  MUX2_X1 U1024 ( .A(n963), .B(n962), .S(n131), .Z(n964) );
  MUX2_X1 U1025 ( .A(n964), .B(n961), .S(n110), .Z(n965) );
  MUX2_X1 U1026 ( .A(\DRAM_mem[14][26] ), .B(\DRAM_mem[30][26] ), .S(n167), 
        .Z(n966) );
  MUX2_X1 U1027 ( .A(\DRAM_mem[6][26] ), .B(\DRAM_mem[22][26] ), .S(n167), .Z(
        n967) );
  MUX2_X1 U1028 ( .A(n967), .B(n966), .S(n131), .Z(n968) );
  MUX2_X1 U1029 ( .A(\DRAM_mem[10][26] ), .B(\DRAM_mem[26][26] ), .S(n167), 
        .Z(n969) );
  MUX2_X1 U1030 ( .A(\DRAM_mem[2][26] ), .B(\DRAM_mem[18][26] ), .S(n167), .Z(
        n970) );
  MUX2_X1 U1031 ( .A(n970), .B(n969), .S(n131), .Z(n971) );
  MUX2_X1 U1032 ( .A(n971), .B(n968), .S(n110), .Z(n972) );
  MUX2_X1 U1033 ( .A(n972), .B(n965), .S(Addr[0]), .Z(n973) );
  MUX2_X1 U1034 ( .A(\DRAM_mem[13][26] ), .B(\DRAM_mem[29][26] ), .S(n167), 
        .Z(n974) );
  MUX2_X1 U1035 ( .A(\DRAM_mem[5][26] ), .B(\DRAM_mem[21][26] ), .S(n167), .Z(
        n975) );
  MUX2_X1 U1036 ( .A(n975), .B(n974), .S(n131), .Z(n976) );
  MUX2_X1 U1037 ( .A(\DRAM_mem[9][26] ), .B(\DRAM_mem[25][26] ), .S(n167), .Z(
        n977) );
  MUX2_X1 U1038 ( .A(\DRAM_mem[1][26] ), .B(\DRAM_mem[17][26] ), .S(n167), .Z(
        n978) );
  MUX2_X1 U1039 ( .A(n978), .B(n977), .S(n131), .Z(n979) );
  MUX2_X1 U1040 ( .A(n979), .B(n976), .S(n110), .Z(n980) );
  MUX2_X1 U1041 ( .A(\DRAM_mem[12][26] ), .B(\DRAM_mem[28][26] ), .S(n167), 
        .Z(n981) );
  MUX2_X1 U1042 ( .A(\DRAM_mem[4][26] ), .B(\DRAM_mem[20][26] ), .S(n167), .Z(
        n982) );
  MUX2_X1 U1043 ( .A(n982), .B(n981), .S(n131), .Z(n983) );
  MUX2_X1 U1044 ( .A(\DRAM_mem[8][26] ), .B(\DRAM_mem[24][26] ), .S(n167), .Z(
        n984) );
  MUX2_X1 U1045 ( .A(\DRAM_mem[0][26] ), .B(\DRAM_mem[16][26] ), .S(n167), .Z(
        n985) );
  MUX2_X1 U1046 ( .A(n985), .B(n984), .S(n131), .Z(n986) );
  MUX2_X1 U1047 ( .A(n986), .B(n983), .S(n110), .Z(n987) );
  MUX2_X1 U1048 ( .A(n987), .B(n980), .S(Addr[0]), .Z(n988) );
  MUX2_X1 U1049 ( .A(n988), .B(n973), .S(Addr[1]), .Z(N391) );
  MUX2_X1 U1050 ( .A(\DRAM_mem[15][27] ), .B(\DRAM_mem[31][27] ), .S(n168), 
        .Z(n989) );
  MUX2_X1 U1051 ( .A(\DRAM_mem[7][27] ), .B(\DRAM_mem[23][27] ), .S(n168), .Z(
        n990) );
  MUX2_X1 U1052 ( .A(n990), .B(n989), .S(n117), .Z(n991) );
  MUX2_X1 U1053 ( .A(\DRAM_mem[11][27] ), .B(\DRAM_mem[27][27] ), .S(n168), 
        .Z(n992) );
  MUX2_X1 U1054 ( .A(\DRAM_mem[3][27] ), .B(\DRAM_mem[19][27] ), .S(n168), .Z(
        n993) );
  MUX2_X1 U1055 ( .A(n993), .B(n992), .S(n116), .Z(n994) );
  MUX2_X1 U1056 ( .A(n994), .B(n991), .S(n111), .Z(n995) );
  MUX2_X1 U1057 ( .A(\DRAM_mem[14][27] ), .B(\DRAM_mem[30][27] ), .S(n168), 
        .Z(n996) );
  MUX2_X1 U1058 ( .A(\DRAM_mem[6][27] ), .B(\DRAM_mem[22][27] ), .S(n168), .Z(
        n997) );
  MUX2_X1 U1059 ( .A(n997), .B(n996), .S(n115), .Z(n998) );
  MUX2_X1 U1060 ( .A(\DRAM_mem[10][27] ), .B(\DRAM_mem[26][27] ), .S(n168), 
        .Z(n999) );
  MUX2_X1 U1061 ( .A(\DRAM_mem[2][27] ), .B(\DRAM_mem[18][27] ), .S(n168), .Z(
        n1000) );
  MUX2_X1 U1062 ( .A(n1000), .B(n999), .S(n114), .Z(n1001) );
  MUX2_X1 U1063 ( .A(n1001), .B(n998), .S(n111), .Z(n1002) );
  MUX2_X1 U1064 ( .A(n1002), .B(n995), .S(Addr[0]), .Z(n1003) );
  MUX2_X1 U1065 ( .A(\DRAM_mem[13][27] ), .B(\DRAM_mem[29][27] ), .S(n168), 
        .Z(n1004) );
  MUX2_X1 U1066 ( .A(\DRAM_mem[5][27] ), .B(\DRAM_mem[21][27] ), .S(n168), .Z(
        n1005) );
  MUX2_X1 U1067 ( .A(n1005), .B(n1004), .S(n131), .Z(n1006) );
  MUX2_X1 U1068 ( .A(\DRAM_mem[9][27] ), .B(\DRAM_mem[25][27] ), .S(n168), .Z(
        n1007) );
  MUX2_X1 U1069 ( .A(\DRAM_mem[1][27] ), .B(\DRAM_mem[17][27] ), .S(n168), .Z(
        n1008) );
  MUX2_X1 U1070 ( .A(n1008), .B(n1007), .S(n130), .Z(n1009) );
  MUX2_X1 U1071 ( .A(n1009), .B(n1006), .S(n111), .Z(n1010) );
  MUX2_X1 U1072 ( .A(\DRAM_mem[12][27] ), .B(\DRAM_mem[28][27] ), .S(n169), 
        .Z(n1011) );
  MUX2_X1 U1073 ( .A(\DRAM_mem[4][27] ), .B(\DRAM_mem[20][27] ), .S(n169), .Z(
        n1012) );
  MUX2_X1 U1074 ( .A(n1012), .B(n1011), .S(n129), .Z(n1013) );
  MUX2_X1 U1075 ( .A(\DRAM_mem[8][27] ), .B(\DRAM_mem[24][27] ), .S(n169), .Z(
        n1014) );
  MUX2_X1 U1076 ( .A(\DRAM_mem[0][27] ), .B(\DRAM_mem[16][27] ), .S(n169), .Z(
        n1015) );
  MUX2_X1 U1077 ( .A(n1015), .B(n1014), .S(n128), .Z(n1016) );
  MUX2_X1 U1078 ( .A(n1016), .B(n1013), .S(n111), .Z(n1017) );
  MUX2_X1 U1079 ( .A(n1017), .B(n1010), .S(Addr[0]), .Z(n1018) );
  MUX2_X1 U1080 ( .A(n1018), .B(n1003), .S(Addr[1]), .Z(N390) );
  MUX2_X1 U1081 ( .A(\DRAM_mem[15][28] ), .B(\DRAM_mem[31][28] ), .S(n169), 
        .Z(n1019) );
  MUX2_X1 U1082 ( .A(\DRAM_mem[7][28] ), .B(\DRAM_mem[23][28] ), .S(n169), .Z(
        n1020) );
  MUX2_X1 U1083 ( .A(n1020), .B(n1019), .S(n127), .Z(n1021) );
  MUX2_X1 U1084 ( .A(\DRAM_mem[11][28] ), .B(\DRAM_mem[27][28] ), .S(n169), 
        .Z(n1022) );
  MUX2_X1 U1085 ( .A(\DRAM_mem[3][28] ), .B(\DRAM_mem[19][28] ), .S(n169), .Z(
        n1023) );
  MUX2_X1 U1086 ( .A(n1023), .B(n1022), .S(n126), .Z(n1024) );
  MUX2_X1 U1087 ( .A(n1024), .B(n1021), .S(n111), .Z(n1025) );
  MUX2_X1 U1088 ( .A(\DRAM_mem[14][28] ), .B(\DRAM_mem[30][28] ), .S(n169), 
        .Z(n1026) );
  MUX2_X1 U1089 ( .A(\DRAM_mem[6][28] ), .B(\DRAM_mem[22][28] ), .S(n169), .Z(
        n1027) );
  MUX2_X1 U1090 ( .A(n1027), .B(n1026), .S(n125), .Z(n1028) );
  MUX2_X1 U1091 ( .A(\DRAM_mem[10][28] ), .B(\DRAM_mem[26][28] ), .S(n169), 
        .Z(n1029) );
  MUX2_X1 U1092 ( .A(\DRAM_mem[2][28] ), .B(\DRAM_mem[18][28] ), .S(n169), .Z(
        n1030) );
  MUX2_X1 U1093 ( .A(n1030), .B(n1029), .S(n124), .Z(n1031) );
  MUX2_X1 U1094 ( .A(n1031), .B(n1028), .S(n111), .Z(n1032) );
  MUX2_X1 U1095 ( .A(n1032), .B(n1025), .S(Addr[0]), .Z(n1033) );
  MUX2_X1 U1096 ( .A(\DRAM_mem[13][28] ), .B(\DRAM_mem[29][28] ), .S(n170), 
        .Z(n1034) );
  MUX2_X1 U1097 ( .A(\DRAM_mem[5][28] ), .B(\DRAM_mem[21][28] ), .S(n170), .Z(
        n1035) );
  MUX2_X1 U1098 ( .A(n1035), .B(n1034), .S(n123), .Z(n1036) );
  MUX2_X1 U1099 ( .A(\DRAM_mem[9][28] ), .B(\DRAM_mem[25][28] ), .S(n170), .Z(
        n1037) );
  MUX2_X1 U1100 ( .A(\DRAM_mem[1][28] ), .B(\DRAM_mem[17][28] ), .S(n170), .Z(
        n1038) );
  MUX2_X1 U1101 ( .A(n1038), .B(n1037), .S(n122), .Z(n1039) );
  MUX2_X1 U1102 ( .A(n1039), .B(n1036), .S(n111), .Z(n1040) );
  MUX2_X1 U1103 ( .A(\DRAM_mem[12][28] ), .B(\DRAM_mem[28][28] ), .S(n170), 
        .Z(n1041) );
  MUX2_X1 U1104 ( .A(\DRAM_mem[4][28] ), .B(\DRAM_mem[20][28] ), .S(n170), .Z(
        n1042) );
  MUX2_X1 U1105 ( .A(n1042), .B(n1041), .S(n121), .Z(n1043) );
  MUX2_X1 U1106 ( .A(\DRAM_mem[8][28] ), .B(\DRAM_mem[24][28] ), .S(n170), .Z(
        n1044) );
  MUX2_X1 U1107 ( .A(\DRAM_mem[0][28] ), .B(\DRAM_mem[16][28] ), .S(n170), .Z(
        n1045) );
  MUX2_X1 U1108 ( .A(n1045), .B(n1044), .S(n120), .Z(n1046) );
  MUX2_X1 U1109 ( .A(n1046), .B(n1043), .S(n111), .Z(n1047) );
  MUX2_X1 U1110 ( .A(n1047), .B(n1040), .S(Addr[0]), .Z(n1048) );
  MUX2_X1 U1111 ( .A(n1048), .B(n1033), .S(Addr[1]), .Z(N389) );
  MUX2_X1 U1112 ( .A(\DRAM_mem[15][29] ), .B(\DRAM_mem[31][29] ), .S(n170), 
        .Z(n1049) );
  MUX2_X1 U1113 ( .A(\DRAM_mem[7][29] ), .B(\DRAM_mem[23][29] ), .S(n170), .Z(
        n1050) );
  MUX2_X1 U1114 ( .A(n1050), .B(n1049), .S(n119), .Z(n1051) );
  MUX2_X1 U1115 ( .A(\DRAM_mem[11][29] ), .B(\DRAM_mem[27][29] ), .S(n170), 
        .Z(n1052) );
  MUX2_X1 U1116 ( .A(\DRAM_mem[3][29] ), .B(\DRAM_mem[19][29] ), .S(n170), .Z(
        n1053) );
  MUX2_X1 U1117 ( .A(n1053), .B(n1052), .S(n118), .Z(n1054) );
  MUX2_X1 U1118 ( .A(n1054), .B(n1051), .S(n111), .Z(n1055) );
  MUX2_X1 U1119 ( .A(\DRAM_mem[14][29] ), .B(\DRAM_mem[30][29] ), .S(n159), 
        .Z(n1056) );
  MUX2_X1 U1120 ( .A(\DRAM_mem[6][29] ), .B(\DRAM_mem[22][29] ), .S(n158), .Z(
        n1057) );
  MUX2_X1 U1121 ( .A(n1057), .B(n1056), .S(n117), .Z(n1058) );
  MUX2_X1 U1122 ( .A(\DRAM_mem[10][29] ), .B(\DRAM_mem[26][29] ), .S(n157), 
        .Z(n1059) );
  MUX2_X1 U1123 ( .A(\DRAM_mem[2][29] ), .B(\DRAM_mem[18][29] ), .S(n156), .Z(
        n1060) );
  MUX2_X1 U1124 ( .A(n1060), .B(n1059), .S(n116), .Z(n1061) );
  MUX2_X1 U1125 ( .A(n1061), .B(n1058), .S(n111), .Z(n1062) );
  MUX2_X1 U1126 ( .A(n1062), .B(n1055), .S(Addr[0]), .Z(n1063) );
  MUX2_X1 U1127 ( .A(\DRAM_mem[13][29] ), .B(\DRAM_mem[29][29] ), .S(n155), 
        .Z(n1064) );
  MUX2_X1 U1128 ( .A(\DRAM_mem[5][29] ), .B(\DRAM_mem[21][29] ), .S(n154), .Z(
        n1065) );
  MUX2_X1 U1129 ( .A(n1065), .B(n1064), .S(n115), .Z(n1066) );
  MUX2_X1 U1130 ( .A(\DRAM_mem[9][29] ), .B(\DRAM_mem[25][29] ), .S(Addr[4]), 
        .Z(n1067) );
  MUX2_X1 U1131 ( .A(\DRAM_mem[1][29] ), .B(\DRAM_mem[17][29] ), .S(n164), .Z(
        n1068) );
  MUX2_X1 U1132 ( .A(n1068), .B(n1067), .S(n114), .Z(n1069) );
  MUX2_X1 U1133 ( .A(n1069), .B(n1066), .S(n111), .Z(n1070) );
  MUX2_X1 U1134 ( .A(\DRAM_mem[12][29] ), .B(\DRAM_mem[28][29] ), .S(n163), 
        .Z(n1071) );
  MUX2_X1 U1135 ( .A(\DRAM_mem[4][29] ), .B(\DRAM_mem[20][29] ), .S(n170), .Z(
        n1072) );
  MUX2_X1 U1136 ( .A(n1072), .B(n1071), .S(Addr[3]), .Z(n1073) );
  MUX2_X1 U1137 ( .A(\DRAM_mem[8][29] ), .B(\DRAM_mem[24][29] ), .S(n169), .Z(
        n1074) );
  MUX2_X1 U1138 ( .A(\DRAM_mem[0][29] ), .B(\DRAM_mem[16][29] ), .S(n168), .Z(
        n1075) );
  MUX2_X1 U1139 ( .A(n1075), .B(n1074), .S(n131), .Z(n1076) );
  MUX2_X1 U1140 ( .A(n1076), .B(n1073), .S(n111), .Z(n1077) );
  MUX2_X1 U1141 ( .A(n1077), .B(n1070), .S(Addr[0]), .Z(n1078) );
  MUX2_X1 U1142 ( .A(n1078), .B(n1063), .S(Addr[1]), .Z(N388) );
  MUX2_X1 U1143 ( .A(\DRAM_mem[15][30] ), .B(\DRAM_mem[31][30] ), .S(n146), 
        .Z(n1079) );
  MUX2_X1 U1144 ( .A(\DRAM_mem[7][30] ), .B(\DRAM_mem[23][30] ), .S(n145), .Z(
        n1080) );
  MUX2_X1 U1145 ( .A(n1080), .B(n1079), .S(n130), .Z(n1081) );
  MUX2_X1 U1146 ( .A(\DRAM_mem[11][30] ), .B(\DRAM_mem[27][30] ), .S(n144), 
        .Z(n1082) );
  MUX2_X1 U1147 ( .A(\DRAM_mem[3][30] ), .B(\DRAM_mem[19][30] ), .S(n143), .Z(
        n1083) );
  MUX2_X1 U1148 ( .A(n1083), .B(n1082), .S(n129), .Z(n1084) );
  MUX2_X1 U1149 ( .A(n1084), .B(n1081), .S(n112), .Z(n1085) );
  MUX2_X1 U1150 ( .A(\DRAM_mem[14][30] ), .B(\DRAM_mem[30][30] ), .S(n142), 
        .Z(n1086) );
  MUX2_X1 U1151 ( .A(\DRAM_mem[6][30] ), .B(\DRAM_mem[22][30] ), .S(n141), .Z(
        n1087) );
  MUX2_X1 U1152 ( .A(n1087), .B(n1086), .S(n128), .Z(n1088) );
  MUX2_X1 U1153 ( .A(\DRAM_mem[10][30] ), .B(\DRAM_mem[26][30] ), .S(n140), 
        .Z(n1089) );
  MUX2_X1 U1154 ( .A(\DRAM_mem[2][30] ), .B(\DRAM_mem[18][30] ), .S(n139), .Z(
        n1090) );
  MUX2_X1 U1155 ( .A(n1090), .B(n1089), .S(n127), .Z(n1091) );
  MUX2_X1 U1156 ( .A(n1091), .B(n1088), .S(n112), .Z(n1092) );
  MUX2_X1 U1157 ( .A(n1092), .B(n1085), .S(Addr[0]), .Z(n1093) );
  MUX2_X1 U1158 ( .A(\DRAM_mem[13][30] ), .B(\DRAM_mem[29][30] ), .S(n138), 
        .Z(n1094) );
  MUX2_X1 U1159 ( .A(\DRAM_mem[5][30] ), .B(\DRAM_mem[21][30] ), .S(n137), .Z(
        n1095) );
  MUX2_X1 U1160 ( .A(n1095), .B(n1094), .S(n126), .Z(n1096) );
  MUX2_X1 U1161 ( .A(\DRAM_mem[9][30] ), .B(\DRAM_mem[25][30] ), .S(n136), .Z(
        n1097) );
  MUX2_X1 U1162 ( .A(\DRAM_mem[1][30] ), .B(\DRAM_mem[17][30] ), .S(n135), .Z(
        n1098) );
  MUX2_X1 U1163 ( .A(n1098), .B(n1097), .S(n125), .Z(n1099) );
  MUX2_X1 U1164 ( .A(n1099), .B(n1096), .S(n112), .Z(n1100) );
  MUX2_X1 U1165 ( .A(\DRAM_mem[12][30] ), .B(\DRAM_mem[28][30] ), .S(n134), 
        .Z(n1101) );
  MUX2_X1 U1166 ( .A(\DRAM_mem[4][30] ), .B(\DRAM_mem[20][30] ), .S(n133), .Z(
        n1102) );
  MUX2_X1 U1167 ( .A(n1102), .B(n1101), .S(n124), .Z(n1103) );
  MUX2_X1 U1168 ( .A(\DRAM_mem[8][30] ), .B(\DRAM_mem[24][30] ), .S(n153), .Z(
        n1104) );
  MUX2_X1 U1169 ( .A(\DRAM_mem[0][30] ), .B(\DRAM_mem[16][30] ), .S(n152), .Z(
        n1105) );
  MUX2_X1 U1170 ( .A(n1105), .B(n1104), .S(Addr[3]), .Z(n1106) );
  MUX2_X1 U1171 ( .A(n1106), .B(n1103), .S(n112), .Z(n1107) );
  MUX2_X1 U1172 ( .A(n1107), .B(n1100), .S(Addr[0]), .Z(n1108) );
  MUX2_X1 U1173 ( .A(n1108), .B(n1093), .S(Addr[1]), .Z(N387) );
  MUX2_X1 U1174 ( .A(\DRAM_mem[15][31] ), .B(\DRAM_mem[31][31] ), .S(n151), 
        .Z(n1109) );
  MUX2_X1 U1175 ( .A(\DRAM_mem[7][31] ), .B(\DRAM_mem[23][31] ), .S(n150), .Z(
        n1110) );
  MUX2_X1 U1176 ( .A(n1110), .B(n1109), .S(Addr[3]), .Z(n1111) );
  MUX2_X1 U1177 ( .A(\DRAM_mem[11][31] ), .B(\DRAM_mem[27][31] ), .S(n149), 
        .Z(n1112) );
  MUX2_X1 U1178 ( .A(\DRAM_mem[3][31] ), .B(\DRAM_mem[19][31] ), .S(n148), .Z(
        n1113) );
  MUX2_X1 U1179 ( .A(n1113), .B(n1112), .S(Addr[3]), .Z(n1114) );
  MUX2_X1 U1180 ( .A(n1114), .B(n1111), .S(n112), .Z(n1115) );
  MUX2_X1 U1181 ( .A(\DRAM_mem[14][31] ), .B(\DRAM_mem[30][31] ), .S(n147), 
        .Z(n1116) );
  MUX2_X1 U1182 ( .A(\DRAM_mem[6][31] ), .B(\DRAM_mem[22][31] ), .S(n167), .Z(
        n1117) );
  MUX2_X1 U1183 ( .A(n1117), .B(n1116), .S(Addr[3]), .Z(n1118) );
  MUX2_X1 U1184 ( .A(\DRAM_mem[10][31] ), .B(\DRAM_mem[26][31] ), .S(n166), 
        .Z(n1119) );
  MUX2_X1 U1185 ( .A(\DRAM_mem[2][31] ), .B(\DRAM_mem[18][31] ), .S(n165), .Z(
        n1120) );
  MUX2_X1 U1186 ( .A(n1120), .B(n1119), .S(Addr[3]), .Z(n1121) );
  MUX2_X1 U1187 ( .A(n1121), .B(n1118), .S(n112), .Z(n1122) );
  MUX2_X1 U1188 ( .A(n1122), .B(n1115), .S(Addr[0]), .Z(n1123) );
  MUX2_X1 U1189 ( .A(\DRAM_mem[13][31] ), .B(\DRAM_mem[29][31] ), .S(n162), 
        .Z(n1124) );
  MUX2_X1 U1190 ( .A(\DRAM_mem[5][31] ), .B(\DRAM_mem[21][31] ), .S(n161), .Z(
        n1125) );
  MUX2_X1 U1191 ( .A(n1125), .B(n1124), .S(Addr[3]), .Z(n1126) );
  MUX2_X1 U1192 ( .A(\DRAM_mem[9][31] ), .B(\DRAM_mem[25][31] ), .S(n160), .Z(
        n1127) );
  MUX2_X1 U1193 ( .A(\DRAM_mem[1][31] ), .B(\DRAM_mem[17][31] ), .S(n159), .Z(
        n1128) );
  MUX2_X1 U1194 ( .A(n1128), .B(n1127), .S(Addr[3]), .Z(n1129) );
  MUX2_X1 U1195 ( .A(n1129), .B(n1126), .S(n112), .Z(n1130) );
  MUX2_X1 U1196 ( .A(\DRAM_mem[12][31] ), .B(\DRAM_mem[28][31] ), .S(n158), 
        .Z(n1131) );
  MUX2_X1 U1197 ( .A(\DRAM_mem[4][31] ), .B(\DRAM_mem[20][31] ), .S(n157), .Z(
        n1132) );
  MUX2_X1 U1198 ( .A(n1132), .B(n1131), .S(Addr[3]), .Z(n1133) );
  MUX2_X1 U1199 ( .A(\DRAM_mem[8][31] ), .B(\DRAM_mem[24][31] ), .S(n156), .Z(
        n1134) );
  MUX2_X1 U1200 ( .A(\DRAM_mem[0][31] ), .B(\DRAM_mem[16][31] ), .S(n155), .Z(
        n1135) );
  MUX2_X1 U1201 ( .A(n1135), .B(n1134), .S(Addr[3]), .Z(n1136) );
  MUX2_X1 U1202 ( .A(n1136), .B(n1133), .S(n112), .Z(n1137) );
  MUX2_X1 U1203 ( .A(n1137), .B(n1130), .S(Addr[0]), .Z(n1138) );
  MUX2_X1 U1204 ( .A(n1138), .B(n1123), .S(Addr[1]), .Z(N386) );
  INV_X1 U1205 ( .A(Rst), .ZN(n2309) );
  MUX2_X1 U1206 ( .A(\DRAM_mem[0][31] ), .B(n1139), .S(n1140), .Z(n2180) );
  MUX2_X1 U1207 ( .A(\DRAM_mem[0][30] ), .B(n1141), .S(n1140), .Z(n2179) );
  MUX2_X1 U1208 ( .A(\DRAM_mem[0][29] ), .B(n1142), .S(n1140), .Z(n2178) );
  MUX2_X1 U1209 ( .A(\DRAM_mem[0][28] ), .B(n1143), .S(n1140), .Z(n2177) );
  MUX2_X1 U1210 ( .A(\DRAM_mem[0][27] ), .B(n1144), .S(n1140), .Z(n2176) );
  MUX2_X1 U1211 ( .A(\DRAM_mem[0][26] ), .B(n1145), .S(n1140), .Z(n2175) );
  MUX2_X1 U1212 ( .A(\DRAM_mem[0][25] ), .B(n1146), .S(n1140), .Z(n2174) );
  MUX2_X1 U1213 ( .A(\DRAM_mem[0][24] ), .B(n1147), .S(n1140), .Z(n2173) );
  MUX2_X1 U1214 ( .A(\DRAM_mem[0][23] ), .B(n1148), .S(n1140), .Z(n2172) );
  MUX2_X1 U1215 ( .A(\DRAM_mem[0][22] ), .B(n1149), .S(n1140), .Z(n2171) );
  MUX2_X1 U1216 ( .A(\DRAM_mem[0][21] ), .B(n1150), .S(n1140), .Z(n2170) );
  MUX2_X1 U1217 ( .A(\DRAM_mem[0][20] ), .B(n1151), .S(n1140), .Z(n2169) );
  MUX2_X1 U1218 ( .A(\DRAM_mem[0][19] ), .B(n1152), .S(n1140), .Z(n2168) );
  MUX2_X1 U1219 ( .A(\DRAM_mem[0][18] ), .B(n1153), .S(n1140), .Z(n2167) );
  MUX2_X1 U1220 ( .A(\DRAM_mem[0][17] ), .B(n1154), .S(n1140), .Z(n2166) );
  MUX2_X1 U1221 ( .A(\DRAM_mem[0][16] ), .B(n1155), .S(n1140), .Z(n2165) );
  MUX2_X1 U1222 ( .A(\DRAM_mem[0][15] ), .B(n1156), .S(n1140), .Z(n2164) );
  MUX2_X1 U1223 ( .A(\DRAM_mem[0][14] ), .B(n2181), .S(n1140), .Z(n2163) );
  MUX2_X1 U1224 ( .A(\DRAM_mem[0][13] ), .B(n2182), .S(n1140), .Z(n2162) );
  MUX2_X1 U1225 ( .A(\DRAM_mem[0][12] ), .B(n2183), .S(n1140), .Z(n2161) );
  MUX2_X1 U1226 ( .A(\DRAM_mem[0][11] ), .B(n2184), .S(n1140), .Z(n2160) );
  MUX2_X1 U1227 ( .A(\DRAM_mem[0][10] ), .B(n2185), .S(n1140), .Z(n2159) );
  MUX2_X1 U1228 ( .A(\DRAM_mem[0][9] ), .B(n2186), .S(n1140), .Z(n2158) );
  MUX2_X1 U1229 ( .A(\DRAM_mem[0][8] ), .B(n2187), .S(n1140), .Z(n2157) );
  MUX2_X1 U1230 ( .A(\DRAM_mem[0][7] ), .B(n2188), .S(n1140), .Z(n2156) );
  MUX2_X1 U1231 ( .A(\DRAM_mem[0][6] ), .B(n2189), .S(n1140), .Z(n2155) );
  MUX2_X1 U1232 ( .A(\DRAM_mem[0][5] ), .B(n2190), .S(n1140), .Z(n2154) );
  MUX2_X1 U1233 ( .A(\DRAM_mem[0][4] ), .B(n2191), .S(n1140), .Z(n2153) );
  MUX2_X1 U1234 ( .A(\DRAM_mem[0][3] ), .B(n2192), .S(n1140), .Z(n2152) );
  MUX2_X1 U1235 ( .A(\DRAM_mem[0][2] ), .B(n2193), .S(n1140), .Z(n2151) );
  MUX2_X1 U1236 ( .A(\DRAM_mem[0][1] ), .B(n2194), .S(n1140), .Z(n2150) );
  MUX2_X1 U1237 ( .A(\DRAM_mem[0][0] ), .B(n2195), .S(n1140), .Z(n2149) );
  MUX2_X1 U1238 ( .A(\DRAM_mem[1][31] ), .B(n1139), .S(n2198), .Z(n2148) );
  MUX2_X1 U1239 ( .A(\DRAM_mem[1][30] ), .B(n1141), .S(n2198), .Z(n2147) );
  MUX2_X1 U1240 ( .A(\DRAM_mem[1][29] ), .B(n1142), .S(n2198), .Z(n2146) );
  MUX2_X1 U1241 ( .A(\DRAM_mem[1][28] ), .B(n1143), .S(n2198), .Z(n2145) );
  MUX2_X1 U1242 ( .A(\DRAM_mem[1][27] ), .B(n1144), .S(n2198), .Z(n2144) );
  MUX2_X1 U1243 ( .A(\DRAM_mem[1][26] ), .B(n1145), .S(n2198), .Z(n2143) );
  MUX2_X1 U1244 ( .A(\DRAM_mem[1][25] ), .B(n1146), .S(n2198), .Z(n2142) );
  MUX2_X1 U1245 ( .A(\DRAM_mem[1][24] ), .B(n1147), .S(n2198), .Z(n2141) );
  MUX2_X1 U1246 ( .A(\DRAM_mem[1][23] ), .B(n1148), .S(n2198), .Z(n2140) );
  MUX2_X1 U1247 ( .A(\DRAM_mem[1][22] ), .B(n1149), .S(n2198), .Z(n2139) );
  MUX2_X1 U1248 ( .A(\DRAM_mem[1][21] ), .B(n1150), .S(n2198), .Z(n2138) );
  MUX2_X1 U1249 ( .A(\DRAM_mem[1][20] ), .B(n1151), .S(n2198), .Z(n2137) );
  MUX2_X1 U1250 ( .A(\DRAM_mem[1][19] ), .B(n1152), .S(n2198), .Z(n2136) );
  MUX2_X1 U1251 ( .A(\DRAM_mem[1][18] ), .B(n1153), .S(n2198), .Z(n2135) );
  MUX2_X1 U1252 ( .A(\DRAM_mem[1][17] ), .B(n1154), .S(n2198), .Z(n2134) );
  MUX2_X1 U1253 ( .A(\DRAM_mem[1][16] ), .B(n1155), .S(n2198), .Z(n2133) );
  MUX2_X1 U1254 ( .A(\DRAM_mem[1][15] ), .B(n1156), .S(n2198), .Z(n2132) );
  MUX2_X1 U1255 ( .A(\DRAM_mem[1][14] ), .B(n2181), .S(n2198), .Z(n2131) );
  MUX2_X1 U1256 ( .A(\DRAM_mem[1][13] ), .B(n2182), .S(n2198), .Z(n2130) );
  MUX2_X1 U1257 ( .A(\DRAM_mem[1][12] ), .B(n2183), .S(n2198), .Z(n2129) );
  MUX2_X1 U1258 ( .A(\DRAM_mem[1][11] ), .B(n2184), .S(n2198), .Z(n2128) );
  MUX2_X1 U1259 ( .A(\DRAM_mem[1][10] ), .B(n2185), .S(n2198), .Z(n2127) );
  MUX2_X1 U1260 ( .A(\DRAM_mem[1][9] ), .B(n2186), .S(n2198), .Z(n2126) );
  MUX2_X1 U1261 ( .A(\DRAM_mem[1][8] ), .B(n2187), .S(n2198), .Z(n2125) );
  MUX2_X1 U1262 ( .A(\DRAM_mem[1][7] ), .B(n2188), .S(n2198), .Z(n2124) );
  MUX2_X1 U1263 ( .A(\DRAM_mem[1][6] ), .B(n2189), .S(n2198), .Z(n2123) );
  MUX2_X1 U1264 ( .A(\DRAM_mem[1][5] ), .B(n2190), .S(n2198), .Z(n2122) );
  MUX2_X1 U1265 ( .A(\DRAM_mem[1][4] ), .B(n2191), .S(n2198), .Z(n2121) );
  MUX2_X1 U1266 ( .A(\DRAM_mem[1][3] ), .B(n2192), .S(n2198), .Z(n2120) );
  MUX2_X1 U1267 ( .A(\DRAM_mem[1][2] ), .B(n2193), .S(n2198), .Z(n2119) );
  MUX2_X1 U1268 ( .A(\DRAM_mem[1][1] ), .B(n2194), .S(n2198), .Z(n2118) );
  MUX2_X1 U1269 ( .A(\DRAM_mem[1][0] ), .B(n2195), .S(n2198), .Z(n2117) );
  MUX2_X1 U1270 ( .A(\DRAM_mem[2][31] ), .B(n1139), .S(n2200), .Z(n2116) );
  MUX2_X1 U1271 ( .A(\DRAM_mem[2][30] ), .B(n1141), .S(n2200), .Z(n2115) );
  MUX2_X1 U1272 ( .A(\DRAM_mem[2][29] ), .B(n1142), .S(n2200), .Z(n2114) );
  MUX2_X1 U1273 ( .A(\DRAM_mem[2][28] ), .B(n1143), .S(n2200), .Z(n2113) );
  MUX2_X1 U1274 ( .A(\DRAM_mem[2][27] ), .B(n1144), .S(n2200), .Z(n2112) );
  MUX2_X1 U1275 ( .A(\DRAM_mem[2][26] ), .B(n1145), .S(n2200), .Z(n2111) );
  MUX2_X1 U1276 ( .A(\DRAM_mem[2][25] ), .B(n1146), .S(n2200), .Z(n2110) );
  MUX2_X1 U1277 ( .A(\DRAM_mem[2][24] ), .B(n1147), .S(n2200), .Z(n2109) );
  MUX2_X1 U1278 ( .A(\DRAM_mem[2][23] ), .B(n1148), .S(n2200), .Z(n2108) );
  MUX2_X1 U1279 ( .A(\DRAM_mem[2][22] ), .B(n1149), .S(n2200), .Z(n2107) );
  MUX2_X1 U1280 ( .A(\DRAM_mem[2][21] ), .B(n1150), .S(n2200), .Z(n2106) );
  MUX2_X1 U1281 ( .A(\DRAM_mem[2][20] ), .B(n1151), .S(n2200), .Z(n2105) );
  MUX2_X1 U1282 ( .A(\DRAM_mem[2][19] ), .B(n1152), .S(n2200), .Z(n2104) );
  MUX2_X1 U1283 ( .A(\DRAM_mem[2][18] ), .B(n1153), .S(n2200), .Z(n2103) );
  MUX2_X1 U1284 ( .A(\DRAM_mem[2][17] ), .B(n1154), .S(n2200), .Z(n2102) );
  MUX2_X1 U1285 ( .A(\DRAM_mem[2][16] ), .B(n1155), .S(n2200), .Z(n2101) );
  MUX2_X1 U1286 ( .A(\DRAM_mem[2][15] ), .B(n1156), .S(n2200), .Z(n2100) );
  MUX2_X1 U1287 ( .A(\DRAM_mem[2][14] ), .B(n2181), .S(n2200), .Z(n2099) );
  MUX2_X1 U1288 ( .A(\DRAM_mem[2][13] ), .B(n2182), .S(n2200), .Z(n2098) );
  MUX2_X1 U1289 ( .A(\DRAM_mem[2][12] ), .B(n2183), .S(n2200), .Z(n2097) );
  MUX2_X1 U1290 ( .A(\DRAM_mem[2][11] ), .B(n2184), .S(n2200), .Z(n2096) );
  MUX2_X1 U1291 ( .A(\DRAM_mem[2][10] ), .B(n2185), .S(n2200), .Z(n2095) );
  MUX2_X1 U1292 ( .A(\DRAM_mem[2][9] ), .B(n2186), .S(n2200), .Z(n2094) );
  MUX2_X1 U1293 ( .A(\DRAM_mem[2][8] ), .B(n2187), .S(n2200), .Z(n2093) );
  MUX2_X1 U1294 ( .A(\DRAM_mem[2][7] ), .B(n2188), .S(n2200), .Z(n2092) );
  MUX2_X1 U1295 ( .A(\DRAM_mem[2][6] ), .B(n2189), .S(n2200), .Z(n2091) );
  MUX2_X1 U1296 ( .A(\DRAM_mem[2][5] ), .B(n2190), .S(n2200), .Z(n2090) );
  MUX2_X1 U1297 ( .A(\DRAM_mem[2][4] ), .B(n2191), .S(n2200), .Z(n2089) );
  MUX2_X1 U1298 ( .A(\DRAM_mem[2][3] ), .B(n2192), .S(n2200), .Z(n2088) );
  MUX2_X1 U1299 ( .A(\DRAM_mem[2][2] ), .B(n2193), .S(n2200), .Z(n2087) );
  MUX2_X1 U1300 ( .A(\DRAM_mem[2][1] ), .B(n2194), .S(n2200), .Z(n2086) );
  MUX2_X1 U1301 ( .A(\DRAM_mem[2][0] ), .B(n2195), .S(n2200), .Z(n2085) );
  MUX2_X1 U1302 ( .A(\DRAM_mem[3][31] ), .B(n1139), .S(n2202), .Z(n2084) );
  MUX2_X1 U1303 ( .A(\DRAM_mem[3][30] ), .B(n1141), .S(n2202), .Z(n2083) );
  MUX2_X1 U1304 ( .A(\DRAM_mem[3][29] ), .B(n1142), .S(n2202), .Z(n2082) );
  MUX2_X1 U1305 ( .A(\DRAM_mem[3][28] ), .B(n1143), .S(n2202), .Z(n2081) );
  MUX2_X1 U1306 ( .A(\DRAM_mem[3][27] ), .B(n1144), .S(n2202), .Z(n2080) );
  MUX2_X1 U1307 ( .A(\DRAM_mem[3][26] ), .B(n1145), .S(n2202), .Z(n2079) );
  MUX2_X1 U1308 ( .A(\DRAM_mem[3][25] ), .B(n1146), .S(n2202), .Z(n2078) );
  MUX2_X1 U1309 ( .A(\DRAM_mem[3][24] ), .B(n1147), .S(n2202), .Z(n2077) );
  MUX2_X1 U1310 ( .A(\DRAM_mem[3][23] ), .B(n1148), .S(n2202), .Z(n2076) );
  MUX2_X1 U1311 ( .A(\DRAM_mem[3][22] ), .B(n1149), .S(n2202), .Z(n2075) );
  MUX2_X1 U1312 ( .A(\DRAM_mem[3][21] ), .B(n1150), .S(n2202), .Z(n2074) );
  MUX2_X1 U1313 ( .A(\DRAM_mem[3][20] ), .B(n1151), .S(n2202), .Z(n2073) );
  MUX2_X1 U1314 ( .A(\DRAM_mem[3][19] ), .B(n1152), .S(n2202), .Z(n2072) );
  MUX2_X1 U1315 ( .A(\DRAM_mem[3][18] ), .B(n1153), .S(n2202), .Z(n2071) );
  MUX2_X1 U1316 ( .A(\DRAM_mem[3][17] ), .B(n1154), .S(n2202), .Z(n2070) );
  MUX2_X1 U1317 ( .A(\DRAM_mem[3][16] ), .B(n1155), .S(n2202), .Z(n2069) );
  MUX2_X1 U1318 ( .A(\DRAM_mem[3][15] ), .B(n1156), .S(n2202), .Z(n2068) );
  MUX2_X1 U1319 ( .A(\DRAM_mem[3][14] ), .B(n2181), .S(n2202), .Z(n2067) );
  MUX2_X1 U1320 ( .A(\DRAM_mem[3][13] ), .B(n2182), .S(n2202), .Z(n2066) );
  MUX2_X1 U1321 ( .A(\DRAM_mem[3][12] ), .B(n2183), .S(n2202), .Z(n2065) );
  MUX2_X1 U1322 ( .A(\DRAM_mem[3][11] ), .B(n2184), .S(n2202), .Z(n2064) );
  MUX2_X1 U1323 ( .A(\DRAM_mem[3][10] ), .B(n2185), .S(n2202), .Z(n2063) );
  MUX2_X1 U1324 ( .A(\DRAM_mem[3][9] ), .B(n2186), .S(n2202), .Z(n2062) );
  MUX2_X1 U1325 ( .A(\DRAM_mem[3][8] ), .B(n2187), .S(n2202), .Z(n2061) );
  MUX2_X1 U1326 ( .A(\DRAM_mem[3][7] ), .B(n2188), .S(n2202), .Z(n2060) );
  MUX2_X1 U1327 ( .A(\DRAM_mem[3][6] ), .B(n2189), .S(n2202), .Z(n2059) );
  MUX2_X1 U1328 ( .A(\DRAM_mem[3][5] ), .B(n2190), .S(n2202), .Z(n2058) );
  MUX2_X1 U1329 ( .A(\DRAM_mem[3][4] ), .B(n2191), .S(n2202), .Z(n2057) );
  MUX2_X1 U1330 ( .A(\DRAM_mem[3][3] ), .B(n2192), .S(n2202), .Z(n2056) );
  MUX2_X1 U1331 ( .A(\DRAM_mem[3][2] ), .B(n2193), .S(n2202), .Z(n2055) );
  MUX2_X1 U1332 ( .A(\DRAM_mem[3][1] ), .B(n2194), .S(n2202), .Z(n2054) );
  MUX2_X1 U1333 ( .A(\DRAM_mem[3][0] ), .B(n2195), .S(n2202), .Z(n2053) );
  MUX2_X1 U1334 ( .A(\DRAM_mem[4][31] ), .B(n1139), .S(n2204), .Z(n2052) );
  MUX2_X1 U1335 ( .A(\DRAM_mem[4][30] ), .B(n1141), .S(n2204), .Z(n2051) );
  MUX2_X1 U1336 ( .A(\DRAM_mem[4][29] ), .B(n1142), .S(n2204), .Z(n2050) );
  MUX2_X1 U1337 ( .A(\DRAM_mem[4][28] ), .B(n1143), .S(n2204), .Z(n2049) );
  MUX2_X1 U1338 ( .A(\DRAM_mem[4][27] ), .B(n1144), .S(n2204), .Z(n2048) );
  MUX2_X1 U1339 ( .A(\DRAM_mem[4][26] ), .B(n1145), .S(n2204), .Z(n2047) );
  MUX2_X1 U1340 ( .A(\DRAM_mem[4][25] ), .B(n1146), .S(n2204), .Z(n2046) );
  MUX2_X1 U1341 ( .A(\DRAM_mem[4][24] ), .B(n1147), .S(n2204), .Z(n2045) );
  MUX2_X1 U1342 ( .A(\DRAM_mem[4][23] ), .B(n1148), .S(n2204), .Z(n2044) );
  MUX2_X1 U1343 ( .A(\DRAM_mem[4][22] ), .B(n1149), .S(n2204), .Z(n2043) );
  MUX2_X1 U1344 ( .A(\DRAM_mem[4][21] ), .B(n1150), .S(n2204), .Z(n2042) );
  MUX2_X1 U1345 ( .A(\DRAM_mem[4][20] ), .B(n1151), .S(n2204), .Z(n2041) );
  MUX2_X1 U1346 ( .A(\DRAM_mem[4][19] ), .B(n1152), .S(n2204), .Z(n2040) );
  MUX2_X1 U1347 ( .A(\DRAM_mem[4][18] ), .B(n1153), .S(n2204), .Z(n2039) );
  MUX2_X1 U1348 ( .A(\DRAM_mem[4][17] ), .B(n1154), .S(n2204), .Z(n2038) );
  MUX2_X1 U1349 ( .A(\DRAM_mem[4][16] ), .B(n1155), .S(n2204), .Z(n2037) );
  MUX2_X1 U1350 ( .A(\DRAM_mem[4][15] ), .B(n1156), .S(n2204), .Z(n2036) );
  MUX2_X1 U1351 ( .A(\DRAM_mem[4][14] ), .B(n2181), .S(n2204), .Z(n2035) );
  MUX2_X1 U1352 ( .A(\DRAM_mem[4][13] ), .B(n2182), .S(n2204), .Z(n2034) );
  MUX2_X1 U1353 ( .A(\DRAM_mem[4][12] ), .B(n2183), .S(n2204), .Z(n2033) );
  MUX2_X1 U1354 ( .A(\DRAM_mem[4][11] ), .B(n2184), .S(n2204), .Z(n2032) );
  MUX2_X1 U1355 ( .A(\DRAM_mem[4][10] ), .B(n2185), .S(n2204), .Z(n2031) );
  MUX2_X1 U1356 ( .A(\DRAM_mem[4][9] ), .B(n2186), .S(n2204), .Z(n2030) );
  MUX2_X1 U1357 ( .A(\DRAM_mem[4][8] ), .B(n2187), .S(n2204), .Z(n2029) );
  MUX2_X1 U1358 ( .A(\DRAM_mem[4][7] ), .B(n2188), .S(n2204), .Z(n2028) );
  MUX2_X1 U1359 ( .A(\DRAM_mem[4][6] ), .B(n2189), .S(n2204), .Z(n2027) );
  MUX2_X1 U1360 ( .A(\DRAM_mem[4][5] ), .B(n2190), .S(n2204), .Z(n2026) );
  MUX2_X1 U1361 ( .A(\DRAM_mem[4][4] ), .B(n2191), .S(n2204), .Z(n2025) );
  MUX2_X1 U1362 ( .A(\DRAM_mem[4][3] ), .B(n2192), .S(n2204), .Z(n2024) );
  MUX2_X1 U1363 ( .A(\DRAM_mem[4][2] ), .B(n2193), .S(n2204), .Z(n2023) );
  MUX2_X1 U1364 ( .A(\DRAM_mem[4][1] ), .B(n2194), .S(n2204), .Z(n2022) );
  MUX2_X1 U1365 ( .A(\DRAM_mem[4][0] ), .B(n2195), .S(n2204), .Z(n2021) );
  MUX2_X1 U1366 ( .A(\DRAM_mem[5][31] ), .B(n1139), .S(n2206), .Z(n2020) );
  MUX2_X1 U1367 ( .A(\DRAM_mem[5][30] ), .B(n1141), .S(n2206), .Z(n2019) );
  MUX2_X1 U1368 ( .A(\DRAM_mem[5][29] ), .B(n1142), .S(n2206), .Z(n2018) );
  MUX2_X1 U1369 ( .A(\DRAM_mem[5][28] ), .B(n1143), .S(n2206), .Z(n2017) );
  MUX2_X1 U1370 ( .A(\DRAM_mem[5][27] ), .B(n1144), .S(n2206), .Z(n2016) );
  MUX2_X1 U1371 ( .A(\DRAM_mem[5][26] ), .B(n1145), .S(n2206), .Z(n2015) );
  MUX2_X1 U1372 ( .A(\DRAM_mem[5][25] ), .B(n1146), .S(n2206), .Z(n2014) );
  MUX2_X1 U1373 ( .A(\DRAM_mem[5][24] ), .B(n1147), .S(n2206), .Z(n2013) );
  MUX2_X1 U1374 ( .A(\DRAM_mem[5][23] ), .B(n1148), .S(n2206), .Z(n2012) );
  MUX2_X1 U1375 ( .A(\DRAM_mem[5][22] ), .B(n1149), .S(n2206), .Z(n2011) );
  MUX2_X1 U1376 ( .A(\DRAM_mem[5][21] ), .B(n1150), .S(n2206), .Z(n2010) );
  MUX2_X1 U1377 ( .A(\DRAM_mem[5][20] ), .B(n1151), .S(n2206), .Z(n2009) );
  MUX2_X1 U1378 ( .A(\DRAM_mem[5][19] ), .B(n1152), .S(n2206), .Z(n2008) );
  MUX2_X1 U1379 ( .A(\DRAM_mem[5][18] ), .B(n1153), .S(n2206), .Z(n2007) );
  MUX2_X1 U1380 ( .A(\DRAM_mem[5][17] ), .B(n1154), .S(n2206), .Z(n2006) );
  MUX2_X1 U1381 ( .A(\DRAM_mem[5][16] ), .B(n1155), .S(n2206), .Z(n2005) );
  MUX2_X1 U1382 ( .A(\DRAM_mem[5][15] ), .B(n1156), .S(n2206), .Z(n2004) );
  MUX2_X1 U1383 ( .A(\DRAM_mem[5][14] ), .B(n2181), .S(n2206), .Z(n2003) );
  MUX2_X1 U1384 ( .A(\DRAM_mem[5][13] ), .B(n2182), .S(n2206), .Z(n2002) );
  MUX2_X1 U1385 ( .A(\DRAM_mem[5][12] ), .B(n2183), .S(n2206), .Z(n2001) );
  MUX2_X1 U1386 ( .A(\DRAM_mem[5][11] ), .B(n2184), .S(n2206), .Z(n2000) );
  MUX2_X1 U1387 ( .A(\DRAM_mem[5][10] ), .B(n2185), .S(n2206), .Z(n1999) );
  MUX2_X1 U1388 ( .A(\DRAM_mem[5][9] ), .B(n2186), .S(n2206), .Z(n1998) );
  MUX2_X1 U1389 ( .A(\DRAM_mem[5][8] ), .B(n2187), .S(n2206), .Z(n1997) );
  MUX2_X1 U1390 ( .A(\DRAM_mem[5][7] ), .B(n2188), .S(n2206), .Z(n1996) );
  MUX2_X1 U1391 ( .A(\DRAM_mem[5][6] ), .B(n2189), .S(n2206), .Z(n1995) );
  MUX2_X1 U1392 ( .A(\DRAM_mem[5][5] ), .B(n2190), .S(n2206), .Z(n1994) );
  MUX2_X1 U1393 ( .A(\DRAM_mem[5][4] ), .B(n2191), .S(n2206), .Z(n1993) );
  MUX2_X1 U1394 ( .A(\DRAM_mem[5][3] ), .B(n2192), .S(n2206), .Z(n1992) );
  MUX2_X1 U1395 ( .A(\DRAM_mem[5][2] ), .B(n2193), .S(n2206), .Z(n1991) );
  MUX2_X1 U1396 ( .A(\DRAM_mem[5][1] ), .B(n2194), .S(n2206), .Z(n1990) );
  MUX2_X1 U1397 ( .A(\DRAM_mem[5][0] ), .B(n2195), .S(n2206), .Z(n1989) );
  MUX2_X1 U1398 ( .A(\DRAM_mem[6][31] ), .B(n1139), .S(n2208), .Z(n1988) );
  MUX2_X1 U1399 ( .A(\DRAM_mem[6][30] ), .B(n1141), .S(n2208), .Z(n1987) );
  MUX2_X1 U1400 ( .A(\DRAM_mem[6][29] ), .B(n1142), .S(n2208), .Z(n1986) );
  MUX2_X1 U1401 ( .A(\DRAM_mem[6][28] ), .B(n1143), .S(n2208), .Z(n1985) );
  MUX2_X1 U1402 ( .A(\DRAM_mem[6][27] ), .B(n1144), .S(n2208), .Z(n1984) );
  MUX2_X1 U1403 ( .A(\DRAM_mem[6][26] ), .B(n1145), .S(n2208), .Z(n1983) );
  MUX2_X1 U1404 ( .A(\DRAM_mem[6][25] ), .B(n1146), .S(n2208), .Z(n1982) );
  MUX2_X1 U1405 ( .A(\DRAM_mem[6][24] ), .B(n1147), .S(n2208), .Z(n1981) );
  MUX2_X1 U1406 ( .A(\DRAM_mem[6][23] ), .B(n1148), .S(n2208), .Z(n1980) );
  MUX2_X1 U1407 ( .A(\DRAM_mem[6][22] ), .B(n1149), .S(n2208), .Z(n1979) );
  MUX2_X1 U1408 ( .A(\DRAM_mem[6][21] ), .B(n1150), .S(n2208), .Z(n1978) );
  MUX2_X1 U1409 ( .A(\DRAM_mem[6][20] ), .B(n1151), .S(n2208), .Z(n1977) );
  MUX2_X1 U1410 ( .A(\DRAM_mem[6][19] ), .B(n1152), .S(n2208), .Z(n1976) );
  MUX2_X1 U1411 ( .A(\DRAM_mem[6][18] ), .B(n1153), .S(n2208), .Z(n1975) );
  MUX2_X1 U1412 ( .A(\DRAM_mem[6][17] ), .B(n1154), .S(n2208), .Z(n1974) );
  MUX2_X1 U1413 ( .A(\DRAM_mem[6][16] ), .B(n1155), .S(n2208), .Z(n1973) );
  MUX2_X1 U1414 ( .A(\DRAM_mem[6][15] ), .B(n1156), .S(n2208), .Z(n1972) );
  MUX2_X1 U1415 ( .A(\DRAM_mem[6][14] ), .B(n2181), .S(n2208), .Z(n1971) );
  MUX2_X1 U1416 ( .A(\DRAM_mem[6][13] ), .B(n2182), .S(n2208), .Z(n1970) );
  MUX2_X1 U1417 ( .A(\DRAM_mem[6][12] ), .B(n2183), .S(n2208), .Z(n1969) );
  MUX2_X1 U1418 ( .A(\DRAM_mem[6][11] ), .B(n2184), .S(n2208), .Z(n1968) );
  MUX2_X1 U1419 ( .A(\DRAM_mem[6][10] ), .B(n2185), .S(n2208), .Z(n1967) );
  MUX2_X1 U1420 ( .A(\DRAM_mem[6][9] ), .B(n2186), .S(n2208), .Z(n1966) );
  MUX2_X1 U1421 ( .A(\DRAM_mem[6][8] ), .B(n2187), .S(n2208), .Z(n1965) );
  MUX2_X1 U1422 ( .A(\DRAM_mem[6][7] ), .B(n2188), .S(n2208), .Z(n1964) );
  MUX2_X1 U1423 ( .A(\DRAM_mem[6][6] ), .B(n2189), .S(n2208), .Z(n1963) );
  MUX2_X1 U1424 ( .A(\DRAM_mem[6][5] ), .B(n2190), .S(n2208), .Z(n1962) );
  MUX2_X1 U1425 ( .A(\DRAM_mem[6][4] ), .B(n2191), .S(n2208), .Z(n1961) );
  MUX2_X1 U1426 ( .A(\DRAM_mem[6][3] ), .B(n2192), .S(n2208), .Z(n1960) );
  MUX2_X1 U1427 ( .A(\DRAM_mem[6][2] ), .B(n2193), .S(n2208), .Z(n1959) );
  MUX2_X1 U1428 ( .A(\DRAM_mem[6][1] ), .B(n2194), .S(n2208), .Z(n1958) );
  MUX2_X1 U1429 ( .A(\DRAM_mem[6][0] ), .B(n2195), .S(n2208), .Z(n1957) );
  MUX2_X1 U1430 ( .A(\DRAM_mem[7][31] ), .B(n1139), .S(n2210), .Z(n1956) );
  MUX2_X1 U1431 ( .A(\DRAM_mem[7][30] ), .B(n1141), .S(n2210), .Z(n1955) );
  MUX2_X1 U1432 ( .A(\DRAM_mem[7][29] ), .B(n1142), .S(n2210), .Z(n1954) );
  MUX2_X1 U1433 ( .A(\DRAM_mem[7][28] ), .B(n1143), .S(n2210), .Z(n1953) );
  MUX2_X1 U1434 ( .A(\DRAM_mem[7][27] ), .B(n1144), .S(n2210), .Z(n1952) );
  MUX2_X1 U1435 ( .A(\DRAM_mem[7][26] ), .B(n1145), .S(n2210), .Z(n1951) );
  MUX2_X1 U1436 ( .A(\DRAM_mem[7][25] ), .B(n1146), .S(n2210), .Z(n1950) );
  MUX2_X1 U1437 ( .A(\DRAM_mem[7][24] ), .B(n1147), .S(n2210), .Z(n1949) );
  MUX2_X1 U1438 ( .A(\DRAM_mem[7][23] ), .B(n1148), .S(n2210), .Z(n1948) );
  MUX2_X1 U1439 ( .A(\DRAM_mem[7][22] ), .B(n1149), .S(n2210), .Z(n1947) );
  MUX2_X1 U1440 ( .A(\DRAM_mem[7][21] ), .B(n1150), .S(n2210), .Z(n1946) );
  MUX2_X1 U1441 ( .A(\DRAM_mem[7][20] ), .B(n1151), .S(n2210), .Z(n1945) );
  MUX2_X1 U1442 ( .A(\DRAM_mem[7][19] ), .B(n1152), .S(n2210), .Z(n1944) );
  MUX2_X1 U1443 ( .A(\DRAM_mem[7][18] ), .B(n1153), .S(n2210), .Z(n1943) );
  MUX2_X1 U1444 ( .A(\DRAM_mem[7][17] ), .B(n1154), .S(n2210), .Z(n1942) );
  MUX2_X1 U1445 ( .A(\DRAM_mem[7][16] ), .B(n1155), .S(n2210), .Z(n1941) );
  MUX2_X1 U1446 ( .A(\DRAM_mem[7][15] ), .B(n1156), .S(n2210), .Z(n1940) );
  MUX2_X1 U1447 ( .A(\DRAM_mem[7][14] ), .B(n2181), .S(n2210), .Z(n1939) );
  MUX2_X1 U1448 ( .A(\DRAM_mem[7][13] ), .B(n2182), .S(n2210), .Z(n1938) );
  MUX2_X1 U1449 ( .A(\DRAM_mem[7][12] ), .B(n2183), .S(n2210), .Z(n1937) );
  MUX2_X1 U1450 ( .A(\DRAM_mem[7][11] ), .B(n2184), .S(n2210), .Z(n1936) );
  MUX2_X1 U1451 ( .A(\DRAM_mem[7][10] ), .B(n2185), .S(n2210), .Z(n1935) );
  MUX2_X1 U1452 ( .A(\DRAM_mem[7][9] ), .B(n2186), .S(n2210), .Z(n1934) );
  MUX2_X1 U1453 ( .A(\DRAM_mem[7][8] ), .B(n2187), .S(n2210), .Z(n1933) );
  MUX2_X1 U1454 ( .A(\DRAM_mem[7][7] ), .B(n2188), .S(n2210), .Z(n1932) );
  MUX2_X1 U1455 ( .A(\DRAM_mem[7][6] ), .B(n2189), .S(n2210), .Z(n1931) );
  MUX2_X1 U1456 ( .A(\DRAM_mem[7][5] ), .B(n2190), .S(n2210), .Z(n1930) );
  MUX2_X1 U1457 ( .A(\DRAM_mem[7][4] ), .B(n2191), .S(n2210), .Z(n1929) );
  MUX2_X1 U1458 ( .A(\DRAM_mem[7][3] ), .B(n2192), .S(n2210), .Z(n1928) );
  MUX2_X1 U1459 ( .A(\DRAM_mem[7][2] ), .B(n2193), .S(n2210), .Z(n1927) );
  MUX2_X1 U1460 ( .A(\DRAM_mem[7][1] ), .B(n2194), .S(n2210), .Z(n1926) );
  MUX2_X1 U1461 ( .A(\DRAM_mem[7][0] ), .B(n2195), .S(n2210), .Z(n1925) );
  AND3_X1 U1462 ( .A1(n132), .A2(n177), .A3(n2212), .ZN(n2197) );
  MUX2_X1 U1463 ( .A(\DRAM_mem[8][31] ), .B(n1139), .S(n2213), .Z(n1924) );
  MUX2_X1 U1464 ( .A(\DRAM_mem[8][30] ), .B(n1141), .S(n2213), .Z(n1923) );
  MUX2_X1 U1465 ( .A(\DRAM_mem[8][29] ), .B(n1142), .S(n2213), .Z(n1922) );
  MUX2_X1 U1466 ( .A(\DRAM_mem[8][28] ), .B(n1143), .S(n2213), .Z(n1921) );
  MUX2_X1 U1467 ( .A(\DRAM_mem[8][27] ), .B(n1144), .S(n2213), .Z(n1920) );
  MUX2_X1 U1468 ( .A(\DRAM_mem[8][26] ), .B(n1145), .S(n2213), .Z(n1919) );
  MUX2_X1 U1469 ( .A(\DRAM_mem[8][25] ), .B(n1146), .S(n2213), .Z(n1918) );
  MUX2_X1 U1470 ( .A(\DRAM_mem[8][24] ), .B(n1147), .S(n2213), .Z(n1917) );
  MUX2_X1 U1471 ( .A(\DRAM_mem[8][23] ), .B(n1148), .S(n2213), .Z(n1916) );
  MUX2_X1 U1472 ( .A(\DRAM_mem[8][22] ), .B(n1149), .S(n2213), .Z(n1915) );
  MUX2_X1 U1473 ( .A(\DRAM_mem[8][21] ), .B(n1150), .S(n2213), .Z(n1914) );
  MUX2_X1 U1474 ( .A(\DRAM_mem[8][20] ), .B(n1151), .S(n2213), .Z(n1913) );
  MUX2_X1 U1475 ( .A(\DRAM_mem[8][19] ), .B(n1152), .S(n2213), .Z(n1912) );
  MUX2_X1 U1476 ( .A(\DRAM_mem[8][18] ), .B(n1153), .S(n2213), .Z(n1911) );
  MUX2_X1 U1477 ( .A(\DRAM_mem[8][17] ), .B(n1154), .S(n2213), .Z(n1910) );
  MUX2_X1 U1478 ( .A(\DRAM_mem[8][16] ), .B(n1155), .S(n2213), .Z(n1909) );
  MUX2_X1 U1479 ( .A(\DRAM_mem[8][15] ), .B(n1156), .S(n2213), .Z(n1908) );
  MUX2_X1 U1480 ( .A(\DRAM_mem[8][14] ), .B(n2181), .S(n2213), .Z(n1907) );
  MUX2_X1 U1481 ( .A(\DRAM_mem[8][13] ), .B(n2182), .S(n2213), .Z(n1906) );
  MUX2_X1 U1482 ( .A(\DRAM_mem[8][12] ), .B(n2183), .S(n2213), .Z(n1905) );
  MUX2_X1 U1483 ( .A(\DRAM_mem[8][11] ), .B(n2184), .S(n2213), .Z(n1904) );
  MUX2_X1 U1484 ( .A(\DRAM_mem[8][10] ), .B(n2185), .S(n2213), .Z(n1903) );
  MUX2_X1 U1485 ( .A(\DRAM_mem[8][9] ), .B(n2186), .S(n2213), .Z(n1902) );
  MUX2_X1 U1486 ( .A(\DRAM_mem[8][8] ), .B(n2187), .S(n2213), .Z(n1901) );
  MUX2_X1 U1487 ( .A(\DRAM_mem[8][7] ), .B(n2188), .S(n2213), .Z(n1900) );
  MUX2_X1 U1488 ( .A(\DRAM_mem[8][6] ), .B(n2189), .S(n2213), .Z(n1899) );
  MUX2_X1 U1489 ( .A(\DRAM_mem[8][5] ), .B(n2190), .S(n2213), .Z(n1898) );
  MUX2_X1 U1490 ( .A(\DRAM_mem[8][4] ), .B(n2191), .S(n2213), .Z(n1897) );
  MUX2_X1 U1491 ( .A(\DRAM_mem[8][3] ), .B(n2192), .S(n2213), .Z(n1896) );
  MUX2_X1 U1492 ( .A(\DRAM_mem[8][2] ), .B(n2193), .S(n2213), .Z(n1895) );
  MUX2_X1 U1493 ( .A(\DRAM_mem[8][1] ), .B(n2194), .S(n2213), .Z(n1894) );
  MUX2_X1 U1494 ( .A(\DRAM_mem[8][0] ), .B(n2195), .S(n2213), .Z(n1893) );
  MUX2_X1 U1495 ( .A(\DRAM_mem[9][31] ), .B(n1139), .S(n2215), .Z(n1892) );
  MUX2_X1 U1496 ( .A(\DRAM_mem[9][30] ), .B(n1141), .S(n2215), .Z(n1891) );
  MUX2_X1 U1497 ( .A(\DRAM_mem[9][29] ), .B(n1142), .S(n2215), .Z(n1890) );
  MUX2_X1 U1498 ( .A(\DRAM_mem[9][28] ), .B(n1143), .S(n2215), .Z(n1889) );
  MUX2_X1 U1499 ( .A(\DRAM_mem[9][27] ), .B(n1144), .S(n2215), .Z(n1888) );
  MUX2_X1 U1500 ( .A(\DRAM_mem[9][26] ), .B(n1145), .S(n2215), .Z(n1887) );
  MUX2_X1 U1501 ( .A(\DRAM_mem[9][25] ), .B(n1146), .S(n2215), .Z(n1886) );
  MUX2_X1 U1502 ( .A(\DRAM_mem[9][24] ), .B(n1147), .S(n2215), .Z(n1885) );
  MUX2_X1 U1503 ( .A(\DRAM_mem[9][23] ), .B(n1148), .S(n2215), .Z(n1884) );
  MUX2_X1 U1504 ( .A(\DRAM_mem[9][22] ), .B(n1149), .S(n2215), .Z(n1883) );
  MUX2_X1 U1505 ( .A(\DRAM_mem[9][21] ), .B(n1150), .S(n2215), .Z(n1882) );
  MUX2_X1 U1506 ( .A(\DRAM_mem[9][20] ), .B(n1151), .S(n2215), .Z(n1881) );
  MUX2_X1 U1507 ( .A(\DRAM_mem[9][19] ), .B(n1152), .S(n2215), .Z(n1880) );
  MUX2_X1 U1508 ( .A(\DRAM_mem[9][18] ), .B(n1153), .S(n2215), .Z(n1879) );
  MUX2_X1 U1509 ( .A(\DRAM_mem[9][17] ), .B(n1154), .S(n2215), .Z(n1878) );
  MUX2_X1 U1510 ( .A(\DRAM_mem[9][16] ), .B(n1155), .S(n2215), .Z(n1877) );
  MUX2_X1 U1511 ( .A(\DRAM_mem[9][15] ), .B(n1156), .S(n2215), .Z(n1876) );
  MUX2_X1 U1512 ( .A(\DRAM_mem[9][14] ), .B(n2181), .S(n2215), .Z(n1875) );
  MUX2_X1 U1513 ( .A(\DRAM_mem[9][13] ), .B(n2182), .S(n2215), .Z(n1874) );
  MUX2_X1 U1514 ( .A(\DRAM_mem[9][12] ), .B(n2183), .S(n2215), .Z(n1873) );
  MUX2_X1 U1515 ( .A(\DRAM_mem[9][11] ), .B(n2184), .S(n2215), .Z(n1872) );
  MUX2_X1 U1516 ( .A(\DRAM_mem[9][10] ), .B(n2185), .S(n2215), .Z(n1871) );
  MUX2_X1 U1517 ( .A(\DRAM_mem[9][9] ), .B(n2186), .S(n2215), .Z(n1870) );
  MUX2_X1 U1518 ( .A(\DRAM_mem[9][8] ), .B(n2187), .S(n2215), .Z(n1869) );
  MUX2_X1 U1519 ( .A(\DRAM_mem[9][7] ), .B(n2188), .S(n2215), .Z(n1868) );
  MUX2_X1 U1520 ( .A(\DRAM_mem[9][6] ), .B(n2189), .S(n2215), .Z(n1867) );
  MUX2_X1 U1521 ( .A(\DRAM_mem[9][5] ), .B(n2190), .S(n2215), .Z(n1866) );
  MUX2_X1 U1522 ( .A(\DRAM_mem[9][4] ), .B(n2191), .S(n2215), .Z(n1865) );
  MUX2_X1 U1523 ( .A(\DRAM_mem[9][3] ), .B(n2192), .S(n2215), .Z(n1864) );
  MUX2_X1 U1524 ( .A(\DRAM_mem[9][2] ), .B(n2193), .S(n2215), .Z(n1863) );
  MUX2_X1 U1525 ( .A(\DRAM_mem[9][1] ), .B(n2194), .S(n2215), .Z(n1862) );
  MUX2_X1 U1526 ( .A(\DRAM_mem[9][0] ), .B(n2195), .S(n2215), .Z(n1861) );
  MUX2_X1 U1527 ( .A(\DRAM_mem[10][31] ), .B(n1139), .S(n2216), .Z(n1860) );
  MUX2_X1 U1528 ( .A(\DRAM_mem[10][30] ), .B(n1141), .S(n2216), .Z(n1859) );
  MUX2_X1 U1529 ( .A(\DRAM_mem[10][29] ), .B(n1142), .S(n2216), .Z(n1858) );
  MUX2_X1 U1530 ( .A(\DRAM_mem[10][28] ), .B(n1143), .S(n2216), .Z(n1857) );
  MUX2_X1 U1531 ( .A(\DRAM_mem[10][27] ), .B(n1144), .S(n2216), .Z(n1856) );
  MUX2_X1 U1532 ( .A(\DRAM_mem[10][26] ), .B(n1145), .S(n2216), .Z(n1855) );
  MUX2_X1 U1533 ( .A(\DRAM_mem[10][25] ), .B(n1146), .S(n2216), .Z(n1854) );
  MUX2_X1 U1534 ( .A(\DRAM_mem[10][24] ), .B(n1147), .S(n2216), .Z(n1853) );
  MUX2_X1 U1535 ( .A(\DRAM_mem[10][23] ), .B(n1148), .S(n2216), .Z(n1852) );
  MUX2_X1 U1536 ( .A(\DRAM_mem[10][22] ), .B(n1149), .S(n2216), .Z(n1851) );
  MUX2_X1 U1537 ( .A(\DRAM_mem[10][21] ), .B(n1150), .S(n2216), .Z(n1850) );
  MUX2_X1 U1538 ( .A(\DRAM_mem[10][20] ), .B(n1151), .S(n2216), .Z(n1849) );
  MUX2_X1 U1539 ( .A(\DRAM_mem[10][19] ), .B(n1152), .S(n2216), .Z(n1848) );
  MUX2_X1 U1540 ( .A(\DRAM_mem[10][18] ), .B(n1153), .S(n2216), .Z(n1847) );
  MUX2_X1 U1541 ( .A(\DRAM_mem[10][17] ), .B(n1154), .S(n2216), .Z(n1846) );
  MUX2_X1 U1542 ( .A(\DRAM_mem[10][16] ), .B(n1155), .S(n2216), .Z(n1845) );
  MUX2_X1 U1543 ( .A(\DRAM_mem[10][15] ), .B(n1156), .S(n2216), .Z(n1844) );
  MUX2_X1 U1544 ( .A(\DRAM_mem[10][14] ), .B(n2181), .S(n2216), .Z(n1843) );
  MUX2_X1 U1545 ( .A(\DRAM_mem[10][13] ), .B(n2182), .S(n2216), .Z(n1842) );
  MUX2_X1 U1546 ( .A(\DRAM_mem[10][12] ), .B(n2183), .S(n2216), .Z(n1841) );
  MUX2_X1 U1547 ( .A(\DRAM_mem[10][11] ), .B(n2184), .S(n2216), .Z(n1840) );
  MUX2_X1 U1548 ( .A(\DRAM_mem[10][10] ), .B(n2185), .S(n2216), .Z(n1839) );
  MUX2_X1 U1549 ( .A(\DRAM_mem[10][9] ), .B(n2186), .S(n2216), .Z(n1838) );
  MUX2_X1 U1550 ( .A(\DRAM_mem[10][8] ), .B(n2187), .S(n2216), .Z(n1837) );
  MUX2_X1 U1551 ( .A(\DRAM_mem[10][7] ), .B(n2188), .S(n2216), .Z(n1836) );
  MUX2_X1 U1552 ( .A(\DRAM_mem[10][6] ), .B(n2189), .S(n2216), .Z(n1835) );
  MUX2_X1 U1553 ( .A(\DRAM_mem[10][5] ), .B(n2190), .S(n2216), .Z(n1834) );
  MUX2_X1 U1554 ( .A(\DRAM_mem[10][4] ), .B(n2191), .S(n2216), .Z(n1833) );
  MUX2_X1 U1555 ( .A(\DRAM_mem[10][3] ), .B(n2192), .S(n2216), .Z(n1832) );
  MUX2_X1 U1556 ( .A(\DRAM_mem[10][2] ), .B(n2193), .S(n2216), .Z(n1831) );
  MUX2_X1 U1557 ( .A(\DRAM_mem[10][1] ), .B(n2194), .S(n2216), .Z(n1830) );
  MUX2_X1 U1558 ( .A(\DRAM_mem[10][0] ), .B(n2195), .S(n2216), .Z(n1829) );
  MUX2_X1 U1559 ( .A(\DRAM_mem[11][31] ), .B(n1139), .S(n2217), .Z(n1828) );
  MUX2_X1 U1560 ( .A(\DRAM_mem[11][30] ), .B(n1141), .S(n2217), .Z(n1827) );
  MUX2_X1 U1561 ( .A(\DRAM_mem[11][29] ), .B(n1142), .S(n2217), .Z(n1826) );
  MUX2_X1 U1562 ( .A(\DRAM_mem[11][28] ), .B(n1143), .S(n2217), .Z(n1825) );
  MUX2_X1 U1563 ( .A(\DRAM_mem[11][27] ), .B(n1144), .S(n2217), .Z(n1824) );
  MUX2_X1 U1564 ( .A(\DRAM_mem[11][26] ), .B(n1145), .S(n2217), .Z(n1823) );
  MUX2_X1 U1565 ( .A(\DRAM_mem[11][25] ), .B(n1146), .S(n2217), .Z(n1822) );
  MUX2_X1 U1566 ( .A(\DRAM_mem[11][24] ), .B(n1147), .S(n2217), .Z(n1821) );
  MUX2_X1 U1567 ( .A(\DRAM_mem[11][23] ), .B(n1148), .S(n2217), .Z(n1820) );
  MUX2_X1 U1568 ( .A(\DRAM_mem[11][22] ), .B(n1149), .S(n2217), .Z(n1819) );
  MUX2_X1 U1569 ( .A(\DRAM_mem[11][21] ), .B(n1150), .S(n2217), .Z(n1818) );
  MUX2_X1 U1570 ( .A(\DRAM_mem[11][20] ), .B(n1151), .S(n2217), .Z(n1817) );
  MUX2_X1 U1571 ( .A(\DRAM_mem[11][19] ), .B(n1152), .S(n2217), .Z(n1816) );
  MUX2_X1 U1572 ( .A(\DRAM_mem[11][18] ), .B(n1153), .S(n2217), .Z(n1815) );
  MUX2_X1 U1573 ( .A(\DRAM_mem[11][17] ), .B(n1154), .S(n2217), .Z(n1814) );
  MUX2_X1 U1574 ( .A(\DRAM_mem[11][16] ), .B(n1155), .S(n2217), .Z(n1813) );
  MUX2_X1 U1575 ( .A(\DRAM_mem[11][15] ), .B(n1156), .S(n2217), .Z(n1812) );
  MUX2_X1 U1576 ( .A(\DRAM_mem[11][14] ), .B(n2181), .S(n2217), .Z(n1811) );
  MUX2_X1 U1577 ( .A(\DRAM_mem[11][13] ), .B(n2182), .S(n2217), .Z(n1810) );
  MUX2_X1 U1578 ( .A(\DRAM_mem[11][12] ), .B(n2183), .S(n2217), .Z(n1809) );
  MUX2_X1 U1579 ( .A(\DRAM_mem[11][11] ), .B(n2184), .S(n2217), .Z(n1808) );
  MUX2_X1 U1580 ( .A(\DRAM_mem[11][10] ), .B(n2185), .S(n2217), .Z(n1807) );
  MUX2_X1 U1581 ( .A(\DRAM_mem[11][9] ), .B(n2186), .S(n2217), .Z(n1806) );
  MUX2_X1 U1582 ( .A(\DRAM_mem[11][8] ), .B(n2187), .S(n2217), .Z(n1805) );
  MUX2_X1 U1583 ( .A(\DRAM_mem[11][7] ), .B(n2188), .S(n2217), .Z(n1804) );
  MUX2_X1 U1584 ( .A(\DRAM_mem[11][6] ), .B(n2189), .S(n2217), .Z(n1803) );
  MUX2_X1 U1585 ( .A(\DRAM_mem[11][5] ), .B(n2190), .S(n2217), .Z(n1802) );
  MUX2_X1 U1586 ( .A(\DRAM_mem[11][4] ), .B(n2191), .S(n2217), .Z(n1801) );
  MUX2_X1 U1587 ( .A(\DRAM_mem[11][3] ), .B(n2192), .S(n2217), .Z(n1800) );
  MUX2_X1 U1588 ( .A(\DRAM_mem[11][2] ), .B(n2193), .S(n2217), .Z(n1799) );
  MUX2_X1 U1589 ( .A(\DRAM_mem[11][1] ), .B(n2194), .S(n2217), .Z(n1798) );
  MUX2_X1 U1590 ( .A(\DRAM_mem[11][0] ), .B(n2195), .S(n2217), .Z(n1797) );
  MUX2_X1 U1591 ( .A(\DRAM_mem[12][31] ), .B(n1139), .S(n2218), .Z(n1796) );
  MUX2_X1 U1592 ( .A(\DRAM_mem[12][30] ), .B(n1141), .S(n2218), .Z(n1795) );
  MUX2_X1 U1593 ( .A(\DRAM_mem[12][29] ), .B(n1142), .S(n2218), .Z(n1794) );
  MUX2_X1 U1594 ( .A(\DRAM_mem[12][28] ), .B(n1143), .S(n2218), .Z(n1793) );
  MUX2_X1 U1595 ( .A(\DRAM_mem[12][27] ), .B(n1144), .S(n2218), .Z(n1792) );
  MUX2_X1 U1596 ( .A(\DRAM_mem[12][26] ), .B(n1145), .S(n2218), .Z(n1791) );
  MUX2_X1 U1597 ( .A(\DRAM_mem[12][25] ), .B(n1146), .S(n2218), .Z(n1790) );
  MUX2_X1 U1598 ( .A(\DRAM_mem[12][24] ), .B(n1147), .S(n2218), .Z(n1789) );
  MUX2_X1 U1599 ( .A(\DRAM_mem[12][23] ), .B(n1148), .S(n2218), .Z(n1788) );
  MUX2_X1 U1600 ( .A(\DRAM_mem[12][22] ), .B(n1149), .S(n2218), .Z(n1787) );
  MUX2_X1 U1601 ( .A(\DRAM_mem[12][21] ), .B(n1150), .S(n2218), .Z(n1786) );
  MUX2_X1 U1602 ( .A(\DRAM_mem[12][20] ), .B(n1151), .S(n2218), .Z(n1785) );
  MUX2_X1 U1603 ( .A(\DRAM_mem[12][19] ), .B(n1152), .S(n2218), .Z(n1784) );
  MUX2_X1 U1604 ( .A(\DRAM_mem[12][18] ), .B(n1153), .S(n2218), .Z(n1783) );
  MUX2_X1 U1605 ( .A(\DRAM_mem[12][17] ), .B(n1154), .S(n2218), .Z(n1782) );
  MUX2_X1 U1606 ( .A(\DRAM_mem[12][16] ), .B(n1155), .S(n2218), .Z(n1781) );
  MUX2_X1 U1607 ( .A(\DRAM_mem[12][15] ), .B(n1156), .S(n2218), .Z(n1780) );
  MUX2_X1 U1608 ( .A(\DRAM_mem[12][14] ), .B(n2181), .S(n2218), .Z(n1779) );
  MUX2_X1 U1609 ( .A(\DRAM_mem[12][13] ), .B(n2182), .S(n2218), .Z(n1778) );
  MUX2_X1 U1610 ( .A(\DRAM_mem[12][12] ), .B(n2183), .S(n2218), .Z(n1777) );
  MUX2_X1 U1611 ( .A(\DRAM_mem[12][11] ), .B(n2184), .S(n2218), .Z(n1776) );
  MUX2_X1 U1612 ( .A(\DRAM_mem[12][10] ), .B(n2185), .S(n2218), .Z(n1775) );
  MUX2_X1 U1613 ( .A(\DRAM_mem[12][9] ), .B(n2186), .S(n2218), .Z(n1774) );
  MUX2_X1 U1614 ( .A(\DRAM_mem[12][8] ), .B(n2187), .S(n2218), .Z(n1773) );
  MUX2_X1 U1615 ( .A(\DRAM_mem[12][7] ), .B(n2188), .S(n2218), .Z(n1772) );
  MUX2_X1 U1616 ( .A(\DRAM_mem[12][6] ), .B(n2189), .S(n2218), .Z(n1771) );
  MUX2_X1 U1617 ( .A(\DRAM_mem[12][5] ), .B(n2190), .S(n2218), .Z(n1770) );
  MUX2_X1 U1618 ( .A(\DRAM_mem[12][4] ), .B(n2191), .S(n2218), .Z(n1769) );
  MUX2_X1 U1619 ( .A(\DRAM_mem[12][3] ), .B(n2192), .S(n2218), .Z(n1768) );
  MUX2_X1 U1620 ( .A(\DRAM_mem[12][2] ), .B(n2193), .S(n2218), .Z(n1767) );
  MUX2_X1 U1621 ( .A(\DRAM_mem[12][1] ), .B(n2194), .S(n2218), .Z(n1766) );
  MUX2_X1 U1622 ( .A(\DRAM_mem[12][0] ), .B(n2195), .S(n2218), .Z(n1765) );
  MUX2_X1 U1623 ( .A(\DRAM_mem[13][31] ), .B(n1139), .S(n2219), .Z(n1764) );
  MUX2_X1 U1624 ( .A(\DRAM_mem[13][30] ), .B(n1141), .S(n2219), .Z(n1763) );
  MUX2_X1 U1625 ( .A(\DRAM_mem[13][29] ), .B(n1142), .S(n2219), .Z(n1762) );
  MUX2_X1 U1626 ( .A(\DRAM_mem[13][28] ), .B(n1143), .S(n2219), .Z(n1761) );
  MUX2_X1 U1627 ( .A(\DRAM_mem[13][27] ), .B(n1144), .S(n2219), .Z(n1760) );
  MUX2_X1 U1628 ( .A(\DRAM_mem[13][26] ), .B(n1145), .S(n2219), .Z(n1759) );
  MUX2_X1 U1629 ( .A(\DRAM_mem[13][25] ), .B(n1146), .S(n2219), .Z(n1758) );
  MUX2_X1 U1630 ( .A(\DRAM_mem[13][24] ), .B(n1147), .S(n2219), .Z(n1757) );
  MUX2_X1 U1631 ( .A(\DRAM_mem[13][23] ), .B(n1148), .S(n2219), .Z(n1756) );
  MUX2_X1 U1632 ( .A(\DRAM_mem[13][22] ), .B(n1149), .S(n2219), .Z(n1755) );
  MUX2_X1 U1633 ( .A(\DRAM_mem[13][21] ), .B(n1150), .S(n2219), .Z(n1754) );
  MUX2_X1 U1634 ( .A(\DRAM_mem[13][20] ), .B(n1151), .S(n2219), .Z(n1753) );
  MUX2_X1 U1635 ( .A(\DRAM_mem[13][19] ), .B(n1152), .S(n2219), .Z(n1752) );
  MUX2_X1 U1636 ( .A(\DRAM_mem[13][18] ), .B(n1153), .S(n2219), .Z(n1751) );
  MUX2_X1 U1637 ( .A(\DRAM_mem[13][17] ), .B(n1154), .S(n2219), .Z(n1750) );
  MUX2_X1 U1638 ( .A(\DRAM_mem[13][16] ), .B(n1155), .S(n2219), .Z(n1749) );
  MUX2_X1 U1639 ( .A(\DRAM_mem[13][15] ), .B(n1156), .S(n2219), .Z(n1748) );
  MUX2_X1 U1640 ( .A(\DRAM_mem[13][14] ), .B(n2181), .S(n2219), .Z(n1747) );
  MUX2_X1 U1641 ( .A(\DRAM_mem[13][13] ), .B(n2182), .S(n2219), .Z(n1746) );
  MUX2_X1 U1642 ( .A(\DRAM_mem[13][12] ), .B(n2183), .S(n2219), .Z(n1745) );
  MUX2_X1 U1643 ( .A(\DRAM_mem[13][11] ), .B(n2184), .S(n2219), .Z(n1744) );
  MUX2_X1 U1644 ( .A(\DRAM_mem[13][10] ), .B(n2185), .S(n2219), .Z(n1743) );
  MUX2_X1 U1645 ( .A(\DRAM_mem[13][9] ), .B(n2186), .S(n2219), .Z(n1742) );
  MUX2_X1 U1646 ( .A(\DRAM_mem[13][8] ), .B(n2187), .S(n2219), .Z(n1741) );
  MUX2_X1 U1647 ( .A(\DRAM_mem[13][7] ), .B(n2188), .S(n2219), .Z(n1740) );
  MUX2_X1 U1648 ( .A(\DRAM_mem[13][6] ), .B(n2189), .S(n2219), .Z(n1739) );
  MUX2_X1 U1649 ( .A(\DRAM_mem[13][5] ), .B(n2190), .S(n2219), .Z(n1738) );
  MUX2_X1 U1650 ( .A(\DRAM_mem[13][4] ), .B(n2191), .S(n2219), .Z(n1737) );
  MUX2_X1 U1651 ( .A(\DRAM_mem[13][3] ), .B(n2192), .S(n2219), .Z(n1736) );
  MUX2_X1 U1652 ( .A(\DRAM_mem[13][2] ), .B(n2193), .S(n2219), .Z(n1735) );
  MUX2_X1 U1653 ( .A(\DRAM_mem[13][1] ), .B(n2194), .S(n2219), .Z(n1734) );
  MUX2_X1 U1654 ( .A(\DRAM_mem[13][0] ), .B(n2195), .S(n2219), .Z(n1733) );
  MUX2_X1 U1655 ( .A(\DRAM_mem[14][31] ), .B(n1139), .S(n2220), .Z(n1732) );
  MUX2_X1 U1656 ( .A(\DRAM_mem[14][30] ), .B(n1141), .S(n2220), .Z(n1731) );
  MUX2_X1 U1657 ( .A(\DRAM_mem[14][29] ), .B(n1142), .S(n2220), .Z(n1730) );
  MUX2_X1 U1658 ( .A(\DRAM_mem[14][28] ), .B(n1143), .S(n2220), .Z(n1729) );
  MUX2_X1 U1659 ( .A(\DRAM_mem[14][27] ), .B(n1144), .S(n2220), .Z(n1728) );
  MUX2_X1 U1660 ( .A(\DRAM_mem[14][26] ), .B(n1145), .S(n2220), .Z(n1727) );
  MUX2_X1 U1661 ( .A(\DRAM_mem[14][25] ), .B(n1146), .S(n2220), .Z(n1726) );
  MUX2_X1 U1662 ( .A(\DRAM_mem[14][24] ), .B(n1147), .S(n2220), .Z(n1725) );
  MUX2_X1 U1663 ( .A(\DRAM_mem[14][23] ), .B(n1148), .S(n2220), .Z(n1724) );
  MUX2_X1 U1664 ( .A(\DRAM_mem[14][22] ), .B(n1149), .S(n2220), .Z(n1723) );
  MUX2_X1 U1665 ( .A(\DRAM_mem[14][21] ), .B(n1150), .S(n2220), .Z(n1722) );
  MUX2_X1 U1666 ( .A(\DRAM_mem[14][20] ), .B(n1151), .S(n2220), .Z(n1721) );
  MUX2_X1 U1667 ( .A(\DRAM_mem[14][19] ), .B(n1152), .S(n2220), .Z(n1720) );
  MUX2_X1 U1668 ( .A(\DRAM_mem[14][18] ), .B(n1153), .S(n2220), .Z(n1719) );
  MUX2_X1 U1669 ( .A(\DRAM_mem[14][17] ), .B(n1154), .S(n2220), .Z(n1718) );
  MUX2_X1 U1670 ( .A(\DRAM_mem[14][16] ), .B(n1155), .S(n2220), .Z(n1717) );
  MUX2_X1 U1671 ( .A(\DRAM_mem[14][15] ), .B(n1156), .S(n2220), .Z(n1716) );
  MUX2_X1 U1672 ( .A(\DRAM_mem[14][14] ), .B(n2181), .S(n2220), .Z(n1715) );
  MUX2_X1 U1673 ( .A(\DRAM_mem[14][13] ), .B(n2182), .S(n2220), .Z(n1714) );
  MUX2_X1 U1674 ( .A(\DRAM_mem[14][12] ), .B(n2183), .S(n2220), .Z(n1713) );
  MUX2_X1 U1675 ( .A(\DRAM_mem[14][11] ), .B(n2184), .S(n2220), .Z(n1712) );
  MUX2_X1 U1676 ( .A(\DRAM_mem[14][10] ), .B(n2185), .S(n2220), .Z(n1711) );
  MUX2_X1 U1677 ( .A(\DRAM_mem[14][9] ), .B(n2186), .S(n2220), .Z(n1710) );
  MUX2_X1 U1678 ( .A(\DRAM_mem[14][8] ), .B(n2187), .S(n2220), .Z(n1709) );
  MUX2_X1 U1679 ( .A(\DRAM_mem[14][7] ), .B(n2188), .S(n2220), .Z(n1708) );
  MUX2_X1 U1680 ( .A(\DRAM_mem[14][6] ), .B(n2189), .S(n2220), .Z(n1707) );
  MUX2_X1 U1681 ( .A(\DRAM_mem[14][5] ), .B(n2190), .S(n2220), .Z(n1706) );
  MUX2_X1 U1682 ( .A(\DRAM_mem[14][4] ), .B(n2191), .S(n2220), .Z(n1705) );
  MUX2_X1 U1683 ( .A(\DRAM_mem[14][3] ), .B(n2192), .S(n2220), .Z(n1704) );
  MUX2_X1 U1684 ( .A(\DRAM_mem[14][2] ), .B(n2193), .S(n2220), .Z(n1703) );
  MUX2_X1 U1685 ( .A(\DRAM_mem[14][1] ), .B(n2194), .S(n2220), .Z(n1702) );
  MUX2_X1 U1686 ( .A(\DRAM_mem[14][0] ), .B(n2195), .S(n2220), .Z(n1701) );
  MUX2_X1 U1687 ( .A(\DRAM_mem[15][31] ), .B(n1139), .S(n2221), .Z(n1700) );
  MUX2_X1 U1688 ( .A(\DRAM_mem[15][30] ), .B(n1141), .S(n2221), .Z(n1699) );
  MUX2_X1 U1689 ( .A(\DRAM_mem[15][29] ), .B(n1142), .S(n2221), .Z(n1698) );
  MUX2_X1 U1690 ( .A(\DRAM_mem[15][28] ), .B(n1143), .S(n2221), .Z(n1697) );
  MUX2_X1 U1691 ( .A(\DRAM_mem[15][27] ), .B(n1144), .S(n2221), .Z(n1696) );
  MUX2_X1 U1692 ( .A(\DRAM_mem[15][26] ), .B(n1145), .S(n2221), .Z(n1695) );
  MUX2_X1 U1693 ( .A(\DRAM_mem[15][25] ), .B(n1146), .S(n2221), .Z(n1694) );
  MUX2_X1 U1694 ( .A(\DRAM_mem[15][24] ), .B(n1147), .S(n2221), .Z(n1693) );
  MUX2_X1 U1695 ( .A(\DRAM_mem[15][23] ), .B(n1148), .S(n2221), .Z(n1692) );
  MUX2_X1 U1696 ( .A(\DRAM_mem[15][22] ), .B(n1149), .S(n2221), .Z(n1691) );
  MUX2_X1 U1697 ( .A(\DRAM_mem[15][21] ), .B(n1150), .S(n2221), .Z(n1690) );
  MUX2_X1 U1698 ( .A(\DRAM_mem[15][20] ), .B(n1151), .S(n2221), .Z(n1689) );
  MUX2_X1 U1699 ( .A(\DRAM_mem[15][19] ), .B(n1152), .S(n2221), .Z(n1688) );
  MUX2_X1 U1700 ( .A(\DRAM_mem[15][18] ), .B(n1153), .S(n2221), .Z(n1687) );
  MUX2_X1 U1701 ( .A(\DRAM_mem[15][17] ), .B(n1154), .S(n2221), .Z(n1686) );
  MUX2_X1 U1702 ( .A(\DRAM_mem[15][16] ), .B(n1155), .S(n2221), .Z(n1685) );
  MUX2_X1 U1703 ( .A(\DRAM_mem[15][15] ), .B(n1156), .S(n2221), .Z(n1684) );
  MUX2_X1 U1704 ( .A(\DRAM_mem[15][14] ), .B(n2181), .S(n2221), .Z(n1683) );
  MUX2_X1 U1705 ( .A(\DRAM_mem[15][13] ), .B(n2182), .S(n2221), .Z(n1682) );
  MUX2_X1 U1706 ( .A(\DRAM_mem[15][12] ), .B(n2183), .S(n2221), .Z(n1681) );
  MUX2_X1 U1707 ( .A(\DRAM_mem[15][11] ), .B(n2184), .S(n2221), .Z(n1680) );
  MUX2_X1 U1708 ( .A(\DRAM_mem[15][10] ), .B(n2185), .S(n2221), .Z(n1679) );
  MUX2_X1 U1709 ( .A(\DRAM_mem[15][9] ), .B(n2186), .S(n2221), .Z(n1678) );
  MUX2_X1 U1710 ( .A(\DRAM_mem[15][8] ), .B(n2187), .S(n2221), .Z(n1677) );
  MUX2_X1 U1711 ( .A(\DRAM_mem[15][7] ), .B(n2188), .S(n2221), .Z(n1676) );
  MUX2_X1 U1712 ( .A(\DRAM_mem[15][6] ), .B(n2189), .S(n2221), .Z(n1675) );
  MUX2_X1 U1713 ( .A(\DRAM_mem[15][5] ), .B(n2190), .S(n2221), .Z(n1674) );
  MUX2_X1 U1714 ( .A(\DRAM_mem[15][4] ), .B(n2191), .S(n2221), .Z(n1673) );
  MUX2_X1 U1715 ( .A(\DRAM_mem[15][3] ), .B(n2192), .S(n2221), .Z(n1672) );
  MUX2_X1 U1716 ( .A(\DRAM_mem[15][2] ), .B(n2193), .S(n2221), .Z(n1671) );
  MUX2_X1 U1717 ( .A(\DRAM_mem[15][1] ), .B(n2194), .S(n2221), .Z(n1670) );
  MUX2_X1 U1718 ( .A(\DRAM_mem[15][0] ), .B(n2195), .S(n2221), .Z(n1669) );
  AND3_X1 U1719 ( .A1(n2212), .A2(n177), .A3(Addr[3]), .ZN(n2214) );
  MUX2_X1 U1720 ( .A(\DRAM_mem[16][31] ), .B(n1139), .S(n2222), .Z(n1668) );
  MUX2_X1 U1721 ( .A(\DRAM_mem[16][30] ), .B(n1141), .S(n2222), .Z(n1667) );
  MUX2_X1 U1722 ( .A(\DRAM_mem[16][29] ), .B(n1142), .S(n2222), .Z(n1666) );
  MUX2_X1 U1723 ( .A(\DRAM_mem[16][28] ), .B(n1143), .S(n2222), .Z(n1665) );
  MUX2_X1 U1724 ( .A(\DRAM_mem[16][27] ), .B(n1144), .S(n2222), .Z(n1664) );
  MUX2_X1 U1725 ( .A(\DRAM_mem[16][26] ), .B(n1145), .S(n2222), .Z(n1663) );
  MUX2_X1 U1726 ( .A(\DRAM_mem[16][25] ), .B(n1146), .S(n2222), .Z(n1662) );
  MUX2_X1 U1727 ( .A(\DRAM_mem[16][24] ), .B(n1147), .S(n2222), .Z(n1661) );
  MUX2_X1 U1728 ( .A(\DRAM_mem[16][23] ), .B(n1148), .S(n2222), .Z(n1660) );
  MUX2_X1 U1729 ( .A(\DRAM_mem[16][22] ), .B(n1149), .S(n2222), .Z(n1659) );
  MUX2_X1 U1730 ( .A(\DRAM_mem[16][21] ), .B(n1150), .S(n2222), .Z(n1658) );
  MUX2_X1 U1731 ( .A(\DRAM_mem[16][20] ), .B(n1151), .S(n2222), .Z(n1657) );
  MUX2_X1 U1732 ( .A(\DRAM_mem[16][19] ), .B(n1152), .S(n2222), .Z(n1656) );
  MUX2_X1 U1733 ( .A(\DRAM_mem[16][18] ), .B(n1153), .S(n2222), .Z(n1655) );
  MUX2_X1 U1734 ( .A(\DRAM_mem[16][17] ), .B(n1154), .S(n2222), .Z(n1654) );
  MUX2_X1 U1735 ( .A(\DRAM_mem[16][16] ), .B(n1155), .S(n2222), .Z(n1653) );
  MUX2_X1 U1736 ( .A(\DRAM_mem[16][15] ), .B(n1156), .S(n2222), .Z(n1652) );
  MUX2_X1 U1737 ( .A(\DRAM_mem[16][14] ), .B(n2181), .S(n2222), .Z(n1651) );
  MUX2_X1 U1738 ( .A(\DRAM_mem[16][13] ), .B(n2182), .S(n2222), .Z(n1650) );
  MUX2_X1 U1739 ( .A(\DRAM_mem[16][12] ), .B(n2183), .S(n2222), .Z(n1649) );
  MUX2_X1 U1740 ( .A(\DRAM_mem[16][11] ), .B(n2184), .S(n2222), .Z(n1648) );
  MUX2_X1 U1741 ( .A(\DRAM_mem[16][10] ), .B(n2185), .S(n2222), .Z(n1647) );
  MUX2_X1 U1742 ( .A(\DRAM_mem[16][9] ), .B(n2186), .S(n2222), .Z(n1646) );
  MUX2_X1 U1743 ( .A(\DRAM_mem[16][8] ), .B(n2187), .S(n2222), .Z(n1645) );
  MUX2_X1 U1744 ( .A(\DRAM_mem[16][7] ), .B(n2188), .S(n2222), .Z(n1644) );
  MUX2_X1 U1745 ( .A(\DRAM_mem[16][6] ), .B(n2189), .S(n2222), .Z(n1643) );
  MUX2_X1 U1746 ( .A(\DRAM_mem[16][5] ), .B(n2190), .S(n2222), .Z(n1642) );
  MUX2_X1 U1747 ( .A(\DRAM_mem[16][4] ), .B(n2191), .S(n2222), .Z(n1641) );
  MUX2_X1 U1748 ( .A(\DRAM_mem[16][3] ), .B(n2192), .S(n2222), .Z(n1640) );
  MUX2_X1 U1749 ( .A(\DRAM_mem[16][2] ), .B(n2193), .S(n2222), .Z(n1639) );
  MUX2_X1 U1750 ( .A(\DRAM_mem[16][1] ), .B(n2194), .S(n2222), .Z(n1638) );
  MUX2_X1 U1751 ( .A(\DRAM_mem[16][0] ), .B(n2195), .S(n2222), .Z(n1637) );
  MUX2_X1 U1752 ( .A(\DRAM_mem[17][31] ), .B(n1139), .S(n2224), .Z(n1636) );
  MUX2_X1 U1753 ( .A(\DRAM_mem[17][30] ), .B(n1141), .S(n2224), .Z(n1635) );
  MUX2_X1 U1754 ( .A(\DRAM_mem[17][29] ), .B(n1142), .S(n2224), .Z(n1634) );
  MUX2_X1 U1755 ( .A(\DRAM_mem[17][28] ), .B(n1143), .S(n2224), .Z(n1633) );
  MUX2_X1 U1756 ( .A(\DRAM_mem[17][27] ), .B(n1144), .S(n2224), .Z(n1632) );
  MUX2_X1 U1757 ( .A(\DRAM_mem[17][26] ), .B(n1145), .S(n2224), .Z(n1631) );
  MUX2_X1 U1758 ( .A(\DRAM_mem[17][25] ), .B(n1146), .S(n2224), .Z(n1630) );
  MUX2_X1 U1759 ( .A(\DRAM_mem[17][24] ), .B(n1147), .S(n2224), .Z(n1629) );
  MUX2_X1 U1760 ( .A(\DRAM_mem[17][23] ), .B(n1148), .S(n2224), .Z(n1628) );
  MUX2_X1 U1761 ( .A(\DRAM_mem[17][22] ), .B(n1149), .S(n2224), .Z(n1627) );
  MUX2_X1 U1762 ( .A(\DRAM_mem[17][21] ), .B(n1150), .S(n2224), .Z(n1626) );
  MUX2_X1 U1763 ( .A(\DRAM_mem[17][20] ), .B(n1151), .S(n2224), .Z(n1625) );
  MUX2_X1 U1764 ( .A(\DRAM_mem[17][19] ), .B(n1152), .S(n2224), .Z(n1624) );
  MUX2_X1 U1765 ( .A(\DRAM_mem[17][18] ), .B(n1153), .S(n2224), .Z(n1623) );
  MUX2_X1 U1766 ( .A(\DRAM_mem[17][17] ), .B(n1154), .S(n2224), .Z(n1622) );
  MUX2_X1 U1767 ( .A(\DRAM_mem[17][16] ), .B(n1155), .S(n2224), .Z(n1621) );
  MUX2_X1 U1768 ( .A(\DRAM_mem[17][15] ), .B(n1156), .S(n2224), .Z(n1620) );
  MUX2_X1 U1769 ( .A(\DRAM_mem[17][14] ), .B(n2181), .S(n2224), .Z(n1619) );
  MUX2_X1 U1770 ( .A(\DRAM_mem[17][13] ), .B(n2182), .S(n2224), .Z(n1618) );
  MUX2_X1 U1771 ( .A(\DRAM_mem[17][12] ), .B(n2183), .S(n2224), .Z(n1617) );
  MUX2_X1 U1772 ( .A(\DRAM_mem[17][11] ), .B(n2184), .S(n2224), .Z(n1616) );
  MUX2_X1 U1773 ( .A(\DRAM_mem[17][10] ), .B(n2185), .S(n2224), .Z(n1615) );
  MUX2_X1 U1774 ( .A(\DRAM_mem[17][9] ), .B(n2186), .S(n2224), .Z(n1614) );
  MUX2_X1 U1775 ( .A(\DRAM_mem[17][8] ), .B(n2187), .S(n2224), .Z(n1613) );
  MUX2_X1 U1776 ( .A(\DRAM_mem[17][7] ), .B(n2188), .S(n2224), .Z(n1612) );
  MUX2_X1 U1777 ( .A(\DRAM_mem[17][6] ), .B(n2189), .S(n2224), .Z(n1611) );
  MUX2_X1 U1778 ( .A(\DRAM_mem[17][5] ), .B(n2190), .S(n2224), .Z(n1610) );
  MUX2_X1 U1779 ( .A(\DRAM_mem[17][4] ), .B(n2191), .S(n2224), .Z(n1609) );
  MUX2_X1 U1780 ( .A(\DRAM_mem[17][3] ), .B(n2192), .S(n2224), .Z(n1608) );
  MUX2_X1 U1781 ( .A(\DRAM_mem[17][2] ), .B(n2193), .S(n2224), .Z(n1607) );
  MUX2_X1 U1782 ( .A(\DRAM_mem[17][1] ), .B(n2194), .S(n2224), .Z(n1606) );
  MUX2_X1 U1783 ( .A(\DRAM_mem[17][0] ), .B(n2195), .S(n2224), .Z(n1605) );
  MUX2_X1 U1784 ( .A(\DRAM_mem[18][31] ), .B(n1139), .S(n2225), .Z(n1604) );
  MUX2_X1 U1785 ( .A(\DRAM_mem[18][30] ), .B(n1141), .S(n2225), .Z(n1603) );
  MUX2_X1 U1786 ( .A(\DRAM_mem[18][29] ), .B(n1142), .S(n2225), .Z(n1602) );
  MUX2_X1 U1787 ( .A(\DRAM_mem[18][28] ), .B(n1143), .S(n2225), .Z(n1601) );
  MUX2_X1 U1788 ( .A(\DRAM_mem[18][27] ), .B(n1144), .S(n2225), .Z(n1600) );
  MUX2_X1 U1789 ( .A(\DRAM_mem[18][26] ), .B(n1145), .S(n2225), .Z(n1599) );
  MUX2_X1 U1790 ( .A(\DRAM_mem[18][25] ), .B(n1146), .S(n2225), .Z(n1598) );
  MUX2_X1 U1791 ( .A(\DRAM_mem[18][24] ), .B(n1147), .S(n2225), .Z(n1597) );
  MUX2_X1 U1792 ( .A(\DRAM_mem[18][23] ), .B(n1148), .S(n2225), .Z(n1596) );
  MUX2_X1 U1793 ( .A(\DRAM_mem[18][22] ), .B(n1149), .S(n2225), .Z(n1595) );
  MUX2_X1 U1794 ( .A(\DRAM_mem[18][21] ), .B(n1150), .S(n2225), .Z(n1594) );
  MUX2_X1 U1795 ( .A(\DRAM_mem[18][20] ), .B(n1151), .S(n2225), .Z(n1593) );
  MUX2_X1 U1796 ( .A(\DRAM_mem[18][19] ), .B(n1152), .S(n2225), .Z(n1592) );
  MUX2_X1 U1797 ( .A(\DRAM_mem[18][18] ), .B(n1153), .S(n2225), .Z(n1591) );
  MUX2_X1 U1798 ( .A(\DRAM_mem[18][17] ), .B(n1154), .S(n2225), .Z(n1590) );
  MUX2_X1 U1799 ( .A(\DRAM_mem[18][16] ), .B(n1155), .S(n2225), .Z(n1589) );
  MUX2_X1 U1800 ( .A(\DRAM_mem[18][15] ), .B(n1156), .S(n2225), .Z(n1588) );
  MUX2_X1 U1801 ( .A(\DRAM_mem[18][14] ), .B(n2181), .S(n2225), .Z(n1587) );
  MUX2_X1 U1802 ( .A(\DRAM_mem[18][13] ), .B(n2182), .S(n2225), .Z(n1586) );
  MUX2_X1 U1803 ( .A(\DRAM_mem[18][12] ), .B(n2183), .S(n2225), .Z(n1585) );
  MUX2_X1 U1804 ( .A(\DRAM_mem[18][11] ), .B(n2184), .S(n2225), .Z(n1584) );
  MUX2_X1 U1805 ( .A(\DRAM_mem[18][10] ), .B(n2185), .S(n2225), .Z(n1583) );
  MUX2_X1 U1806 ( .A(\DRAM_mem[18][9] ), .B(n2186), .S(n2225), .Z(n1582) );
  MUX2_X1 U1807 ( .A(\DRAM_mem[18][8] ), .B(n2187), .S(n2225), .Z(n1581) );
  MUX2_X1 U1808 ( .A(\DRAM_mem[18][7] ), .B(n2188), .S(n2225), .Z(n1580) );
  MUX2_X1 U1809 ( .A(\DRAM_mem[18][6] ), .B(n2189), .S(n2225), .Z(n1579) );
  MUX2_X1 U1810 ( .A(\DRAM_mem[18][5] ), .B(n2190), .S(n2225), .Z(n1578) );
  MUX2_X1 U1811 ( .A(\DRAM_mem[18][4] ), .B(n2191), .S(n2225), .Z(n1577) );
  MUX2_X1 U1812 ( .A(\DRAM_mem[18][3] ), .B(n2192), .S(n2225), .Z(n1576) );
  MUX2_X1 U1813 ( .A(\DRAM_mem[18][2] ), .B(n2193), .S(n2225), .Z(n1575) );
  MUX2_X1 U1814 ( .A(\DRAM_mem[18][1] ), .B(n2194), .S(n2225), .Z(n1574) );
  MUX2_X1 U1815 ( .A(\DRAM_mem[18][0] ), .B(n2195), .S(n2225), .Z(n1573) );
  MUX2_X1 U1816 ( .A(\DRAM_mem[19][31] ), .B(n1139), .S(n2226), .Z(n1572) );
  MUX2_X1 U1817 ( .A(\DRAM_mem[19][30] ), .B(n1141), .S(n2226), .Z(n1571) );
  MUX2_X1 U1818 ( .A(\DRAM_mem[19][29] ), .B(n1142), .S(n2226), .Z(n1570) );
  MUX2_X1 U1819 ( .A(\DRAM_mem[19][28] ), .B(n1143), .S(n2226), .Z(n1569) );
  MUX2_X1 U1820 ( .A(\DRAM_mem[19][27] ), .B(n1144), .S(n2226), .Z(n1568) );
  MUX2_X1 U1821 ( .A(\DRAM_mem[19][26] ), .B(n1145), .S(n2226), .Z(n1567) );
  MUX2_X1 U1822 ( .A(\DRAM_mem[19][25] ), .B(n1146), .S(n2226), .Z(n1566) );
  MUX2_X1 U1823 ( .A(\DRAM_mem[19][24] ), .B(n1147), .S(n2226), .Z(n1565) );
  MUX2_X1 U1824 ( .A(\DRAM_mem[19][23] ), .B(n1148), .S(n2226), .Z(n1564) );
  MUX2_X1 U1825 ( .A(\DRAM_mem[19][22] ), .B(n1149), .S(n2226), .Z(n1563) );
  MUX2_X1 U1826 ( .A(\DRAM_mem[19][21] ), .B(n1150), .S(n2226), .Z(n1562) );
  MUX2_X1 U1827 ( .A(\DRAM_mem[19][20] ), .B(n1151), .S(n2226), .Z(n1561) );
  MUX2_X1 U1828 ( .A(\DRAM_mem[19][19] ), .B(n1152), .S(n2226), .Z(n1560) );
  MUX2_X1 U1829 ( .A(\DRAM_mem[19][18] ), .B(n1153), .S(n2226), .Z(n1559) );
  MUX2_X1 U1830 ( .A(\DRAM_mem[19][17] ), .B(n1154), .S(n2226), .Z(n1558) );
  MUX2_X1 U1831 ( .A(\DRAM_mem[19][16] ), .B(n1155), .S(n2226), .Z(n1557) );
  MUX2_X1 U1832 ( .A(\DRAM_mem[19][15] ), .B(n1156), .S(n2226), .Z(n1556) );
  MUX2_X1 U1833 ( .A(\DRAM_mem[19][14] ), .B(n2181), .S(n2226), .Z(n1555) );
  MUX2_X1 U1834 ( .A(\DRAM_mem[19][13] ), .B(n2182), .S(n2226), .Z(n1554) );
  MUX2_X1 U1835 ( .A(\DRAM_mem[19][12] ), .B(n2183), .S(n2226), .Z(n1553) );
  MUX2_X1 U1836 ( .A(\DRAM_mem[19][11] ), .B(n2184), .S(n2226), .Z(n1552) );
  MUX2_X1 U1837 ( .A(\DRAM_mem[19][10] ), .B(n2185), .S(n2226), .Z(n1551) );
  MUX2_X1 U1838 ( .A(\DRAM_mem[19][9] ), .B(n2186), .S(n2226), .Z(n1550) );
  MUX2_X1 U1839 ( .A(\DRAM_mem[19][8] ), .B(n2187), .S(n2226), .Z(n1549) );
  MUX2_X1 U1840 ( .A(\DRAM_mem[19][7] ), .B(n2188), .S(n2226), .Z(n1548) );
  MUX2_X1 U1841 ( .A(\DRAM_mem[19][6] ), .B(n2189), .S(n2226), .Z(n1547) );
  MUX2_X1 U1842 ( .A(\DRAM_mem[19][5] ), .B(n2190), .S(n2226), .Z(n1546) );
  MUX2_X1 U1843 ( .A(\DRAM_mem[19][4] ), .B(n2191), .S(n2226), .Z(n1545) );
  MUX2_X1 U1844 ( .A(\DRAM_mem[19][3] ), .B(n2192), .S(n2226), .Z(n1544) );
  MUX2_X1 U1845 ( .A(\DRAM_mem[19][2] ), .B(n2193), .S(n2226), .Z(n1543) );
  MUX2_X1 U1846 ( .A(\DRAM_mem[19][1] ), .B(n2194), .S(n2226), .Z(n1542) );
  MUX2_X1 U1847 ( .A(\DRAM_mem[19][0] ), .B(n2195), .S(n2226), .Z(n1541) );
  MUX2_X1 U1848 ( .A(\DRAM_mem[20][31] ), .B(n1139), .S(n2227), .Z(n1540) );
  MUX2_X1 U1849 ( .A(\DRAM_mem[20][30] ), .B(n1141), .S(n2227), .Z(n1539) );
  MUX2_X1 U1850 ( .A(\DRAM_mem[20][29] ), .B(n1142), .S(n2227), .Z(n1538) );
  MUX2_X1 U1851 ( .A(\DRAM_mem[20][28] ), .B(n1143), .S(n2227), .Z(n1537) );
  MUX2_X1 U1852 ( .A(\DRAM_mem[20][27] ), .B(n1144), .S(n2227), .Z(n1536) );
  MUX2_X1 U1853 ( .A(\DRAM_mem[20][26] ), .B(n1145), .S(n2227), .Z(n1535) );
  MUX2_X1 U1854 ( .A(\DRAM_mem[20][25] ), .B(n1146), .S(n2227), .Z(n1534) );
  MUX2_X1 U1855 ( .A(\DRAM_mem[20][24] ), .B(n1147), .S(n2227), .Z(n1533) );
  MUX2_X1 U1856 ( .A(\DRAM_mem[20][23] ), .B(n1148), .S(n2227), .Z(n1532) );
  MUX2_X1 U1857 ( .A(\DRAM_mem[20][22] ), .B(n1149), .S(n2227), .Z(n1531) );
  MUX2_X1 U1858 ( .A(\DRAM_mem[20][21] ), .B(n1150), .S(n2227), .Z(n1530) );
  MUX2_X1 U1859 ( .A(\DRAM_mem[20][20] ), .B(n1151), .S(n2227), .Z(n1529) );
  MUX2_X1 U1860 ( .A(\DRAM_mem[20][19] ), .B(n1152), .S(n2227), .Z(n1528) );
  MUX2_X1 U1861 ( .A(\DRAM_mem[20][18] ), .B(n1153), .S(n2227), .Z(n1527) );
  MUX2_X1 U1862 ( .A(\DRAM_mem[20][17] ), .B(n1154), .S(n2227), .Z(n1526) );
  MUX2_X1 U1863 ( .A(\DRAM_mem[20][16] ), .B(n1155), .S(n2227), .Z(n1525) );
  MUX2_X1 U1864 ( .A(\DRAM_mem[20][15] ), .B(n1156), .S(n2227), .Z(n1524) );
  MUX2_X1 U1865 ( .A(\DRAM_mem[20][14] ), .B(n2181), .S(n2227), .Z(n1523) );
  MUX2_X1 U1866 ( .A(\DRAM_mem[20][13] ), .B(n2182), .S(n2227), .Z(n1522) );
  MUX2_X1 U1867 ( .A(\DRAM_mem[20][12] ), .B(n2183), .S(n2227), .Z(n1521) );
  MUX2_X1 U1868 ( .A(\DRAM_mem[20][11] ), .B(n2184), .S(n2227), .Z(n1520) );
  MUX2_X1 U1869 ( .A(\DRAM_mem[20][10] ), .B(n2185), .S(n2227), .Z(n1519) );
  MUX2_X1 U1870 ( .A(\DRAM_mem[20][9] ), .B(n2186), .S(n2227), .Z(n1518) );
  MUX2_X1 U1871 ( .A(\DRAM_mem[20][8] ), .B(n2187), .S(n2227), .Z(n1517) );
  MUX2_X1 U1872 ( .A(\DRAM_mem[20][7] ), .B(n2188), .S(n2227), .Z(n1516) );
  MUX2_X1 U1873 ( .A(\DRAM_mem[20][6] ), .B(n2189), .S(n2227), .Z(n1515) );
  MUX2_X1 U1874 ( .A(\DRAM_mem[20][5] ), .B(n2190), .S(n2227), .Z(n1514) );
  MUX2_X1 U1875 ( .A(\DRAM_mem[20][4] ), .B(n2191), .S(n2227), .Z(n1513) );
  MUX2_X1 U1876 ( .A(\DRAM_mem[20][3] ), .B(n2192), .S(n2227), .Z(n1512) );
  MUX2_X1 U1877 ( .A(\DRAM_mem[20][2] ), .B(n2193), .S(n2227), .Z(n1511) );
  MUX2_X1 U1878 ( .A(\DRAM_mem[20][1] ), .B(n2194), .S(n2227), .Z(n1510) );
  MUX2_X1 U1879 ( .A(\DRAM_mem[20][0] ), .B(n2195), .S(n2227), .Z(n1509) );
  MUX2_X1 U1880 ( .A(\DRAM_mem[21][31] ), .B(n1139), .S(n2228), .Z(n1508) );
  MUX2_X1 U1881 ( .A(\DRAM_mem[21][30] ), .B(n1141), .S(n2228), .Z(n1507) );
  MUX2_X1 U1882 ( .A(\DRAM_mem[21][29] ), .B(n1142), .S(n2228), .Z(n1506) );
  MUX2_X1 U1883 ( .A(\DRAM_mem[21][28] ), .B(n1143), .S(n2228), .Z(n1505) );
  MUX2_X1 U1884 ( .A(\DRAM_mem[21][27] ), .B(n1144), .S(n2228), .Z(n1504) );
  MUX2_X1 U1885 ( .A(\DRAM_mem[21][26] ), .B(n1145), .S(n2228), .Z(n1503) );
  MUX2_X1 U1886 ( .A(\DRAM_mem[21][25] ), .B(n1146), .S(n2228), .Z(n1502) );
  MUX2_X1 U1887 ( .A(\DRAM_mem[21][24] ), .B(n1147), .S(n2228), .Z(n1501) );
  MUX2_X1 U1888 ( .A(\DRAM_mem[21][23] ), .B(n1148), .S(n2228), .Z(n1500) );
  MUX2_X1 U1889 ( .A(\DRAM_mem[21][22] ), .B(n1149), .S(n2228), .Z(n1499) );
  MUX2_X1 U1890 ( .A(\DRAM_mem[21][21] ), .B(n1150), .S(n2228), .Z(n1498) );
  MUX2_X1 U1891 ( .A(\DRAM_mem[21][20] ), .B(n1151), .S(n2228), .Z(n1497) );
  MUX2_X1 U1892 ( .A(\DRAM_mem[21][19] ), .B(n1152), .S(n2228), .Z(n1496) );
  MUX2_X1 U1893 ( .A(\DRAM_mem[21][18] ), .B(n1153), .S(n2228), .Z(n1495) );
  MUX2_X1 U1894 ( .A(\DRAM_mem[21][17] ), .B(n1154), .S(n2228), .Z(n1494) );
  MUX2_X1 U1895 ( .A(\DRAM_mem[21][16] ), .B(n1155), .S(n2228), .Z(n1493) );
  MUX2_X1 U1896 ( .A(\DRAM_mem[21][15] ), .B(n1156), .S(n2228), .Z(n1492) );
  MUX2_X1 U1897 ( .A(\DRAM_mem[21][14] ), .B(n2181), .S(n2228), .Z(n1491) );
  MUX2_X1 U1898 ( .A(\DRAM_mem[21][13] ), .B(n2182), .S(n2228), .Z(n1490) );
  MUX2_X1 U1899 ( .A(\DRAM_mem[21][12] ), .B(n2183), .S(n2228), .Z(n1489) );
  MUX2_X1 U1900 ( .A(\DRAM_mem[21][11] ), .B(n2184), .S(n2228), .Z(n1488) );
  MUX2_X1 U1901 ( .A(\DRAM_mem[21][10] ), .B(n2185), .S(n2228), .Z(n1487) );
  MUX2_X1 U1902 ( .A(\DRAM_mem[21][9] ), .B(n2186), .S(n2228), .Z(n1486) );
  MUX2_X1 U1903 ( .A(\DRAM_mem[21][8] ), .B(n2187), .S(n2228), .Z(n1485) );
  MUX2_X1 U1904 ( .A(\DRAM_mem[21][7] ), .B(n2188), .S(n2228), .Z(n1484) );
  MUX2_X1 U1905 ( .A(\DRAM_mem[21][6] ), .B(n2189), .S(n2228), .Z(n1483) );
  MUX2_X1 U1906 ( .A(\DRAM_mem[21][5] ), .B(n2190), .S(n2228), .Z(n1482) );
  MUX2_X1 U1907 ( .A(\DRAM_mem[21][4] ), .B(n2191), .S(n2228), .Z(n1481) );
  MUX2_X1 U1908 ( .A(\DRAM_mem[21][3] ), .B(n2192), .S(n2228), .Z(n1480) );
  MUX2_X1 U1909 ( .A(\DRAM_mem[21][2] ), .B(n2193), .S(n2228), .Z(n1479) );
  MUX2_X1 U1910 ( .A(\DRAM_mem[21][1] ), .B(n2194), .S(n2228), .Z(n1478) );
  MUX2_X1 U1911 ( .A(\DRAM_mem[21][0] ), .B(n2195), .S(n2228), .Z(n1477) );
  MUX2_X1 U1912 ( .A(\DRAM_mem[22][31] ), .B(n1139), .S(n2229), .Z(n1476) );
  MUX2_X1 U1913 ( .A(\DRAM_mem[22][30] ), .B(n1141), .S(n2229), .Z(n1475) );
  MUX2_X1 U1914 ( .A(\DRAM_mem[22][29] ), .B(n1142), .S(n2229), .Z(n1474) );
  MUX2_X1 U1915 ( .A(\DRAM_mem[22][28] ), .B(n1143), .S(n2229), .Z(n1473) );
  MUX2_X1 U1916 ( .A(\DRAM_mem[22][27] ), .B(n1144), .S(n2229), .Z(n1472) );
  MUX2_X1 U1917 ( .A(\DRAM_mem[22][26] ), .B(n1145), .S(n2229), .Z(n1471) );
  MUX2_X1 U1918 ( .A(\DRAM_mem[22][25] ), .B(n1146), .S(n2229), .Z(n1470) );
  MUX2_X1 U1919 ( .A(\DRAM_mem[22][24] ), .B(n1147), .S(n2229), .Z(n1469) );
  MUX2_X1 U1920 ( .A(\DRAM_mem[22][23] ), .B(n1148), .S(n2229), .Z(n1468) );
  MUX2_X1 U1921 ( .A(\DRAM_mem[22][22] ), .B(n1149), .S(n2229), .Z(n1467) );
  MUX2_X1 U1922 ( .A(\DRAM_mem[22][21] ), .B(n1150), .S(n2229), .Z(n1466) );
  MUX2_X1 U1923 ( .A(\DRAM_mem[22][20] ), .B(n1151), .S(n2229), .Z(n1465) );
  MUX2_X1 U1924 ( .A(\DRAM_mem[22][19] ), .B(n1152), .S(n2229), .Z(n1464) );
  MUX2_X1 U1925 ( .A(\DRAM_mem[22][18] ), .B(n1153), .S(n2229), .Z(n1463) );
  MUX2_X1 U1926 ( .A(\DRAM_mem[22][17] ), .B(n1154), .S(n2229), .Z(n1462) );
  MUX2_X1 U1927 ( .A(\DRAM_mem[22][16] ), .B(n1155), .S(n2229), .Z(n1461) );
  MUX2_X1 U1928 ( .A(\DRAM_mem[22][15] ), .B(n1156), .S(n2229), .Z(n1460) );
  MUX2_X1 U1929 ( .A(\DRAM_mem[22][14] ), .B(n2181), .S(n2229), .Z(n1459) );
  MUX2_X1 U1930 ( .A(\DRAM_mem[22][13] ), .B(n2182), .S(n2229), .Z(n1458) );
  MUX2_X1 U1931 ( .A(\DRAM_mem[22][12] ), .B(n2183), .S(n2229), .Z(n1457) );
  MUX2_X1 U1932 ( .A(\DRAM_mem[22][11] ), .B(n2184), .S(n2229), .Z(n1456) );
  MUX2_X1 U1933 ( .A(\DRAM_mem[22][10] ), .B(n2185), .S(n2229), .Z(n1455) );
  MUX2_X1 U1934 ( .A(\DRAM_mem[22][9] ), .B(n2186), .S(n2229), .Z(n1454) );
  MUX2_X1 U1935 ( .A(\DRAM_mem[22][8] ), .B(n2187), .S(n2229), .Z(n1453) );
  MUX2_X1 U1936 ( .A(\DRAM_mem[22][7] ), .B(n2188), .S(n2229), .Z(n1452) );
  MUX2_X1 U1937 ( .A(\DRAM_mem[22][6] ), .B(n2189), .S(n2229), .Z(n1451) );
  MUX2_X1 U1938 ( .A(\DRAM_mem[22][5] ), .B(n2190), .S(n2229), .Z(n1450) );
  MUX2_X1 U1939 ( .A(\DRAM_mem[22][4] ), .B(n2191), .S(n2229), .Z(n1449) );
  MUX2_X1 U1940 ( .A(\DRAM_mem[22][3] ), .B(n2192), .S(n2229), .Z(n1448) );
  MUX2_X1 U1941 ( .A(\DRAM_mem[22][2] ), .B(n2193), .S(n2229), .Z(n1447) );
  MUX2_X1 U1942 ( .A(\DRAM_mem[22][1] ), .B(n2194), .S(n2229), .Z(n1446) );
  MUX2_X1 U1943 ( .A(\DRAM_mem[22][0] ), .B(n2195), .S(n2229), .Z(n1445) );
  MUX2_X1 U1944 ( .A(\DRAM_mem[23][31] ), .B(n1139), .S(n2230), .Z(n1444) );
  MUX2_X1 U1945 ( .A(\DRAM_mem[23][30] ), .B(n1141), .S(n2230), .Z(n1443) );
  MUX2_X1 U1946 ( .A(\DRAM_mem[23][29] ), .B(n1142), .S(n2230), .Z(n1442) );
  MUX2_X1 U1947 ( .A(\DRAM_mem[23][28] ), .B(n1143), .S(n2230), .Z(n1441) );
  MUX2_X1 U1948 ( .A(\DRAM_mem[23][27] ), .B(n1144), .S(n2230), .Z(n1440) );
  MUX2_X1 U1949 ( .A(\DRAM_mem[23][26] ), .B(n1145), .S(n2230), .Z(n1439) );
  MUX2_X1 U1950 ( .A(\DRAM_mem[23][25] ), .B(n1146), .S(n2230), .Z(n1438) );
  MUX2_X1 U1951 ( .A(\DRAM_mem[23][24] ), .B(n1147), .S(n2230), .Z(n1437) );
  MUX2_X1 U1952 ( .A(\DRAM_mem[23][23] ), .B(n1148), .S(n2230), .Z(n1436) );
  MUX2_X1 U1953 ( .A(\DRAM_mem[23][22] ), .B(n1149), .S(n2230), .Z(n1435) );
  MUX2_X1 U1954 ( .A(\DRAM_mem[23][21] ), .B(n1150), .S(n2230), .Z(n1434) );
  MUX2_X1 U1955 ( .A(\DRAM_mem[23][20] ), .B(n1151), .S(n2230), .Z(n1433) );
  MUX2_X1 U1956 ( .A(\DRAM_mem[23][19] ), .B(n1152), .S(n2230), .Z(n1432) );
  MUX2_X1 U1957 ( .A(\DRAM_mem[23][18] ), .B(n1153), .S(n2230), .Z(n1431) );
  MUX2_X1 U1958 ( .A(\DRAM_mem[23][17] ), .B(n1154), .S(n2230), .Z(n1430) );
  MUX2_X1 U1959 ( .A(\DRAM_mem[23][16] ), .B(n1155), .S(n2230), .Z(n1429) );
  MUX2_X1 U1960 ( .A(\DRAM_mem[23][15] ), .B(n1156), .S(n2230), .Z(n1428) );
  MUX2_X1 U1961 ( .A(\DRAM_mem[23][14] ), .B(n2181), .S(n2230), .Z(n1427) );
  MUX2_X1 U1962 ( .A(\DRAM_mem[23][13] ), .B(n2182), .S(n2230), .Z(n1426) );
  MUX2_X1 U1963 ( .A(\DRAM_mem[23][12] ), .B(n2183), .S(n2230), .Z(n1425) );
  MUX2_X1 U1964 ( .A(\DRAM_mem[23][11] ), .B(n2184), .S(n2230), .Z(n1424) );
  MUX2_X1 U1965 ( .A(\DRAM_mem[23][10] ), .B(n2185), .S(n2230), .Z(n1423) );
  MUX2_X1 U1966 ( .A(\DRAM_mem[23][9] ), .B(n2186), .S(n2230), .Z(n1422) );
  MUX2_X1 U1967 ( .A(\DRAM_mem[23][8] ), .B(n2187), .S(n2230), .Z(n1421) );
  MUX2_X1 U1968 ( .A(\DRAM_mem[23][7] ), .B(n2188), .S(n2230), .Z(n1420) );
  MUX2_X1 U1969 ( .A(\DRAM_mem[23][6] ), .B(n2189), .S(n2230), .Z(n1419) );
  MUX2_X1 U1970 ( .A(\DRAM_mem[23][5] ), .B(n2190), .S(n2230), .Z(n1418) );
  MUX2_X1 U1971 ( .A(\DRAM_mem[23][4] ), .B(n2191), .S(n2230), .Z(n1417) );
  MUX2_X1 U1972 ( .A(\DRAM_mem[23][3] ), .B(n2192), .S(n2230), .Z(n1416) );
  MUX2_X1 U1973 ( .A(\DRAM_mem[23][2] ), .B(n2193), .S(n2230), .Z(n1415) );
  MUX2_X1 U1974 ( .A(\DRAM_mem[23][1] ), .B(n2194), .S(n2230), .Z(n1414) );
  MUX2_X1 U1975 ( .A(\DRAM_mem[23][0] ), .B(n2195), .S(n2230), .Z(n1413) );
  AND3_X1 U1976 ( .A1(n2212), .A2(n132), .A3(n164), .ZN(n2223) );
  MUX2_X1 U1977 ( .A(\DRAM_mem[24][31] ), .B(n1139), .S(n2231), .Z(n1412) );
  MUX2_X1 U1978 ( .A(\DRAM_mem[24][30] ), .B(n1141), .S(n2231), .Z(n1411) );
  MUX2_X1 U1979 ( .A(\DRAM_mem[24][29] ), .B(n1142), .S(n2231), .Z(n1410) );
  MUX2_X1 U1980 ( .A(\DRAM_mem[24][28] ), .B(n1143), .S(n2231), .Z(n1409) );
  MUX2_X1 U1981 ( .A(\DRAM_mem[24][27] ), .B(n1144), .S(n2231), .Z(n1408) );
  MUX2_X1 U1982 ( .A(\DRAM_mem[24][26] ), .B(n1145), .S(n2231), .Z(n1407) );
  MUX2_X1 U1983 ( .A(\DRAM_mem[24][25] ), .B(n1146), .S(n2231), .Z(n1406) );
  MUX2_X1 U1984 ( .A(\DRAM_mem[24][24] ), .B(n1147), .S(n2231), .Z(n1405) );
  MUX2_X1 U1985 ( .A(\DRAM_mem[24][23] ), .B(n1148), .S(n2231), .Z(n1404) );
  MUX2_X1 U1986 ( .A(\DRAM_mem[24][22] ), .B(n1149), .S(n2231), .Z(n1403) );
  MUX2_X1 U1987 ( .A(\DRAM_mem[24][21] ), .B(n1150), .S(n2231), .Z(n1402) );
  MUX2_X1 U1988 ( .A(\DRAM_mem[24][20] ), .B(n1151), .S(n2231), .Z(n1401) );
  MUX2_X1 U1989 ( .A(\DRAM_mem[24][19] ), .B(n1152), .S(n2231), .Z(n1400) );
  MUX2_X1 U1990 ( .A(\DRAM_mem[24][18] ), .B(n1153), .S(n2231), .Z(n1399) );
  MUX2_X1 U1991 ( .A(\DRAM_mem[24][17] ), .B(n1154), .S(n2231), .Z(n1398) );
  MUX2_X1 U1992 ( .A(\DRAM_mem[24][16] ), .B(n1155), .S(n2231), .Z(n1397) );
  MUX2_X1 U1993 ( .A(\DRAM_mem[24][15] ), .B(n1156), .S(n2231), .Z(n1396) );
  MUX2_X1 U1994 ( .A(\DRAM_mem[24][14] ), .B(n2181), .S(n2231), .Z(n1395) );
  MUX2_X1 U1995 ( .A(\DRAM_mem[24][13] ), .B(n2182), .S(n2231), .Z(n1394) );
  MUX2_X1 U1996 ( .A(\DRAM_mem[24][12] ), .B(n2183), .S(n2231), .Z(n1393) );
  MUX2_X1 U1997 ( .A(\DRAM_mem[24][11] ), .B(n2184), .S(n2231), .Z(n1392) );
  MUX2_X1 U1998 ( .A(\DRAM_mem[24][10] ), .B(n2185), .S(n2231), .Z(n1391) );
  MUX2_X1 U1999 ( .A(\DRAM_mem[24][9] ), .B(n2186), .S(n2231), .Z(n1390) );
  MUX2_X1 U2000 ( .A(\DRAM_mem[24][8] ), .B(n2187), .S(n2231), .Z(n1389) );
  MUX2_X1 U2001 ( .A(\DRAM_mem[24][7] ), .B(n2188), .S(n2231), .Z(n1388) );
  MUX2_X1 U2002 ( .A(\DRAM_mem[24][6] ), .B(n2189), .S(n2231), .Z(n1387) );
  MUX2_X1 U2003 ( .A(\DRAM_mem[24][5] ), .B(n2190), .S(n2231), .Z(n1386) );
  MUX2_X1 U2004 ( .A(\DRAM_mem[24][4] ), .B(n2191), .S(n2231), .Z(n1385) );
  MUX2_X1 U2005 ( .A(\DRAM_mem[24][3] ), .B(n2192), .S(n2231), .Z(n1384) );
  MUX2_X1 U2006 ( .A(\DRAM_mem[24][2] ), .B(n2193), .S(n2231), .Z(n1383) );
  MUX2_X1 U2007 ( .A(\DRAM_mem[24][1] ), .B(n2194), .S(n2231), .Z(n1382) );
  MUX2_X1 U2008 ( .A(\DRAM_mem[24][0] ), .B(n2195), .S(n2231), .Z(n1381) );
  NOR3_X1 U2009 ( .A1(Addr[1]), .A2(n112), .A3(Addr[0]), .ZN(n2196) );
  MUX2_X1 U2010 ( .A(\DRAM_mem[25][31] ), .B(n1139), .S(n2233), .Z(n1380) );
  MUX2_X1 U2011 ( .A(\DRAM_mem[25][30] ), .B(n1141), .S(n2233), .Z(n1379) );
  MUX2_X1 U2012 ( .A(\DRAM_mem[25][29] ), .B(n1142), .S(n2233), .Z(n1378) );
  MUX2_X1 U2013 ( .A(\DRAM_mem[25][28] ), .B(n1143), .S(n2233), .Z(n1377) );
  MUX2_X1 U2014 ( .A(\DRAM_mem[25][27] ), .B(n1144), .S(n2233), .Z(n1376) );
  MUX2_X1 U2015 ( .A(\DRAM_mem[25][26] ), .B(n1145), .S(n2233), .Z(n1375) );
  MUX2_X1 U2016 ( .A(\DRAM_mem[25][25] ), .B(n1146), .S(n2233), .Z(n1374) );
  MUX2_X1 U2017 ( .A(\DRAM_mem[25][24] ), .B(n1147), .S(n2233), .Z(n1373) );
  MUX2_X1 U2018 ( .A(\DRAM_mem[25][23] ), .B(n1148), .S(n2233), .Z(n1372) );
  MUX2_X1 U2019 ( .A(\DRAM_mem[25][22] ), .B(n1149), .S(n2233), .Z(n1371) );
  MUX2_X1 U2020 ( .A(\DRAM_mem[25][21] ), .B(n1150), .S(n2233), .Z(n1370) );
  MUX2_X1 U2021 ( .A(\DRAM_mem[25][20] ), .B(n1151), .S(n2233), .Z(n1369) );
  MUX2_X1 U2022 ( .A(\DRAM_mem[25][19] ), .B(n1152), .S(n2233), .Z(n1368) );
  MUX2_X1 U2023 ( .A(\DRAM_mem[25][18] ), .B(n1153), .S(n2233), .Z(n1367) );
  MUX2_X1 U2024 ( .A(\DRAM_mem[25][17] ), .B(n1154), .S(n2233), .Z(n1366) );
  MUX2_X1 U2025 ( .A(\DRAM_mem[25][16] ), .B(n1155), .S(n2233), .Z(n1365) );
  MUX2_X1 U2026 ( .A(\DRAM_mem[25][15] ), .B(n1156), .S(n2233), .Z(n1364) );
  MUX2_X1 U2027 ( .A(\DRAM_mem[25][14] ), .B(n2181), .S(n2233), .Z(n1363) );
  MUX2_X1 U2028 ( .A(\DRAM_mem[25][13] ), .B(n2182), .S(n2233), .Z(n1362) );
  MUX2_X1 U2029 ( .A(\DRAM_mem[25][12] ), .B(n2183), .S(n2233), .Z(n1361) );
  MUX2_X1 U2030 ( .A(\DRAM_mem[25][11] ), .B(n2184), .S(n2233), .Z(n1360) );
  MUX2_X1 U2031 ( .A(\DRAM_mem[25][10] ), .B(n2185), .S(n2233), .Z(n1359) );
  MUX2_X1 U2032 ( .A(\DRAM_mem[25][9] ), .B(n2186), .S(n2233), .Z(n1358) );
  MUX2_X1 U2033 ( .A(\DRAM_mem[25][8] ), .B(n2187), .S(n2233), .Z(n1357) );
  MUX2_X1 U2034 ( .A(\DRAM_mem[25][7] ), .B(n2188), .S(n2233), .Z(n1356) );
  MUX2_X1 U2035 ( .A(\DRAM_mem[25][6] ), .B(n2189), .S(n2233), .Z(n1355) );
  MUX2_X1 U2036 ( .A(\DRAM_mem[25][5] ), .B(n2190), .S(n2233), .Z(n1354) );
  MUX2_X1 U2037 ( .A(\DRAM_mem[25][4] ), .B(n2191), .S(n2233), .Z(n1353) );
  MUX2_X1 U2038 ( .A(\DRAM_mem[25][3] ), .B(n2192), .S(n2233), .Z(n1352) );
  MUX2_X1 U2039 ( .A(\DRAM_mem[25][2] ), .B(n2193), .S(n2233), .Z(n1351) );
  MUX2_X1 U2040 ( .A(\DRAM_mem[25][1] ), .B(n2194), .S(n2233), .Z(n1350) );
  MUX2_X1 U2041 ( .A(\DRAM_mem[25][0] ), .B(n2195), .S(n2233), .Z(n1349) );
  NOR3_X1 U2042 ( .A1(Addr[1]), .A2(n112), .A3(n2234), .ZN(n2199) );
  MUX2_X1 U2043 ( .A(\DRAM_mem[26][31] ), .B(n1139), .S(n2235), .Z(n1348) );
  MUX2_X1 U2044 ( .A(\DRAM_mem[26][30] ), .B(n1141), .S(n2235), .Z(n1347) );
  MUX2_X1 U2045 ( .A(\DRAM_mem[26][29] ), .B(n1142), .S(n2235), .Z(n1346) );
  MUX2_X1 U2046 ( .A(\DRAM_mem[26][28] ), .B(n1143), .S(n2235), .Z(n1345) );
  MUX2_X1 U2047 ( .A(\DRAM_mem[26][27] ), .B(n1144), .S(n2235), .Z(n1344) );
  MUX2_X1 U2048 ( .A(\DRAM_mem[26][26] ), .B(n1145), .S(n2235), .Z(n1343) );
  MUX2_X1 U2049 ( .A(\DRAM_mem[26][25] ), .B(n1146), .S(n2235), .Z(n1342) );
  MUX2_X1 U2050 ( .A(\DRAM_mem[26][24] ), .B(n1147), .S(n2235), .Z(n1341) );
  MUX2_X1 U2051 ( .A(\DRAM_mem[26][23] ), .B(n1148), .S(n2235), .Z(n1340) );
  MUX2_X1 U2052 ( .A(\DRAM_mem[26][22] ), .B(n1149), .S(n2235), .Z(n1339) );
  MUX2_X1 U2053 ( .A(\DRAM_mem[26][21] ), .B(n1150), .S(n2235), .Z(n1338) );
  MUX2_X1 U2054 ( .A(\DRAM_mem[26][20] ), .B(n1151), .S(n2235), .Z(n1337) );
  MUX2_X1 U2055 ( .A(\DRAM_mem[26][19] ), .B(n1152), .S(n2235), .Z(n1336) );
  MUX2_X1 U2056 ( .A(\DRAM_mem[26][18] ), .B(n1153), .S(n2235), .Z(n1335) );
  MUX2_X1 U2057 ( .A(\DRAM_mem[26][17] ), .B(n1154), .S(n2235), .Z(n1334) );
  MUX2_X1 U2058 ( .A(\DRAM_mem[26][16] ), .B(n1155), .S(n2235), .Z(n1333) );
  MUX2_X1 U2059 ( .A(\DRAM_mem[26][15] ), .B(n1156), .S(n2235), .Z(n1332) );
  MUX2_X1 U2060 ( .A(\DRAM_mem[26][14] ), .B(n2181), .S(n2235), .Z(n1331) );
  MUX2_X1 U2061 ( .A(\DRAM_mem[26][13] ), .B(n2182), .S(n2235), .Z(n1330) );
  MUX2_X1 U2062 ( .A(\DRAM_mem[26][12] ), .B(n2183), .S(n2235), .Z(n1329) );
  MUX2_X1 U2063 ( .A(\DRAM_mem[26][11] ), .B(n2184), .S(n2235), .Z(n1328) );
  MUX2_X1 U2064 ( .A(\DRAM_mem[26][10] ), .B(n2185), .S(n2235), .Z(n1327) );
  MUX2_X1 U2065 ( .A(\DRAM_mem[26][9] ), .B(n2186), .S(n2235), .Z(n1326) );
  MUX2_X1 U2066 ( .A(\DRAM_mem[26][8] ), .B(n2187), .S(n2235), .Z(n1325) );
  MUX2_X1 U2067 ( .A(\DRAM_mem[26][7] ), .B(n2188), .S(n2235), .Z(n1324) );
  MUX2_X1 U2068 ( .A(\DRAM_mem[26][6] ), .B(n2189), .S(n2235), .Z(n1323) );
  MUX2_X1 U2069 ( .A(\DRAM_mem[26][5] ), .B(n2190), .S(n2235), .Z(n1322) );
  MUX2_X1 U2070 ( .A(\DRAM_mem[26][4] ), .B(n2191), .S(n2235), .Z(n1321) );
  MUX2_X1 U2071 ( .A(\DRAM_mem[26][3] ), .B(n2192), .S(n2235), .Z(n1320) );
  MUX2_X1 U2072 ( .A(\DRAM_mem[26][2] ), .B(n2193), .S(n2235), .Z(n1319) );
  MUX2_X1 U2073 ( .A(\DRAM_mem[26][1] ), .B(n2194), .S(n2235), .Z(n1318) );
  MUX2_X1 U2074 ( .A(\DRAM_mem[26][0] ), .B(n2195), .S(n2235), .Z(n1317) );
  NOR3_X1 U2075 ( .A1(Addr[0]), .A2(n112), .A3(n2236), .ZN(n2201) );
  MUX2_X1 U2076 ( .A(\DRAM_mem[27][31] ), .B(n1139), .S(n2237), .Z(n1316) );
  MUX2_X1 U2077 ( .A(\DRAM_mem[27][30] ), .B(n1141), .S(n2237), .Z(n1315) );
  MUX2_X1 U2078 ( .A(\DRAM_mem[27][29] ), .B(n1142), .S(n2237), .Z(n1314) );
  MUX2_X1 U2079 ( .A(\DRAM_mem[27][28] ), .B(n1143), .S(n2237), .Z(n1313) );
  MUX2_X1 U2080 ( .A(\DRAM_mem[27][27] ), .B(n1144), .S(n2237), .Z(n1312) );
  MUX2_X1 U2081 ( .A(\DRAM_mem[27][26] ), .B(n1145), .S(n2237), .Z(n1311) );
  MUX2_X1 U2082 ( .A(\DRAM_mem[27][25] ), .B(n1146), .S(n2237), .Z(n1310) );
  MUX2_X1 U2083 ( .A(\DRAM_mem[27][24] ), .B(n1147), .S(n2237), .Z(n1309) );
  MUX2_X1 U2084 ( .A(\DRAM_mem[27][23] ), .B(n1148), .S(n2237), .Z(n1308) );
  MUX2_X1 U2085 ( .A(\DRAM_mem[27][22] ), .B(n1149), .S(n2237), .Z(n1307) );
  MUX2_X1 U2086 ( .A(\DRAM_mem[27][21] ), .B(n1150), .S(n2237), .Z(n1306) );
  MUX2_X1 U2087 ( .A(\DRAM_mem[27][20] ), .B(n1151), .S(n2237), .Z(n1305) );
  MUX2_X1 U2088 ( .A(\DRAM_mem[27][19] ), .B(n1152), .S(n2237), .Z(n1304) );
  MUX2_X1 U2089 ( .A(\DRAM_mem[27][18] ), .B(n1153), .S(n2237), .Z(n1303) );
  MUX2_X1 U2090 ( .A(\DRAM_mem[27][17] ), .B(n1154), .S(n2237), .Z(n1302) );
  MUX2_X1 U2091 ( .A(\DRAM_mem[27][16] ), .B(n1155), .S(n2237), .Z(n1301) );
  MUX2_X1 U2092 ( .A(\DRAM_mem[27][15] ), .B(n1156), .S(n2237), .Z(n1300) );
  MUX2_X1 U2093 ( .A(\DRAM_mem[27][14] ), .B(n2181), .S(n2237), .Z(n1299) );
  MUX2_X1 U2094 ( .A(\DRAM_mem[27][13] ), .B(n2182), .S(n2237), .Z(n1298) );
  MUX2_X1 U2095 ( .A(\DRAM_mem[27][12] ), .B(n2183), .S(n2237), .Z(n1297) );
  MUX2_X1 U2096 ( .A(\DRAM_mem[27][11] ), .B(n2184), .S(n2237), .Z(n1296) );
  MUX2_X1 U2097 ( .A(\DRAM_mem[27][10] ), .B(n2185), .S(n2237), .Z(n1295) );
  MUX2_X1 U2098 ( .A(\DRAM_mem[27][9] ), .B(n2186), .S(n2237), .Z(n1294) );
  MUX2_X1 U2099 ( .A(\DRAM_mem[27][8] ), .B(n2187), .S(n2237), .Z(n1293) );
  MUX2_X1 U2100 ( .A(\DRAM_mem[27][7] ), .B(n2188), .S(n2237), .Z(n1292) );
  MUX2_X1 U2101 ( .A(\DRAM_mem[27][6] ), .B(n2189), .S(n2237), .Z(n1291) );
  MUX2_X1 U2102 ( .A(\DRAM_mem[27][5] ), .B(n2190), .S(n2237), .Z(n1290) );
  MUX2_X1 U2103 ( .A(\DRAM_mem[27][4] ), .B(n2191), .S(n2237), .Z(n1289) );
  MUX2_X1 U2104 ( .A(\DRAM_mem[27][3] ), .B(n2192), .S(n2237), .Z(n1288) );
  MUX2_X1 U2105 ( .A(\DRAM_mem[27][2] ), .B(n2193), .S(n2237), .Z(n1287) );
  MUX2_X1 U2106 ( .A(\DRAM_mem[27][1] ), .B(n2194), .S(n2237), .Z(n1286) );
  MUX2_X1 U2107 ( .A(\DRAM_mem[27][0] ), .B(n2195), .S(n2237), .Z(n1285) );
  NOR3_X1 U2108 ( .A1(n2234), .A2(n112), .A3(n2236), .ZN(n2203) );
  MUX2_X1 U2109 ( .A(\DRAM_mem[28][31] ), .B(n1139), .S(n2238), .Z(n1284) );
  MUX2_X1 U2110 ( .A(\DRAM_mem[28][30] ), .B(n1141), .S(n2238), .Z(n1283) );
  MUX2_X1 U2111 ( .A(\DRAM_mem[28][29] ), .B(n1142), .S(n2238), .Z(n1282) );
  MUX2_X1 U2112 ( .A(\DRAM_mem[28][28] ), .B(n1143), .S(n2238), .Z(n1281) );
  MUX2_X1 U2113 ( .A(\DRAM_mem[28][27] ), .B(n1144), .S(n2238), .Z(n1280) );
  MUX2_X1 U2114 ( .A(\DRAM_mem[28][26] ), .B(n1145), .S(n2238), .Z(n1279) );
  MUX2_X1 U2115 ( .A(\DRAM_mem[28][25] ), .B(n1146), .S(n2238), .Z(n1278) );
  MUX2_X1 U2116 ( .A(\DRAM_mem[28][24] ), .B(n1147), .S(n2238), .Z(n1277) );
  MUX2_X1 U2117 ( .A(\DRAM_mem[28][23] ), .B(n1148), .S(n2238), .Z(n1276) );
  MUX2_X1 U2118 ( .A(\DRAM_mem[28][22] ), .B(n1149), .S(n2238), .Z(n1275) );
  MUX2_X1 U2119 ( .A(\DRAM_mem[28][21] ), .B(n1150), .S(n2238), .Z(n1274) );
  MUX2_X1 U2120 ( .A(\DRAM_mem[28][20] ), .B(n1151), .S(n2238), .Z(n1273) );
  MUX2_X1 U2121 ( .A(\DRAM_mem[28][19] ), .B(n1152), .S(n2238), .Z(n1272) );
  MUX2_X1 U2122 ( .A(\DRAM_mem[28][18] ), .B(n1153), .S(n2238), .Z(n1271) );
  MUX2_X1 U2123 ( .A(\DRAM_mem[28][17] ), .B(n1154), .S(n2238), .Z(n1270) );
  MUX2_X1 U2124 ( .A(\DRAM_mem[28][16] ), .B(n1155), .S(n2238), .Z(n1269) );
  MUX2_X1 U2125 ( .A(\DRAM_mem[28][15] ), .B(n1156), .S(n2238), .Z(n1268) );
  MUX2_X1 U2126 ( .A(\DRAM_mem[28][14] ), .B(n2181), .S(n2238), .Z(n1267) );
  MUX2_X1 U2127 ( .A(\DRAM_mem[28][13] ), .B(n2182), .S(n2238), .Z(n1266) );
  MUX2_X1 U2128 ( .A(\DRAM_mem[28][12] ), .B(n2183), .S(n2238), .Z(n1265) );
  MUX2_X1 U2129 ( .A(\DRAM_mem[28][11] ), .B(n2184), .S(n2238), .Z(n1264) );
  MUX2_X1 U2130 ( .A(\DRAM_mem[28][10] ), .B(n2185), .S(n2238), .Z(n1263) );
  MUX2_X1 U2131 ( .A(\DRAM_mem[28][9] ), .B(n2186), .S(n2238), .Z(n1262) );
  MUX2_X1 U2132 ( .A(\DRAM_mem[28][8] ), .B(n2187), .S(n2238), .Z(n1261) );
  MUX2_X1 U2133 ( .A(\DRAM_mem[28][7] ), .B(n2188), .S(n2238), .Z(n1260) );
  MUX2_X1 U2134 ( .A(\DRAM_mem[28][6] ), .B(n2189), .S(n2238), .Z(n1259) );
  MUX2_X1 U2135 ( .A(\DRAM_mem[28][5] ), .B(n2190), .S(n2238), .Z(n1258) );
  MUX2_X1 U2136 ( .A(\DRAM_mem[28][4] ), .B(n2191), .S(n2238), .Z(n1257) );
  MUX2_X1 U2137 ( .A(\DRAM_mem[28][3] ), .B(n2192), .S(n2238), .Z(n1256) );
  MUX2_X1 U2138 ( .A(\DRAM_mem[28][2] ), .B(n2193), .S(n2238), .Z(n1255) );
  MUX2_X1 U2139 ( .A(\DRAM_mem[28][1] ), .B(n2194), .S(n2238), .Z(n1254) );
  MUX2_X1 U2140 ( .A(\DRAM_mem[28][0] ), .B(n2195), .S(n2238), .Z(n1253) );
  AND3_X1 U2141 ( .A1(n2234), .A2(n2236), .A3(n113), .ZN(n2205) );
  MUX2_X1 U2142 ( .A(\DRAM_mem[29][31] ), .B(n1139), .S(n2239), .Z(n1252) );
  MUX2_X1 U2143 ( .A(\DRAM_mem[29][30] ), .B(n1141), .S(n2239), .Z(n1251) );
  MUX2_X1 U2144 ( .A(\DRAM_mem[29][29] ), .B(n1142), .S(n2239), .Z(n1250) );
  MUX2_X1 U2145 ( .A(\DRAM_mem[29][28] ), .B(n1143), .S(n2239), .Z(n1249) );
  MUX2_X1 U2146 ( .A(\DRAM_mem[29][27] ), .B(n1144), .S(n2239), .Z(n1248) );
  MUX2_X1 U2147 ( .A(\DRAM_mem[29][26] ), .B(n1145), .S(n2239), .Z(n1247) );
  MUX2_X1 U2148 ( .A(\DRAM_mem[29][25] ), .B(n1146), .S(n2239), .Z(n1246) );
  MUX2_X1 U2149 ( .A(\DRAM_mem[29][24] ), .B(n1147), .S(n2239), .Z(n1245) );
  MUX2_X1 U2150 ( .A(\DRAM_mem[29][23] ), .B(n1148), .S(n2239), .Z(n1244) );
  MUX2_X1 U2151 ( .A(\DRAM_mem[29][22] ), .B(n1149), .S(n2239), .Z(n1243) );
  MUX2_X1 U2152 ( .A(\DRAM_mem[29][21] ), .B(n1150), .S(n2239), .Z(n1242) );
  MUX2_X1 U2153 ( .A(\DRAM_mem[29][20] ), .B(n1151), .S(n2239), .Z(n1241) );
  MUX2_X1 U2154 ( .A(\DRAM_mem[29][19] ), .B(n1152), .S(n2239), .Z(n1240) );
  MUX2_X1 U2155 ( .A(\DRAM_mem[29][18] ), .B(n1153), .S(n2239), .Z(n1239) );
  MUX2_X1 U2156 ( .A(\DRAM_mem[29][17] ), .B(n1154), .S(n2239), .Z(n1238) );
  MUX2_X1 U2157 ( .A(\DRAM_mem[29][16] ), .B(n1155), .S(n2239), .Z(n1237) );
  MUX2_X1 U2158 ( .A(\DRAM_mem[29][15] ), .B(n1156), .S(n2239), .Z(n1236) );
  MUX2_X1 U2159 ( .A(\DRAM_mem[29][14] ), .B(n2181), .S(n2239), .Z(n1235) );
  MUX2_X1 U2160 ( .A(\DRAM_mem[29][13] ), .B(n2182), .S(n2239), .Z(n1234) );
  MUX2_X1 U2161 ( .A(\DRAM_mem[29][12] ), .B(n2183), .S(n2239), .Z(n1233) );
  MUX2_X1 U2162 ( .A(\DRAM_mem[29][11] ), .B(n2184), .S(n2239), .Z(n1232) );
  MUX2_X1 U2163 ( .A(\DRAM_mem[29][10] ), .B(n2185), .S(n2239), .Z(n1231) );
  MUX2_X1 U2164 ( .A(\DRAM_mem[29][9] ), .B(n2186), .S(n2239), .Z(n1230) );
  MUX2_X1 U2165 ( .A(\DRAM_mem[29][8] ), .B(n2187), .S(n2239), .Z(n1229) );
  MUX2_X1 U2166 ( .A(\DRAM_mem[29][7] ), .B(n2188), .S(n2239), .Z(n1228) );
  MUX2_X1 U2167 ( .A(\DRAM_mem[29][6] ), .B(n2189), .S(n2239), .Z(n1227) );
  MUX2_X1 U2168 ( .A(\DRAM_mem[29][5] ), .B(n2190), .S(n2239), .Z(n1226) );
  MUX2_X1 U2169 ( .A(\DRAM_mem[29][4] ), .B(n2191), .S(n2239), .Z(n1225) );
  MUX2_X1 U2170 ( .A(\DRAM_mem[29][3] ), .B(n2192), .S(n2239), .Z(n1224) );
  MUX2_X1 U2171 ( .A(\DRAM_mem[29][2] ), .B(n2193), .S(n2239), .Z(n1223) );
  MUX2_X1 U2172 ( .A(\DRAM_mem[29][1] ), .B(n2194), .S(n2239), .Z(n1222) );
  MUX2_X1 U2173 ( .A(\DRAM_mem[29][0] ), .B(n2195), .S(n2239), .Z(n1221) );
  AND3_X1 U2174 ( .A1(Addr[0]), .A2(n2236), .A3(n113), .ZN(n2207) );
  INV_X1 U2175 ( .A(Addr[1]), .ZN(n2236) );
  MUX2_X1 U2176 ( .A(\DRAM_mem[30][31] ), .B(n1139), .S(n2240), .Z(n1220) );
  MUX2_X1 U2177 ( .A(\DRAM_mem[30][30] ), .B(n1141), .S(n2240), .Z(n1219) );
  MUX2_X1 U2178 ( .A(\DRAM_mem[30][29] ), .B(n1142), .S(n2240), .Z(n1218) );
  MUX2_X1 U2179 ( .A(\DRAM_mem[30][28] ), .B(n1143), .S(n2240), .Z(n1217) );
  MUX2_X1 U2180 ( .A(\DRAM_mem[30][27] ), .B(n1144), .S(n2240), .Z(n1216) );
  MUX2_X1 U2181 ( .A(\DRAM_mem[30][26] ), .B(n1145), .S(n2240), .Z(n1215) );
  MUX2_X1 U2182 ( .A(\DRAM_mem[30][25] ), .B(n1146), .S(n2240), .Z(n1214) );
  MUX2_X1 U2183 ( .A(\DRAM_mem[30][24] ), .B(n1147), .S(n2240), .Z(n1213) );
  MUX2_X1 U2184 ( .A(\DRAM_mem[30][23] ), .B(n1148), .S(n2240), .Z(n1212) );
  MUX2_X1 U2185 ( .A(\DRAM_mem[30][22] ), .B(n1149), .S(n2240), .Z(n1211) );
  MUX2_X1 U2186 ( .A(\DRAM_mem[30][21] ), .B(n1150), .S(n2240), .Z(n1210) );
  MUX2_X1 U2187 ( .A(\DRAM_mem[30][20] ), .B(n1151), .S(n2240), .Z(n1209) );
  MUX2_X1 U2188 ( .A(\DRAM_mem[30][19] ), .B(n1152), .S(n2240), .Z(n1208) );
  MUX2_X1 U2189 ( .A(\DRAM_mem[30][18] ), .B(n1153), .S(n2240), .Z(n1207) );
  MUX2_X1 U2190 ( .A(\DRAM_mem[30][17] ), .B(n1154), .S(n2240), .Z(n1206) );
  MUX2_X1 U2191 ( .A(\DRAM_mem[30][16] ), .B(n1155), .S(n2240), .Z(n1205) );
  MUX2_X1 U2192 ( .A(\DRAM_mem[30][15] ), .B(n1156), .S(n2240), .Z(n1204) );
  MUX2_X1 U2193 ( .A(\DRAM_mem[30][14] ), .B(n2181), .S(n2240), .Z(n1203) );
  MUX2_X1 U2194 ( .A(\DRAM_mem[30][13] ), .B(n2182), .S(n2240), .Z(n1202) );
  MUX2_X1 U2195 ( .A(\DRAM_mem[30][12] ), .B(n2183), .S(n2240), .Z(n1201) );
  MUX2_X1 U2196 ( .A(\DRAM_mem[30][11] ), .B(n2184), .S(n2240), .Z(n1200) );
  MUX2_X1 U2197 ( .A(\DRAM_mem[30][10] ), .B(n2185), .S(n2240), .Z(n1199) );
  MUX2_X1 U2198 ( .A(\DRAM_mem[30][9] ), .B(n2186), .S(n2240), .Z(n1198) );
  MUX2_X1 U2199 ( .A(\DRAM_mem[30][8] ), .B(n2187), .S(n2240), .Z(n1197) );
  MUX2_X1 U2200 ( .A(\DRAM_mem[30][7] ), .B(n2188), .S(n2240), .Z(n1196) );
  MUX2_X1 U2201 ( .A(\DRAM_mem[30][6] ), .B(n2189), .S(n2240), .Z(n1195) );
  MUX2_X1 U2202 ( .A(\DRAM_mem[30][5] ), .B(n2190), .S(n2240), .Z(n1194) );
  MUX2_X1 U2203 ( .A(\DRAM_mem[30][4] ), .B(n2191), .S(n2240), .Z(n1193) );
  MUX2_X1 U2204 ( .A(\DRAM_mem[30][3] ), .B(n2192), .S(n2240), .Z(n1192) );
  MUX2_X1 U2205 ( .A(\DRAM_mem[30][2] ), .B(n2193), .S(n2240), .Z(n1191) );
  MUX2_X1 U2206 ( .A(\DRAM_mem[30][1] ), .B(n2194), .S(n2240), .Z(n1190) );
  MUX2_X1 U2207 ( .A(\DRAM_mem[30][0] ), .B(n2195), .S(n2240), .Z(n1189) );
  AND3_X1 U2208 ( .A1(Addr[1]), .A2(n2234), .A3(n113), .ZN(n2209) );
  INV_X1 U2209 ( .A(Addr[0]), .ZN(n2234) );
  MUX2_X1 U2210 ( .A(\DRAM_mem[31][31] ), .B(n1139), .S(n2241), .Z(n1188) );
  INV_X1 U2211 ( .A(n2242), .ZN(n1139) );
  OAI21_X1 U2212 ( .B1(Din[31]), .B2(n2243), .A(n2244), .ZN(n2242) );
  MUX2_X1 U2213 ( .A(\DRAM_mem[31][30] ), .B(n1141), .S(n2241), .Z(n1187) );
  INV_X1 U2214 ( .A(n2245), .ZN(n1141) );
  OAI21_X1 U2215 ( .B1(Din[30]), .B2(n2243), .A(n2244), .ZN(n2245) );
  MUX2_X1 U2216 ( .A(\DRAM_mem[31][29] ), .B(n1142), .S(n2241), .Z(n1186) );
  INV_X1 U2217 ( .A(n2246), .ZN(n1142) );
  OAI21_X1 U2218 ( .B1(Din[29]), .B2(n2243), .A(n2244), .ZN(n2246) );
  MUX2_X1 U2219 ( .A(\DRAM_mem[31][28] ), .B(n1143), .S(n2241), .Z(n1185) );
  INV_X1 U2220 ( .A(n2247), .ZN(n1143) );
  OAI21_X1 U2221 ( .B1(Din[28]), .B2(n2243), .A(n2244), .ZN(n2247) );
  MUX2_X1 U2222 ( .A(\DRAM_mem[31][27] ), .B(n1144), .S(n2241), .Z(n1184) );
  INV_X1 U2223 ( .A(n2248), .ZN(n1144) );
  OAI21_X1 U2224 ( .B1(Din[27]), .B2(n2243), .A(n2244), .ZN(n2248) );
  MUX2_X1 U2225 ( .A(\DRAM_mem[31][26] ), .B(n1145), .S(n2241), .Z(n1183) );
  INV_X1 U2226 ( .A(n2249), .ZN(n1145) );
  OAI21_X1 U2227 ( .B1(Din[26]), .B2(n2243), .A(n2244), .ZN(n2249) );
  MUX2_X1 U2228 ( .A(\DRAM_mem[31][25] ), .B(n1146), .S(n2241), .Z(n1182) );
  INV_X1 U2229 ( .A(n2250), .ZN(n1146) );
  OAI21_X1 U2230 ( .B1(Din[25]), .B2(n2243), .A(n2244), .ZN(n2250) );
  MUX2_X1 U2231 ( .A(\DRAM_mem[31][24] ), .B(n1147), .S(n2241), .Z(n1181) );
  INV_X1 U2232 ( .A(n2251), .ZN(n1147) );
  OAI21_X1 U2233 ( .B1(Din[24]), .B2(n2243), .A(n2244), .ZN(n2251) );
  MUX2_X1 U2234 ( .A(\DRAM_mem[31][23] ), .B(n1148), .S(n2241), .Z(n1180) );
  INV_X1 U2235 ( .A(n2252), .ZN(n1148) );
  OAI21_X1 U2236 ( .B1(Din[23]), .B2(n2243), .A(n2244), .ZN(n2252) );
  MUX2_X1 U2237 ( .A(\DRAM_mem[31][22] ), .B(n1149), .S(n2241), .Z(n1179) );
  INV_X1 U2238 ( .A(n2253), .ZN(n1149) );
  OAI21_X1 U2239 ( .B1(Din[22]), .B2(n2243), .A(n2244), .ZN(n2253) );
  MUX2_X1 U2240 ( .A(\DRAM_mem[31][21] ), .B(n1150), .S(n2241), .Z(n1178) );
  INV_X1 U2241 ( .A(n2254), .ZN(n1150) );
  OAI21_X1 U2242 ( .B1(Din[21]), .B2(n2243), .A(n2244), .ZN(n2254) );
  MUX2_X1 U2243 ( .A(\DRAM_mem[31][20] ), .B(n1151), .S(n2241), .Z(n1177) );
  INV_X1 U2244 ( .A(n2255), .ZN(n1151) );
  OAI21_X1 U2245 ( .B1(Din[20]), .B2(n2243), .A(n2244), .ZN(n2255) );
  MUX2_X1 U2246 ( .A(\DRAM_mem[31][19] ), .B(n1152), .S(n2241), .Z(n1176) );
  INV_X1 U2247 ( .A(n2256), .ZN(n1152) );
  OAI21_X1 U2248 ( .B1(Din[19]), .B2(n2243), .A(n2244), .ZN(n2256) );
  MUX2_X1 U2249 ( .A(\DRAM_mem[31][18] ), .B(n1153), .S(n2241), .Z(n1175) );
  INV_X1 U2250 ( .A(n2257), .ZN(n1153) );
  OAI21_X1 U2251 ( .B1(Din[18]), .B2(n2243), .A(n2244), .ZN(n2257) );
  MUX2_X1 U2252 ( .A(\DRAM_mem[31][17] ), .B(n1154), .S(n2241), .Z(n1174) );
  INV_X1 U2253 ( .A(n2258), .ZN(n1154) );
  OAI21_X1 U2254 ( .B1(Din[17]), .B2(n2243), .A(n2244), .ZN(n2258) );
  MUX2_X1 U2255 ( .A(\DRAM_mem[31][16] ), .B(n1155), .S(n2241), .Z(n1173) );
  INV_X1 U2256 ( .A(n2259), .ZN(n1155) );
  OAI21_X1 U2257 ( .B1(Din[16]), .B2(n2243), .A(n2244), .ZN(n2259) );
  MUX2_X1 U2258 ( .A(\DRAM_mem[31][15] ), .B(n1156), .S(n2241), .Z(n1172) );
  INV_X1 U2259 ( .A(n2260), .ZN(n1156) );
  OAI21_X1 U2260 ( .B1(Din[15]), .B2(n2243), .A(n2244), .ZN(n2260) );
  NAND2_X1 U2261 ( .A1(n2261), .A2(n2262), .ZN(n2244) );
  INV_X1 U2262 ( .A(n2261), .ZN(n2243) );
  AOI21_X1 U2263 ( .B1(n2263), .B2(Din[15]), .A(n2264), .ZN(n2261) );
  MUX2_X1 U2264 ( .A(\DRAM_mem[31][14] ), .B(n2181), .S(n2241), .Z(n1171) );
  INV_X1 U2265 ( .A(n2265), .ZN(n2181) );
  OAI21_X1 U2266 ( .B1(Din[14]), .B2(n2264), .A(n2266), .ZN(n2265) );
  MUX2_X1 U2267 ( .A(\DRAM_mem[31][13] ), .B(n2182), .S(n2241), .Z(n1170) );
  INV_X1 U2268 ( .A(n2267), .ZN(n2182) );
  OAI21_X1 U2269 ( .B1(Din[13]), .B2(n2264), .A(n2266), .ZN(n2267) );
  MUX2_X1 U2270 ( .A(\DRAM_mem[31][12] ), .B(n2183), .S(n2241), .Z(n1169) );
  INV_X1 U2271 ( .A(n2268), .ZN(n2183) );
  OAI21_X1 U2272 ( .B1(Din[12]), .B2(n2264), .A(n2266), .ZN(n2268) );
  MUX2_X1 U2273 ( .A(\DRAM_mem[31][11] ), .B(n2184), .S(n2241), .Z(n1168) );
  INV_X1 U2274 ( .A(n2269), .ZN(n2184) );
  OAI21_X1 U2275 ( .B1(Din[11]), .B2(n2264), .A(n2266), .ZN(n2269) );
  MUX2_X1 U2276 ( .A(\DRAM_mem[31][10] ), .B(n2185), .S(n2241), .Z(n1167) );
  INV_X1 U2277 ( .A(n2270), .ZN(n2185) );
  OAI21_X1 U2278 ( .B1(Din[10]), .B2(n2264), .A(n2266), .ZN(n2270) );
  MUX2_X1 U2279 ( .A(\DRAM_mem[31][9] ), .B(n2186), .S(n2241), .Z(n1166) );
  INV_X1 U2280 ( .A(n2271), .ZN(n2186) );
  OAI21_X1 U2281 ( .B1(Din[9]), .B2(n2264), .A(n2266), .ZN(n2271) );
  MUX2_X1 U2282 ( .A(\DRAM_mem[31][8] ), .B(n2187), .S(n2241), .Z(n1165) );
  INV_X1 U2283 ( .A(n2272), .ZN(n2187) );
  OAI21_X1 U2284 ( .B1(Din[8]), .B2(n2264), .A(n2266), .ZN(n2272) );
  NAND2_X1 U2285 ( .A1(n2273), .A2(n2274), .ZN(n2266) );
  INV_X1 U2286 ( .A(n2274), .ZN(n2264) );
  NAND2_X1 U2287 ( .A1(Din[7]), .A2(n2275), .ZN(n2274) );
  MUX2_X1 U2288 ( .A(\DRAM_mem[31][7] ), .B(n2188), .S(n2241), .Z(n1164) );
  AND2_X1 U2289 ( .A1(Din[7]), .A2(n2276), .ZN(n2188) );
  MUX2_X1 U2290 ( .A(\DRAM_mem[31][6] ), .B(n2189), .S(n2241), .Z(n1163) );
  AND2_X1 U2291 ( .A1(Din[6]), .A2(n2276), .ZN(n2189) );
  MUX2_X1 U2292 ( .A(\DRAM_mem[31][5] ), .B(n2190), .S(n2241), .Z(n1162) );
  AND2_X1 U2293 ( .A1(Din[5]), .A2(n2276), .ZN(n2190) );
  MUX2_X1 U2294 ( .A(\DRAM_mem[31][4] ), .B(n2191), .S(n2241), .Z(n1161) );
  AND2_X1 U2295 ( .A1(Din[4]), .A2(n2276), .ZN(n2191) );
  MUX2_X1 U2296 ( .A(\DRAM_mem[31][3] ), .B(n2192), .S(n2241), .Z(n1160) );
  AND2_X1 U2297 ( .A1(Din[3]), .A2(n2276), .ZN(n2192) );
  MUX2_X1 U2298 ( .A(\DRAM_mem[31][2] ), .B(n2193), .S(n2241), .Z(n1159) );
  AND2_X1 U2299 ( .A1(Din[2]), .A2(n2276), .ZN(n2193) );
  MUX2_X1 U2300 ( .A(\DRAM_mem[31][1] ), .B(n2194), .S(n2241), .Z(n1158) );
  AND2_X1 U2301 ( .A1(Din[1]), .A2(n2276), .ZN(n2194) );
  MUX2_X1 U2302 ( .A(\DRAM_mem[31][0] ), .B(n2195), .S(n2241), .Z(n1157) );
  AND3_X1 U2303 ( .A1(Addr[1]), .A2(Addr[0]), .A3(n113), .ZN(n2211) );
  AND3_X1 U2304 ( .A1(Addr[3]), .A2(n2212), .A3(n163), .ZN(n2232) );
  AND2_X1 U2305 ( .A1(WM), .A2(EN), .ZN(n2212) );
  AND2_X1 U2306 ( .A1(Din[0]), .A2(n2276), .ZN(n2195) );
  NAND2_X1 U2307 ( .A1(n2273), .A2(n2277), .ZN(n2276) );
  INV_X1 U2308 ( .A(n2275), .ZN(n2277) );
  AND2_X1 U2309 ( .A1(RM), .A2(EN), .ZN(N598) );
  OAI21_X1 U2310 ( .B1(n2262), .B2(n2278), .A(n2279), .ZN(N597) );
  INV_X1 U2311 ( .A(N386), .ZN(n2278) );
  OAI21_X1 U2312 ( .B1(n2262), .B2(n2280), .A(n2279), .ZN(N596) );
  INV_X1 U2313 ( .A(N387), .ZN(n2280) );
  OAI21_X1 U2314 ( .B1(n2262), .B2(n2281), .A(n2279), .ZN(N595) );
  INV_X1 U2315 ( .A(N388), .ZN(n2281) );
  OAI21_X1 U2316 ( .B1(n2262), .B2(n2282), .A(n2279), .ZN(N594) );
  INV_X1 U2317 ( .A(N389), .ZN(n2282) );
  OAI21_X1 U2318 ( .B1(n2262), .B2(n2283), .A(n2279), .ZN(N593) );
  INV_X1 U2319 ( .A(N390), .ZN(n2283) );
  OAI21_X1 U2320 ( .B1(n2262), .B2(n2284), .A(n2279), .ZN(N592) );
  INV_X1 U2321 ( .A(N391), .ZN(n2284) );
  OAI21_X1 U2322 ( .B1(n2262), .B2(n2285), .A(n2279), .ZN(N591) );
  INV_X1 U2323 ( .A(N392), .ZN(n2285) );
  OAI21_X1 U2324 ( .B1(n2262), .B2(n2286), .A(n2279), .ZN(N590) );
  INV_X1 U2325 ( .A(N393), .ZN(n2286) );
  OAI21_X1 U2326 ( .B1(n2262), .B2(n2287), .A(n2279), .ZN(N589) );
  INV_X1 U2327 ( .A(N394), .ZN(n2287) );
  OAI21_X1 U2328 ( .B1(n2262), .B2(n2288), .A(n2279), .ZN(N588) );
  INV_X1 U2329 ( .A(N395), .ZN(n2288) );
  OAI21_X1 U2330 ( .B1(n2262), .B2(n2289), .A(n2279), .ZN(N587) );
  INV_X1 U2331 ( .A(N396), .ZN(n2289) );
  OAI21_X1 U2332 ( .B1(n2262), .B2(n2290), .A(n2279), .ZN(N586) );
  INV_X1 U2333 ( .A(N397), .ZN(n2290) );
  OAI21_X1 U2334 ( .B1(n2262), .B2(n2291), .A(n2279), .ZN(N585) );
  INV_X1 U2335 ( .A(N398), .ZN(n2291) );
  OAI21_X1 U2336 ( .B1(n2262), .B2(n2292), .A(n2279), .ZN(N584) );
  INV_X1 U2337 ( .A(N399), .ZN(n2292) );
  OAI21_X1 U2338 ( .B1(n2262), .B2(n2293), .A(n2279), .ZN(N583) );
  INV_X1 U2339 ( .A(N400), .ZN(n2293) );
  OAI21_X1 U2340 ( .B1(n2262), .B2(n2294), .A(n2279), .ZN(N582) );
  INV_X1 U2341 ( .A(N401), .ZN(n2294) );
  INV_X1 U2342 ( .A(n2296), .ZN(n2262) );
  INV_X1 U2343 ( .A(n2297), .ZN(N581) );
  AOI21_X1 U2344 ( .B1(n2298), .B2(N484), .A(n2295), .ZN(n2297) );
  INV_X1 U2345 ( .A(n2299), .ZN(N580) );
  AOI21_X1 U2346 ( .B1(n2298), .B2(N485), .A(n2295), .ZN(n2299) );
  INV_X1 U2347 ( .A(n2300), .ZN(N579) );
  AOI21_X1 U2348 ( .B1(n2298), .B2(N486), .A(n2295), .ZN(n2300) );
  INV_X1 U2349 ( .A(n2301), .ZN(N578) );
  AOI21_X1 U2350 ( .B1(n2298), .B2(N487), .A(n2295), .ZN(n2301) );
  INV_X1 U2351 ( .A(n2302), .ZN(N577) );
  AOI21_X1 U2352 ( .B1(n2298), .B2(N488), .A(n2295), .ZN(n2302) );
  INV_X1 U2353 ( .A(n2303), .ZN(N576) );
  AOI21_X1 U2354 ( .B1(n2298), .B2(N489), .A(n2295), .ZN(n2303) );
  INV_X1 U2355 ( .A(n2304), .ZN(N575) );
  AOI21_X1 U2356 ( .B1(n2298), .B2(N490), .A(n2295), .ZN(n2304) );
  INV_X1 U2357 ( .A(n2305), .ZN(N574) );
  AOI21_X1 U2358 ( .B1(n2298), .B2(N491), .A(n2295), .ZN(n2305) );
  AND2_X1 U2359 ( .A1(N492), .A2(n2275), .ZN(n2295) );
  NOR3_X1 U2360 ( .A1(Sel[1]), .A2(Sel[2]), .A3(n2306), .ZN(n2275) );
  INV_X1 U2361 ( .A(Sel[0]), .ZN(n2306) );
  OAI21_X1 U2362 ( .B1(Sel[0]), .B2(Sel[1]), .A(n2273), .ZN(n2298) );
  NOR2_X1 U2363 ( .A1(n2296), .A2(n2263), .ZN(n2273) );
  NOR3_X1 U2364 ( .A1(Sel[0]), .A2(Sel[2]), .A3(n2307), .ZN(n2263) );
  INV_X1 U2365 ( .A(Sel[1]), .ZN(n2307) );
  NOR3_X1 U2366 ( .A1(Sel[1]), .A2(Sel[2]), .A3(Sel[0]), .ZN(n2296) );
  AND2_X1 U2367 ( .A1(n2308), .A2(N492), .ZN(N573) );
  AND2_X1 U2368 ( .A1(N493), .A2(n2308), .ZN(N572) );
  AND2_X1 U2369 ( .A1(N494), .A2(n2308), .ZN(N571) );
  AND2_X1 U2370 ( .A1(N495), .A2(n2308), .ZN(N570) );
  AND2_X1 U2371 ( .A1(N496), .A2(n2308), .ZN(N569) );
  AND2_X1 U2372 ( .A1(N497), .A2(n2308), .ZN(N568) );
  AND2_X1 U2373 ( .A1(N498), .A2(n2308), .ZN(N567) );
  AND2_X1 U2374 ( .A1(N499), .A2(n2308), .ZN(N566) );
  OAI21_X1 U2375 ( .B1(Sel[1]), .B2(Sel[0]), .A(Sel[2]), .ZN(n2308) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_96 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_95 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_94 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_93 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_92 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_91 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_90 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_89 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_88 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_87 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_86 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_85 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_84 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_83 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_82 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_81 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_80 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_79 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_78 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_77 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_76 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_75 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_74 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_73 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_72 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_71 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_70 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_69 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_68 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_67 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_66 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_65 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_64 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_63 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_62 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_61 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_60 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_59 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_58 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_57 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_56 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_55 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_54 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_53 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_52 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_51 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_50 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_49 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_48 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_47 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_46 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_45 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_44 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_43 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_42 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_41 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_40 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_39 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_38 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_37 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_36 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_35 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_34 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_33 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module MEMU_N32 ( CLK, RST, RM, WM, EN3, S3, S4, MEM_CFG, ALU_OUT, regBout, 
        NPC2in, RD3in, RD3out, WB_DATA );
  input [2:0] MEM_CFG;
  input [31:0] ALU_OUT;
  input [31:0] regBout;
  input [31:0] NPC2in;
  input [4:0] RD3in;
  output [4:0] RD3out;
  output [31:0] WB_DATA;
  input CLK, RST, RM, WM, EN3, S3, S4;

  wire   [31:0] DataMemOut;
  wire   [31:0] wb_prime;
  assign RD3out[4] = RD3in[4];
  assign RD3out[3] = RD3in[3];
  assign RD3out[2] = RD3in[2];
  assign RD3out[1] = RD3in[1];
  assign RD3out[0] = RD3in[0];

  DataMemory_RAM_DEPTH32_WORD_SIZE32 DRAM ( .Rst(RST), .Addr(ALU_OUT), .Din(
        regBout), .Dout(DataMemOut), .Sel(MEM_CFG), .RM(RM), .WM(WM), .EN(EN3), 
        .CLK(CLK) );
  MUX21_GENERIC_NBIT32_2 MUX21_ALMEM ( .A(DataMemOut), .B(ALU_OUT), .SEL(S3), 
        .Y(wb_prime) );
  MUX21_GENERIC_NBIT32_1 MUX21_NPCWB ( .A(NPC2in), .B(wb_prime), .SEL(S4), .Y(
        WB_DATA) );
endmodule


module dlx ( RST, CLK );
  input RST, CLK;
  wire   stall, PC_EN, jump;
  wire   [31:0] IR_IN_CTRL;
  wire   [4:0] rd1_in;
  wire   [4:0] rd1_out;
  wire   [4:0] cw_dec;
  wire   [10:0] cw_ex;
  wire   [8:0] cw_mem;
  wire   [31:0] alu_out;
  wire   [31:0] IR_OUT;
  wire   [31:0] NPC_OUT;
  wire   [4:0] wr_address;
  wire   [31:0] wr_data;
  wire   [31:0] npc1_out;
  wire   [31:0] rega_out;
  wire   [31:0] regb_out;
  wire   [31:0] imm_out;
  wire   [31:0] aluout_regn;
  wire   [31:0] bout_regn;
  wire   [31:0] npc2_out;
  wire   [4:0] rd2out;

  dlx_cu unit_control ( .Clk(CLK), .Rst(RST), .IR_IN(IR_IN_CTRL), 
        .IR_OUT_OPCODE(IR_OUT[31:26]), .RD1_IN(rd1_in), .RD1_OUT(rd1_out), 
        .CW_DECODE(cw_dec), .CW_EXE(cw_ex), .CW_MEMWB(cw_mem), .FETCH_STALL(
        stall) );
  FU_N32 unit_fetch ( .IR_En(PC_EN), .PC_En(PC_EN), .NPC_En(PC_EN), .Clk(CLK), 
        .RST(RST), .COND_REGOUT(jump), .FLUSH(stall), .ALU_OUT(alu_out), 
        .IR_IN(IR_IN_CTRL), .IR_OUT(IR_OUT), .NPC_OUT(NPC_OUT) );
  DU_N32 unit_decode ( .IR_IN(IR_OUT), .NPC(NPC_OUT), .WR_ADDR_RF(wr_address), 
        .DATAIN(wr_data), .EN1(cw_dec[2]), .RF1(cw_dec[4]), .RF2(cw_dec[3]), 
        .WF1(cw_mem[4]), .CLK(CLK), .RST(RST), .SEL_IMM(cw_dec[1:0]), 
        .NPC1_OUT(npc1_out), .regA_OUT(rega_out), .regB_OUT(regb_out), 
        .IMM_OUT(imm_out), .RD1_IN(rd1_in), .RD1_OUT(rd1_out) );
  EXUNIT_N32 unit_execution ( .NPC1(npc1_out), .RD1(rd1_out), .A(rega_out), 
        .B(regb_out), .IMM(imm_out), .S1_A_NPC(cw_ex[10]), .S2_IMM_B(cw_ex[9]), 
        .ALU_OPCODE(cw_ex[5:0]), .CLK(CLK), .RST(RST), .JUMP_EN(cw_ex[7:6]), 
        .EN_REGN_ALU_OUT(cw_ex[8]), .JUMP(jump), .ALUOUT(alu_out), 
        .ALU_OUT_REGN(aluout_regn), .B_OUT_REGN(bout_regn), .NPC2(npc2_out), 
        .RD2_OUT_REGN(rd2out) );
  MEMU_N32 unit_memory ( .CLK(CLK), .RST(RST), .RM(cw_mem[8]), .WM(cw_mem[7]), 
        .EN3(cw_mem[5]), .S3(cw_mem[6]), .S4(cw_mem[3]), .MEM_CFG(cw_mem[2:0]), 
        .ALU_OUT(aluout_regn), .regBout(bout_regn), .NPC2in(npc2_out), .RD3in(
        rd2out), .RD3out(wr_address), .WB_DATA(wr_data) );
  INV_X4 U4 ( .A(stall), .ZN(PC_EN) );
endmodule

