library IEEE;
use IEEE.std_logic_1164.all; 
use WORK.constants.all; 

entity tb is
end tb;

architecture test of tb is
component is
	GENERIC ();
	PORT();
end component;

begin
	
	uut:
	
	process
	begin
	end process;
end test;

