

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Level1 is
  Port ( );
end Level1;

architecture Beh of Level1 is

begin


end Beh;
