package CONSTANTS is
   constant IVDELAY : time := 0.0 ns;
   constant NDDELAY : time := 0.0 ns;
   constant NDDELAYRISE : time := 0.0 ns;
   constant NDDELAYFALL : time := 0.0 ns;
   constant NRDELAY : time := 0.0 ns;
   constant DRCAS : time := 0.0 ns;
   constant DRCAC : time := 0.0 ns;
   constant NumBit : integer := 16;	
   constant NumBitBlock: integer := 2;
   constant TP_MUX : time := 0.0 ns; 	
end CONSTANTS;
