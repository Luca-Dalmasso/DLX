
module DataMemory_RAM_DEPTH32_WORD_SIZE32 ( Rst, Addr, Din, Dout, Sel, RM, WM, 
        EN, CLK );
  input [31:0] Addr;
  input [31:0] Din;
  output [31:0] Dout;
  input [2:0] Sel;
  input Rst, RM, WM, EN, CLK;
  wire   N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576,
         N577, N578, N579, N580, N581, N598, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n13687, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540;

  DLH_X1 \Dout_reg[31]  ( .G(N598), .D(n7404), .Q(Dout[31]) );
  DLH_X1 \Dout_reg[30]  ( .G(N598), .D(n7403), .Q(Dout[30]) );
  DLH_X1 \Dout_reg[29]  ( .G(N598), .D(n7402), .Q(Dout[29]) );
  DLH_X1 \Dout_reg[28]  ( .G(N598), .D(n7401), .Q(Dout[28]) );
  DLH_X1 \Dout_reg[27]  ( .G(N598), .D(n7400), .Q(Dout[27]) );
  DLH_X1 \Dout_reg[26]  ( .G(N598), .D(n7399), .Q(Dout[26]) );
  DLH_X1 \Dout_reg[25]  ( .G(N598), .D(n7398), .Q(Dout[25]) );
  DLH_X1 \Dout_reg[24]  ( .G(N598), .D(n7397), .Q(Dout[24]) );
  DLH_X1 \Dout_reg[23]  ( .G(N598), .D(n7396), .Q(Dout[23]) );
  DLH_X1 \Dout_reg[22]  ( .G(N598), .D(n7395), .Q(Dout[22]) );
  DLH_X1 \Dout_reg[21]  ( .G(N598), .D(n7394), .Q(Dout[21]) );
  DLH_X1 \Dout_reg[20]  ( .G(N598), .D(n7393), .Q(Dout[20]) );
  DLH_X1 \Dout_reg[19]  ( .G(N598), .D(n7392), .Q(Dout[19]) );
  DLH_X1 \Dout_reg[18]  ( .G(N598), .D(n7391), .Q(Dout[18]) );
  DLH_X1 \Dout_reg[17]  ( .G(N598), .D(n7390), .Q(Dout[17]) );
  DLH_X1 \Dout_reg[16]  ( .G(N598), .D(n7389), .Q(Dout[16]) );
  DLH_X1 \Dout_reg[15]  ( .G(N598), .D(N581), .Q(Dout[15]) );
  DLH_X1 \Dout_reg[14]  ( .G(N598), .D(N580), .Q(Dout[14]) );
  DLH_X1 \Dout_reg[13]  ( .G(N598), .D(N579), .Q(Dout[13]) );
  DLH_X1 \Dout_reg[12]  ( .G(N598), .D(N578), .Q(Dout[12]) );
  DLH_X1 \Dout_reg[11]  ( .G(N598), .D(N577), .Q(Dout[11]) );
  DLH_X1 \Dout_reg[10]  ( .G(N598), .D(N576), .Q(Dout[10]) );
  DLH_X1 \Dout_reg[9]  ( .G(N598), .D(N575), .Q(Dout[9]) );
  DLH_X1 \Dout_reg[8]  ( .G(N598), .D(N574), .Q(Dout[8]) );
  DLH_X1 \Dout_reg[7]  ( .G(N598), .D(N573), .Q(Dout[7]) );
  DLH_X1 \Dout_reg[6]  ( .G(N598), .D(N572), .Q(Dout[6]) );
  DLH_X1 \Dout_reg[5]  ( .G(N598), .D(N571), .Q(Dout[5]) );
  DLH_X1 \Dout_reg[4]  ( .G(N598), .D(N570), .Q(Dout[4]) );
  DLH_X1 \Dout_reg[3]  ( .G(N598), .D(N569), .Q(Dout[3]) );
  DLH_X1 \Dout_reg[2]  ( .G(N598), .D(N568), .Q(Dout[2]) );
  DLH_X1 \Dout_reg[1]  ( .G(N598), .D(N567), .Q(Dout[1]) );
  DLH_X1 \Dout_reg[0]  ( .G(N598), .D(N566), .Q(Dout[0]) );
  DFFR_X1 \DRAM_mem_reg[0][31]  ( .D(n2213), .CK(CLK), .RN(n945), .Q(n3039), 
        .QN(n457) );
  DFFR_X1 \DRAM_mem_reg[0][30]  ( .D(n2212), .CK(CLK), .RN(n945), .Q(n3040), 
        .QN(n458) );
  DFFR_X1 \DRAM_mem_reg[0][29]  ( .D(n2211), .CK(CLK), .RN(n945), .Q(n3041), 
        .QN(n459) );
  DFFR_X1 \DRAM_mem_reg[0][28]  ( .D(n2210), .CK(CLK), .RN(n945), .Q(n3042), 
        .QN(n460) );
  DFFR_X1 \DRAM_mem_reg[0][27]  ( .D(n2209), .CK(CLK), .RN(n945), .Q(n3043), 
        .QN(n461) );
  DFFR_X1 \DRAM_mem_reg[0][26]  ( .D(n2208), .CK(CLK), .RN(n945), .Q(n3044), 
        .QN(n462) );
  DFFR_X1 \DRAM_mem_reg[0][25]  ( .D(n2207), .CK(CLK), .RN(n945), .Q(n3045), 
        .QN(n463) );
  DFFR_X1 \DRAM_mem_reg[0][24]  ( .D(n2206), .CK(CLK), .RN(n945), .Q(n3046), 
        .QN(n464) );
  DFFR_X1 \DRAM_mem_reg[0][23]  ( .D(n2205), .CK(CLK), .RN(n945), .Q(n3047), 
        .QN(n465) );
  DFFR_X1 \DRAM_mem_reg[0][22]  ( .D(n2204), .CK(CLK), .RN(n945), .Q(n3048), 
        .QN(n466) );
  DFFR_X1 \DRAM_mem_reg[0][21]  ( .D(n2203), .CK(CLK), .RN(n945), .Q(n3049), 
        .QN(n467) );
  DFFR_X1 \DRAM_mem_reg[0][20]  ( .D(n2202), .CK(CLK), .RN(n945), .Q(n3050), 
        .QN(n468) );
  DFFR_X1 \DRAM_mem_reg[0][19]  ( .D(n2201), .CK(CLK), .RN(n946), .Q(n3051), 
        .QN(n469) );
  DFFR_X1 \DRAM_mem_reg[0][18]  ( .D(n2200), .CK(CLK), .RN(n946), .Q(n3052), 
        .QN(n470) );
  DFFR_X1 \DRAM_mem_reg[0][17]  ( .D(n2199), .CK(CLK), .RN(n946), .Q(n3053), 
        .QN(n471) );
  DFFR_X1 \DRAM_mem_reg[0][16]  ( .D(n2198), .CK(CLK), .RN(n946), .Q(n3054), 
        .QN(n472) );
  DFFR_X1 \DRAM_mem_reg[0][15]  ( .D(n2197), .CK(CLK), .RN(n946), .Q(n126) );
  DFFR_X1 \DRAM_mem_reg[0][14]  ( .D(n2196), .CK(CLK), .RN(n946), .Q(n3055), 
        .QN(n431) );
  DFFR_X1 \DRAM_mem_reg[0][13]  ( .D(n2195), .CK(CLK), .RN(n946), .Q(n3056), 
        .QN(n435) );
  DFFR_X1 \DRAM_mem_reg[0][12]  ( .D(n2194), .CK(CLK), .RN(n946), .Q(n3057), 
        .QN(n439) );
  DFFR_X1 \DRAM_mem_reg[0][11]  ( .D(n2193), .CK(CLK), .RN(n946), .Q(n3058), 
        .QN(n443) );
  DFFR_X1 \DRAM_mem_reg[0][10]  ( .D(n2192), .CK(CLK), .RN(n946), .Q(n3059), 
        .QN(n447) );
  DFFR_X1 \DRAM_mem_reg[0][9]  ( .D(n2191), .CK(CLK), .RN(n946), .Q(n3060), 
        .QN(n451) );
  DFFR_X1 \DRAM_mem_reg[0][8]  ( .D(n2190), .CK(CLK), .RN(n946), .Q(n3061), 
        .QN(n455) );
  DFFR_X1 \DRAM_mem_reg[0][7]  ( .D(n2189), .CK(CLK), .RN(n947), .Q(n825), 
        .QN(n3062) );
  DFFR_X1 \DRAM_mem_reg[0][6]  ( .D(n2188), .CK(CLK), .RN(n947), .Q(n826), 
        .QN(n3063) );
  DFFR_X1 \DRAM_mem_reg[0][5]  ( .D(n2187), .CK(CLK), .RN(n947), .Q(n827), 
        .QN(n3064) );
  DFFR_X1 \DRAM_mem_reg[0][4]  ( .D(n2186), .CK(CLK), .RN(n947), .Q(n828), 
        .QN(n3065) );
  DFFR_X1 \DRAM_mem_reg[0][3]  ( .D(n2185), .CK(CLK), .RN(n947), .Q(n829), 
        .QN(n3066) );
  DFFR_X1 \DRAM_mem_reg[0][2]  ( .D(n2184), .CK(CLK), .RN(n947), .Q(n830), 
        .QN(n3067) );
  DFFR_X1 \DRAM_mem_reg[0][1]  ( .D(n2183), .CK(CLK), .RN(n947), .Q(n831), 
        .QN(n3068) );
  DFFR_X1 \DRAM_mem_reg[0][0]  ( .D(n2182), .CK(CLK), .RN(n947), .Q(n832), 
        .QN(n3069) );
  DFFR_X1 \DRAM_mem_reg[1][31]  ( .D(n2181), .CK(CLK), .RN(n947), .Q(n2885), 
        .QN(n205) );
  DFFR_X1 \DRAM_mem_reg[1][30]  ( .D(n2180), .CK(CLK), .RN(n947), .Q(n2886), 
        .QN(n206) );
  DFFR_X1 \DRAM_mem_reg[1][29]  ( .D(n2179), .CK(CLK), .RN(n947), .Q(n2887), 
        .QN(n207) );
  DFFR_X1 \DRAM_mem_reg[1][28]  ( .D(n2178), .CK(CLK), .RN(n947), .Q(n2888), 
        .QN(n208) );
  DFFR_X1 \DRAM_mem_reg[1][27]  ( .D(n2177), .CK(CLK), .RN(n948), .Q(n2889), 
        .QN(n209) );
  DFFR_X1 \DRAM_mem_reg[1][26]  ( .D(n2176), .CK(CLK), .RN(n948), .Q(n2890), 
        .QN(n210) );
  DFFR_X1 \DRAM_mem_reg[1][25]  ( .D(n2175), .CK(CLK), .RN(n948), .Q(n2891), 
        .QN(n211) );
  DFFR_X1 \DRAM_mem_reg[1][24]  ( .D(n2174), .CK(CLK), .RN(n948), .Q(n2892), 
        .QN(n212) );
  DFFR_X1 \DRAM_mem_reg[1][23]  ( .D(n2173), .CK(CLK), .RN(n948), .Q(n2893), 
        .QN(n213) );
  DFFR_X1 \DRAM_mem_reg[1][22]  ( .D(n2172), .CK(CLK), .RN(n948), .Q(n2894), 
        .QN(n214) );
  DFFR_X1 \DRAM_mem_reg[1][21]  ( .D(n2171), .CK(CLK), .RN(n948), .Q(n2895), 
        .QN(n215) );
  DFFR_X1 \DRAM_mem_reg[1][20]  ( .D(n2170), .CK(CLK), .RN(n948), .Q(n2896), 
        .QN(n216) );
  DFFR_X1 \DRAM_mem_reg[1][19]  ( .D(n2169), .CK(CLK), .RN(n948), .Q(n2897), 
        .QN(n217) );
  DFFR_X1 \DRAM_mem_reg[1][18]  ( .D(n2168), .CK(CLK), .RN(n948), .Q(n2898), 
        .QN(n218) );
  DFFR_X1 \DRAM_mem_reg[1][17]  ( .D(n2167), .CK(CLK), .RN(n948), .Q(n2899), 
        .QN(n219) );
  DFFR_X1 \DRAM_mem_reg[1][16]  ( .D(n2166), .CK(CLK), .RN(n948), .Q(n2900), 
        .QN(n220) );
  DFFR_X1 \DRAM_mem_reg[1][15]  ( .D(n2165), .CK(CLK), .RN(n949), .Q(n124) );
  DFFR_X1 \DRAM_mem_reg[1][14]  ( .D(n2164), .CK(CLK), .RN(n949), .Q(n3070), 
        .QN(n179) );
  DFFR_X1 \DRAM_mem_reg[1][13]  ( .D(n2163), .CK(CLK), .RN(n949), .Q(n3071), 
        .QN(n183) );
  DFFR_X1 \DRAM_mem_reg[1][12]  ( .D(n2162), .CK(CLK), .RN(n949), .Q(n3072), 
        .QN(n187) );
  DFFR_X1 \DRAM_mem_reg[1][11]  ( .D(n2161), .CK(CLK), .RN(n949), .Q(n3073), 
        .QN(n191) );
  DFFR_X1 \DRAM_mem_reg[1][10]  ( .D(n2160), .CK(CLK), .RN(n949), .Q(n3074), 
        .QN(n195) );
  DFFR_X1 \DRAM_mem_reg[1][9]  ( .D(n2159), .CK(CLK), .RN(n949), .Q(n3075), 
        .QN(n199) );
  DFFR_X1 \DRAM_mem_reg[1][8]  ( .D(n2158), .CK(CLK), .RN(n949), .Q(n3076), 
        .QN(n203) );
  DFFR_X1 \DRAM_mem_reg[1][7]  ( .D(n2157), .CK(CLK), .RN(n949), .Q(n721), 
        .QN(n3077) );
  DFFR_X1 \DRAM_mem_reg[1][6]  ( .D(n2156), .CK(CLK), .RN(n949), .Q(n722), 
        .QN(n3078) );
  DFFR_X1 \DRAM_mem_reg[1][5]  ( .D(n2155), .CK(CLK), .RN(n949), .Q(n723), 
        .QN(n3079) );
  DFFR_X1 \DRAM_mem_reg[1][4]  ( .D(n2154), .CK(CLK), .RN(n949), .Q(n724), 
        .QN(n3080) );
  DFFR_X1 \DRAM_mem_reg[1][3]  ( .D(n2153), .CK(CLK), .RN(n950), .Q(n725), 
        .QN(n3081) );
  DFFR_X1 \DRAM_mem_reg[1][2]  ( .D(n2152), .CK(CLK), .RN(n950), .Q(n726), 
        .QN(n3082) );
  DFFR_X1 \DRAM_mem_reg[1][1]  ( .D(n2151), .CK(CLK), .RN(n950), .Q(n727), 
        .QN(n3083) );
  DFFR_X1 \DRAM_mem_reg[1][0]  ( .D(n2150), .CK(CLK), .RN(n950), .Q(n728), 
        .QN(n3084) );
  DFFR_X1 \DRAM_mem_reg[2][31]  ( .D(n2149), .CK(CLK), .RN(n950), .Q(n2901) );
  DFFR_X1 \DRAM_mem_reg[2][30]  ( .D(n2148), .CK(CLK), .RN(n950), .Q(n2902) );
  DFFR_X1 \DRAM_mem_reg[2][29]  ( .D(n2147), .CK(CLK), .RN(n950), .Q(n2903) );
  DFFR_X1 \DRAM_mem_reg[2][28]  ( .D(n2146), .CK(CLK), .RN(n950), .Q(n2904) );
  DFFR_X1 \DRAM_mem_reg[2][27]  ( .D(n2145), .CK(CLK), .RN(n950), .Q(n2905) );
  DFFR_X1 \DRAM_mem_reg[2][26]  ( .D(n2144), .CK(CLK), .RN(n950), .Q(n2906) );
  DFFR_X1 \DRAM_mem_reg[2][25]  ( .D(n2143), .CK(CLK), .RN(n950), .Q(n2907) );
  DFFR_X1 \DRAM_mem_reg[2][24]  ( .D(n2142), .CK(CLK), .RN(n950), .Q(n2908) );
  DFFR_X1 \DRAM_mem_reg[2][23]  ( .D(n2141), .CK(CLK), .RN(n951), .Q(n2909) );
  DFFR_X1 \DRAM_mem_reg[2][22]  ( .D(n2140), .CK(CLK), .RN(n951), .Q(n2910) );
  DFFR_X1 \DRAM_mem_reg[2][21]  ( .D(n2139), .CK(CLK), .RN(n951), .Q(n2911) );
  DFFR_X1 \DRAM_mem_reg[2][20]  ( .D(n2138), .CK(CLK), .RN(n951), .Q(n2912) );
  DFFR_X1 \DRAM_mem_reg[2][19]  ( .D(n2137), .CK(CLK), .RN(n951), .Q(n2913) );
  DFFR_X1 \DRAM_mem_reg[2][18]  ( .D(n2136), .CK(CLK), .RN(n951), .Q(n2914) );
  DFFR_X1 \DRAM_mem_reg[2][17]  ( .D(n2135), .CK(CLK), .RN(n951), .Q(n2915) );
  DFFR_X1 \DRAM_mem_reg[2][16]  ( .D(n2134), .CK(CLK), .RN(n951), .Q(n2916) );
  DFFR_X1 \DRAM_mem_reg[2][15]  ( .D(n2133), .CK(CLK), .RN(n951), .Q(n122) );
  DFFR_X1 \DRAM_mem_reg[2][14]  ( .D(n2132), .CK(CLK), .RN(n951), .Q(n21) );
  DFFR_X1 \DRAM_mem_reg[2][13]  ( .D(n2131), .CK(CLK), .RN(n951), .Q(n29) );
  DFFR_X1 \DRAM_mem_reg[2][12]  ( .D(n2130), .CK(CLK), .RN(n951), .Q(n37) );
  DFFR_X1 \DRAM_mem_reg[2][11]  ( .D(n2129), .CK(CLK), .RN(n952), .Q(n45) );
  DFFR_X1 \DRAM_mem_reg[2][10]  ( .D(n2128), .CK(CLK), .RN(n952), .Q(n53) );
  DFFR_X1 \DRAM_mem_reg[2][9]  ( .D(n2127), .CK(CLK), .RN(n952), .Q(n61) );
  DFFR_X1 \DRAM_mem_reg[2][8]  ( .D(n2126), .CK(CLK), .RN(n952), .Q(n69) );
  DFFR_X1 \DRAM_mem_reg[2][7]  ( .D(n2125), .CK(CLK), .RN(n952), .Q(n2976) );
  DFFR_X1 \DRAM_mem_reg[2][6]  ( .D(n2124), .CK(CLK), .RN(n952), .Q(n2984) );
  DFFR_X1 \DRAM_mem_reg[2][5]  ( .D(n2123), .CK(CLK), .RN(n952), .Q(n2992) );
  DFFR_X1 \DRAM_mem_reg[2][4]  ( .D(n2122), .CK(CLK), .RN(n952), .Q(n3000) );
  DFFR_X1 \DRAM_mem_reg[2][3]  ( .D(n2121), .CK(CLK), .RN(n952), .Q(n3008) );
  DFFR_X1 \DRAM_mem_reg[2][2]  ( .D(n2120), .CK(CLK), .RN(n952), .Q(n3016) );
  DFFR_X1 \DRAM_mem_reg[2][1]  ( .D(n2119), .CK(CLK), .RN(n952), .Q(n3024) );
  DFFR_X1 \DRAM_mem_reg[2][0]  ( .D(n2118), .CK(CLK), .RN(n952), .Q(n3032) );
  DFFR_X1 \DRAM_mem_reg[3][31]  ( .D(n2117), .CK(CLK), .RN(n953), .Q(n161) );
  DFFR_X1 \DRAM_mem_reg[3][30]  ( .D(n2116), .CK(CLK), .RN(n953), .Q(n162) );
  DFFR_X1 \DRAM_mem_reg[3][29]  ( .D(n2115), .CK(CLK), .RN(n953), .Q(n163) );
  DFFR_X1 \DRAM_mem_reg[3][28]  ( .D(n2114), .CK(CLK), .RN(n953), .Q(n164) );
  DFFR_X1 \DRAM_mem_reg[3][27]  ( .D(n2113), .CK(CLK), .RN(n953), .Q(n165) );
  DFFR_X1 \DRAM_mem_reg[3][26]  ( .D(n2112), .CK(CLK), .RN(n953), .Q(n166) );
  DFFR_X1 \DRAM_mem_reg[3][25]  ( .D(n2111), .CK(CLK), .RN(n953), .Q(n167) );
  DFFR_X1 \DRAM_mem_reg[3][24]  ( .D(n2110), .CK(CLK), .RN(n953), .Q(n168) );
  DFFR_X1 \DRAM_mem_reg[3][23]  ( .D(n2109), .CK(CLK), .RN(n953), .Q(n169) );
  DFFR_X1 \DRAM_mem_reg[3][22]  ( .D(n2108), .CK(CLK), .RN(n953), .Q(n170) );
  DFFR_X1 \DRAM_mem_reg[3][21]  ( .D(n2107), .CK(CLK), .RN(n953), .Q(n171) );
  DFFR_X1 \DRAM_mem_reg[3][20]  ( .D(n2106), .CK(CLK), .RN(n953), .Q(n172) );
  DFFR_X1 \DRAM_mem_reg[3][19]  ( .D(n2105), .CK(CLK), .RN(n954), .Q(n173) );
  DFFR_X1 \DRAM_mem_reg[3][18]  ( .D(n2104), .CK(CLK), .RN(n954), .Q(n174) );
  DFFR_X1 \DRAM_mem_reg[3][17]  ( .D(n2103), .CK(CLK), .RN(n954), .Q(n175) );
  DFFR_X1 \DRAM_mem_reg[3][16]  ( .D(n2102), .CK(CLK), .RN(n954), .Q(n176) );
  DFFR_X1 \DRAM_mem_reg[3][15]  ( .D(n2101), .CK(CLK), .RN(n954), .Q(n128) );
  DFFR_X1 \DRAM_mem_reg[3][14]  ( .D(n2100), .CK(CLK), .RN(n954), .Q(n257) );
  DFFR_X1 \DRAM_mem_reg[3][13]  ( .D(n2099), .CK(CLK), .RN(n954), .Q(n265) );
  DFFR_X1 \DRAM_mem_reg[3][12]  ( .D(n2098), .CK(CLK), .RN(n954), .Q(n273) );
  DFFR_X1 \DRAM_mem_reg[3][11]  ( .D(n2097), .CK(CLK), .RN(n954), .Q(n281) );
  DFFR_X1 \DRAM_mem_reg[3][10]  ( .D(n2096), .CK(CLK), .RN(n954), .Q(n289) );
  DFFR_X1 \DRAM_mem_reg[3][9]  ( .D(n2095), .CK(CLK), .RN(n954), .Q(n297) );
  DFFR_X1 \DRAM_mem_reg[3][8]  ( .D(n2094), .CK(CLK), .RN(n954), .Q(n305) );
  DFFR_X1 \DRAM_mem_reg[3][7]  ( .D(n2093), .CK(CLK), .RN(n955), .Q(n2975) );
  DFFR_X1 \DRAM_mem_reg[3][6]  ( .D(n2092), .CK(CLK), .RN(n955), .Q(n2983) );
  DFFR_X1 \DRAM_mem_reg[3][5]  ( .D(n2091), .CK(CLK), .RN(n955), .Q(n2991) );
  DFFR_X1 \DRAM_mem_reg[3][4]  ( .D(n2090), .CK(CLK), .RN(n955), .Q(n2999) );
  DFFR_X1 \DRAM_mem_reg[3][3]  ( .D(n2089), .CK(CLK), .RN(n955), .Q(n3007) );
  DFFR_X1 \DRAM_mem_reg[3][2]  ( .D(n2088), .CK(CLK), .RN(n955), .Q(n3015) );
  DFFR_X1 \DRAM_mem_reg[3][1]  ( .D(n2087), .CK(CLK), .RN(n955), .Q(n3023) );
  DFFR_X1 \DRAM_mem_reg[3][0]  ( .D(n2086), .CK(CLK), .RN(n955), .Q(n3031) );
  DFFR_X1 \DRAM_mem_reg[4][31]  ( .D(n2085), .CK(CLK), .RN(n955), .Q(n73) );
  DFFR_X1 \DRAM_mem_reg[4][30]  ( .D(n2084), .CK(CLK), .RN(n955), .Q(n74) );
  DFFR_X1 \DRAM_mem_reg[4][29]  ( .D(n2083), .CK(CLK), .RN(n955), .Q(n75) );
  DFFR_X1 \DRAM_mem_reg[4][28]  ( .D(n2082), .CK(CLK), .RN(n955), .Q(n76) );
  DFFR_X1 \DRAM_mem_reg[4][27]  ( .D(n2081), .CK(CLK), .RN(n956), .Q(n77) );
  DFFR_X1 \DRAM_mem_reg[4][26]  ( .D(n2080), .CK(CLK), .RN(n956), .Q(n78) );
  DFFR_X1 \DRAM_mem_reg[4][25]  ( .D(n2079), .CK(CLK), .RN(n956), .Q(n79) );
  DFFR_X1 \DRAM_mem_reg[4][24]  ( .D(n2078), .CK(CLK), .RN(n956), .Q(n80) );
  DFFR_X1 \DRAM_mem_reg[4][23]  ( .D(n2077), .CK(CLK), .RN(n956), .Q(n81) );
  DFFR_X1 \DRAM_mem_reg[4][22]  ( .D(n2076), .CK(CLK), .RN(n956), .Q(n82) );
  DFFR_X1 \DRAM_mem_reg[4][21]  ( .D(n2075), .CK(CLK), .RN(n956), .Q(n83) );
  DFFR_X1 \DRAM_mem_reg[4][20]  ( .D(n2074), .CK(CLK), .RN(n956), .Q(n84) );
  DFFR_X1 \DRAM_mem_reg[4][19]  ( .D(n2073), .CK(CLK), .RN(n956), .Q(n85) );
  DFFR_X1 \DRAM_mem_reg[4][18]  ( .D(n2072), .CK(CLK), .RN(n956), .Q(n86) );
  DFFR_X1 \DRAM_mem_reg[4][17]  ( .D(n2071), .CK(CLK), .RN(n956), .Q(n87) );
  DFFR_X1 \DRAM_mem_reg[4][16]  ( .D(n2070), .CK(CLK), .RN(n956), .Q(n88) );
  DFFR_X1 \DRAM_mem_reg[4][15]  ( .D(n2069), .CK(CLK), .RN(n957), .Q(n362) );
  DFFR_X1 \DRAM_mem_reg[4][14]  ( .D(n2068), .CK(CLK), .RN(n957), .Q(n2938), 
        .QN(n432) );
  DFFR_X1 \DRAM_mem_reg[4][13]  ( .D(n2067), .CK(CLK), .RN(n957), .Q(n2944), 
        .QN(n436) );
  DFFR_X1 \DRAM_mem_reg[4][12]  ( .D(n2066), .CK(CLK), .RN(n957), .Q(n2950), 
        .QN(n440) );
  DFFR_X1 \DRAM_mem_reg[4][11]  ( .D(n2065), .CK(CLK), .RN(n957), .Q(n2956), 
        .QN(n444) );
  DFFR_X1 \DRAM_mem_reg[4][10]  ( .D(n2064), .CK(CLK), .RN(n957), .Q(n2962), 
        .QN(n448) );
  DFFR_X1 \DRAM_mem_reg[4][9]  ( .D(n2063), .CK(CLK), .RN(n957), .Q(n2968), 
        .QN(n452) );
  DFFR_X1 \DRAM_mem_reg[4][8]  ( .D(n2062), .CK(CLK), .RN(n957), .Q(n2974), 
        .QN(n456) );
  DFFR_X1 \DRAM_mem_reg[4][7]  ( .D(n2061), .CK(CLK), .RN(n957), .Q(n833), 
        .QN(n3085) );
  DFFR_X1 \DRAM_mem_reg[4][6]  ( .D(n2060), .CK(CLK), .RN(n957), .Q(n834), 
        .QN(n3086) );
  DFFR_X1 \DRAM_mem_reg[4][5]  ( .D(n2059), .CK(CLK), .RN(n957), .Q(n835), 
        .QN(n3087) );
  DFFR_X1 \DRAM_mem_reg[4][4]  ( .D(n2058), .CK(CLK), .RN(n957), .Q(n836), 
        .QN(n3088) );
  DFFR_X1 \DRAM_mem_reg[4][3]  ( .D(n2057), .CK(CLK), .RN(n958), .Q(n837), 
        .QN(n3089) );
  DFFR_X1 \DRAM_mem_reg[4][2]  ( .D(n2056), .CK(CLK), .RN(n958), .Q(n838), 
        .QN(n3090) );
  DFFR_X1 \DRAM_mem_reg[4][1]  ( .D(n2055), .CK(CLK), .RN(n958), .Q(n839), 
        .QN(n3091) );
  DFFR_X1 \DRAM_mem_reg[4][0]  ( .D(n2054), .CK(CLK), .RN(n958), .Q(n840), 
        .QN(n3092) );
  DFFR_X1 \DRAM_mem_reg[5][31]  ( .D(n2053), .CK(CLK), .RN(n958), .Q(n397) );
  DFFR_X1 \DRAM_mem_reg[5][30]  ( .D(n2052), .CK(CLK), .RN(n958), .Q(n398) );
  DFFR_X1 \DRAM_mem_reg[5][29]  ( .D(n2051), .CK(CLK), .RN(n958), .Q(n399) );
  DFFR_X1 \DRAM_mem_reg[5][28]  ( .D(n2050), .CK(CLK), .RN(n958), .Q(n400) );
  DFFR_X1 \DRAM_mem_reg[5][27]  ( .D(n2049), .CK(CLK), .RN(n958), .Q(n401) );
  DFFR_X1 \DRAM_mem_reg[5][26]  ( .D(n2048), .CK(CLK), .RN(n958), .Q(n402) );
  DFFR_X1 \DRAM_mem_reg[5][25]  ( .D(n2047), .CK(CLK), .RN(n958), .Q(n403) );
  DFFR_X1 \DRAM_mem_reg[5][24]  ( .D(n2046), .CK(CLK), .RN(n958), .Q(n404) );
  DFFR_X1 \DRAM_mem_reg[5][23]  ( .D(n2045), .CK(CLK), .RN(n959), .Q(n405) );
  DFFR_X1 \DRAM_mem_reg[5][22]  ( .D(n2044), .CK(CLK), .RN(n959), .Q(n406) );
  DFFR_X1 \DRAM_mem_reg[5][21]  ( .D(n2043), .CK(CLK), .RN(n959), .Q(n407) );
  DFFR_X1 \DRAM_mem_reg[5][20]  ( .D(n2042), .CK(CLK), .RN(n959), .Q(n408) );
  DFFR_X1 \DRAM_mem_reg[5][19]  ( .D(n2041), .CK(CLK), .RN(n959), .Q(n409) );
  DFFR_X1 \DRAM_mem_reg[5][18]  ( .D(n2040), .CK(CLK), .RN(n959), .Q(n410) );
  DFFR_X1 \DRAM_mem_reg[5][17]  ( .D(n2039), .CK(CLK), .RN(n959), .Q(n411) );
  DFFR_X1 \DRAM_mem_reg[5][16]  ( .D(n2038), .CK(CLK), .RN(n959), .Q(n412) );
  DFFR_X1 \DRAM_mem_reg[5][15]  ( .D(n2037), .CK(CLK), .RN(n959), .Q(n360) );
  DFFR_X1 \DRAM_mem_reg[5][14]  ( .D(n2036), .CK(CLK), .RN(n959), .Q(n2937), 
        .QN(n180) );
  DFFR_X1 \DRAM_mem_reg[5][13]  ( .D(n2035), .CK(CLK), .RN(n959), .Q(n2943), 
        .QN(n184) );
  DFFR_X1 \DRAM_mem_reg[5][12]  ( .D(n2034), .CK(CLK), .RN(n959), .Q(n2949), 
        .QN(n188) );
  DFFR_X1 \DRAM_mem_reg[5][11]  ( .D(n2033), .CK(CLK), .RN(n960), .Q(n2955), 
        .QN(n192) );
  DFFR_X1 \DRAM_mem_reg[5][10]  ( .D(n2032), .CK(CLK), .RN(n960), .Q(n2961), 
        .QN(n196) );
  DFFR_X1 \DRAM_mem_reg[5][9]  ( .D(n2031), .CK(CLK), .RN(n960), .Q(n2967), 
        .QN(n200) );
  DFFR_X1 \DRAM_mem_reg[5][8]  ( .D(n2030), .CK(CLK), .RN(n960), .Q(n2973), 
        .QN(n204) );
  DFFR_X1 \DRAM_mem_reg[5][7]  ( .D(n2029), .CK(CLK), .RN(n960), .Q(n729), 
        .QN(n3093) );
  DFFR_X1 \DRAM_mem_reg[5][6]  ( .D(n2028), .CK(CLK), .RN(n960), .Q(n730), 
        .QN(n3094) );
  DFFR_X1 \DRAM_mem_reg[5][5]  ( .D(n2027), .CK(CLK), .RN(n960), .Q(n731), 
        .QN(n3095) );
  DFFR_X1 \DRAM_mem_reg[5][4]  ( .D(n2026), .CK(CLK), .RN(n960), .Q(n732), 
        .QN(n3096) );
  DFFR_X1 \DRAM_mem_reg[5][3]  ( .D(n2025), .CK(CLK), .RN(n960), .Q(n733), 
        .QN(n3097) );
  DFFR_X1 \DRAM_mem_reg[5][2]  ( .D(n2024), .CK(CLK), .RN(n960), .Q(n734), 
        .QN(n3098) );
  DFFR_X1 \DRAM_mem_reg[5][1]  ( .D(n2023), .CK(CLK), .RN(n960), .Q(n735), 
        .QN(n3099) );
  DFFR_X1 \DRAM_mem_reg[5][0]  ( .D(n2022), .CK(CLK), .RN(n960), .Q(n736), 
        .QN(n3100) );
  DFFR_X1 \DRAM_mem_reg[6][31]  ( .D(n2021), .CK(CLK), .RN(n961), .Q(n309) );
  DFFR_X1 \DRAM_mem_reg[6][30]  ( .D(n2020), .CK(CLK), .RN(n961), .Q(n310) );
  DFFR_X1 \DRAM_mem_reg[6][29]  ( .D(n2019), .CK(CLK), .RN(n961), .Q(n311) );
  DFFR_X1 \DRAM_mem_reg[6][28]  ( .D(n2018), .CK(CLK), .RN(n961), .Q(n312) );
  DFFR_X1 \DRAM_mem_reg[6][27]  ( .D(n2017), .CK(CLK), .RN(n961), .Q(n313) );
  DFFR_X1 \DRAM_mem_reg[6][26]  ( .D(n2016), .CK(CLK), .RN(n961), .Q(n314) );
  DFFR_X1 \DRAM_mem_reg[6][25]  ( .D(n2015), .CK(CLK), .RN(n961), .Q(n315) );
  DFFR_X1 \DRAM_mem_reg[6][24]  ( .D(n2014), .CK(CLK), .RN(n961), .Q(n316) );
  DFFR_X1 \DRAM_mem_reg[6][23]  ( .D(n2013), .CK(CLK), .RN(n961), .Q(n317) );
  DFFR_X1 \DRAM_mem_reg[6][22]  ( .D(n2012), .CK(CLK), .RN(n961), .Q(n318) );
  DFFR_X1 \DRAM_mem_reg[6][21]  ( .D(n2011), .CK(CLK), .RN(n961), .Q(n319) );
  DFFR_X1 \DRAM_mem_reg[6][20]  ( .D(n2010), .CK(CLK), .RN(n961), .Q(n320) );
  DFFR_X1 \DRAM_mem_reg[6][19]  ( .D(n2009), .CK(CLK), .RN(n962), .Q(n321) );
  DFFR_X1 \DRAM_mem_reg[6][18]  ( .D(n2008), .CK(CLK), .RN(n962), .Q(n322) );
  DFFR_X1 \DRAM_mem_reg[6][17]  ( .D(n2007), .CK(CLK), .RN(n962), .Q(n323) );
  DFFR_X1 \DRAM_mem_reg[6][16]  ( .D(n2006), .CK(CLK), .RN(n962), .Q(n324) );
  DFFR_X1 \DRAM_mem_reg[6][15]  ( .D(n2005), .CK(CLK), .RN(n962), .Q(n358) );
  DFFR_X1 \DRAM_mem_reg[6][14]  ( .D(n2004), .CK(CLK), .RN(n962), .Q(n22) );
  DFFR_X1 \DRAM_mem_reg[6][13]  ( .D(n2003), .CK(CLK), .RN(n962), .Q(n30) );
  DFFR_X1 \DRAM_mem_reg[6][12]  ( .D(n2002), .CK(CLK), .RN(n962), .Q(n38) );
  DFFR_X1 \DRAM_mem_reg[6][11]  ( .D(n2001), .CK(CLK), .RN(n962), .Q(n46) );
  DFFR_X1 \DRAM_mem_reg[6][10]  ( .D(n2000), .CK(CLK), .RN(n962), .Q(n54) );
  DFFR_X1 \DRAM_mem_reg[6][9]  ( .D(n1999), .CK(CLK), .RN(n962), .Q(n62) );
  DFFR_X1 \DRAM_mem_reg[6][8]  ( .D(n1998), .CK(CLK), .RN(n962), .Q(n70) );
  DFFR_X1 \DRAM_mem_reg[6][7]  ( .D(n1997), .CK(CLK), .RN(n963), .Q(n2978) );
  DFFR_X1 \DRAM_mem_reg[6][6]  ( .D(n1996), .CK(CLK), .RN(n963), .Q(n2986) );
  DFFR_X1 \DRAM_mem_reg[6][5]  ( .D(n1995), .CK(CLK), .RN(n963), .Q(n2994) );
  DFFR_X1 \DRAM_mem_reg[6][4]  ( .D(n1994), .CK(CLK), .RN(n963), .Q(n3002) );
  DFFR_X1 \DRAM_mem_reg[6][3]  ( .D(n1993), .CK(CLK), .RN(n963), .Q(n3010) );
  DFFR_X1 \DRAM_mem_reg[6][2]  ( .D(n1992), .CK(CLK), .RN(n963), .Q(n3018) );
  DFFR_X1 \DRAM_mem_reg[6][1]  ( .D(n1991), .CK(CLK), .RN(n963), .Q(n3026) );
  DFFR_X1 \DRAM_mem_reg[6][0]  ( .D(n1990), .CK(CLK), .RN(n963), .Q(n3034) );
  DFFR_X1 \DRAM_mem_reg[7][31]  ( .D(n1989), .CK(CLK), .RN(n963), .Q(n2917), 
        .QN(n413) );
  DFFR_X1 \DRAM_mem_reg[7][30]  ( .D(n1988), .CK(CLK), .RN(n963), .Q(n2918), 
        .QN(n414) );
  DFFR_X1 \DRAM_mem_reg[7][29]  ( .D(n1987), .CK(CLK), .RN(n963), .Q(n2919), 
        .QN(n415) );
  DFFR_X1 \DRAM_mem_reg[7][28]  ( .D(n1986), .CK(CLK), .RN(n963), .Q(n2920), 
        .QN(n416) );
  DFFR_X1 \DRAM_mem_reg[7][27]  ( .D(n1985), .CK(CLK), .RN(n964), .Q(n2921), 
        .QN(n417) );
  DFFR_X1 \DRAM_mem_reg[7][26]  ( .D(n1984), .CK(CLK), .RN(n964), .Q(n2922), 
        .QN(n418) );
  DFFR_X1 \DRAM_mem_reg[7][25]  ( .D(n1983), .CK(CLK), .RN(n964), .Q(n2923), 
        .QN(n419) );
  DFFR_X1 \DRAM_mem_reg[7][24]  ( .D(n1982), .CK(CLK), .RN(n964), .Q(n2924), 
        .QN(n420) );
  DFFR_X1 \DRAM_mem_reg[7][23]  ( .D(n1981), .CK(CLK), .RN(n964), .Q(n2925), 
        .QN(n421) );
  DFFR_X1 \DRAM_mem_reg[7][22]  ( .D(n1980), .CK(CLK), .RN(n964), .Q(n2926), 
        .QN(n422) );
  DFFR_X1 \DRAM_mem_reg[7][21]  ( .D(n1979), .CK(CLK), .RN(n964), .Q(n2927), 
        .QN(n423) );
  DFFR_X1 \DRAM_mem_reg[7][20]  ( .D(n1978), .CK(CLK), .RN(n964), .Q(n2928), 
        .QN(n424) );
  DFFR_X1 \DRAM_mem_reg[7][19]  ( .D(n1977), .CK(CLK), .RN(n964), .Q(n2929), 
        .QN(n425) );
  DFFR_X1 \DRAM_mem_reg[7][18]  ( .D(n1976), .CK(CLK), .RN(n964), .Q(n2930), 
        .QN(n426) );
  DFFR_X1 \DRAM_mem_reg[7][17]  ( .D(n1975), .CK(CLK), .RN(n964), .Q(n2931), 
        .QN(n427) );
  DFFR_X1 \DRAM_mem_reg[7][16]  ( .D(n1974), .CK(CLK), .RN(n964), .Q(n2932), 
        .QN(n428) );
  DFFR_X1 \DRAM_mem_reg[7][15]  ( .D(n1973), .CK(CLK), .RN(n965), .Q(n364) );
  DFFR_X1 \DRAM_mem_reg[7][14]  ( .D(n1972), .CK(CLK), .RN(n965), .Q(n258) );
  DFFR_X1 \DRAM_mem_reg[7][13]  ( .D(n1971), .CK(CLK), .RN(n965), .Q(n266) );
  DFFR_X1 \DRAM_mem_reg[7][12]  ( .D(n1970), .CK(CLK), .RN(n965), .Q(n274) );
  DFFR_X1 \DRAM_mem_reg[7][11]  ( .D(n1969), .CK(CLK), .RN(n965), .Q(n282) );
  DFFR_X1 \DRAM_mem_reg[7][10]  ( .D(n1968), .CK(CLK), .RN(n965), .Q(n290) );
  DFFR_X1 \DRAM_mem_reg[7][9]  ( .D(n1967), .CK(CLK), .RN(n965), .Q(n298) );
  DFFR_X1 \DRAM_mem_reg[7][8]  ( .D(n1966), .CK(CLK), .RN(n965), .Q(n306) );
  DFFR_X1 \DRAM_mem_reg[7][7]  ( .D(n1965), .CK(CLK), .RN(n965), .Q(n2977) );
  DFFR_X1 \DRAM_mem_reg[7][6]  ( .D(n1964), .CK(CLK), .RN(n965), .Q(n2985) );
  DFFR_X1 \DRAM_mem_reg[7][5]  ( .D(n1963), .CK(CLK), .RN(n965), .Q(n2993) );
  DFFR_X1 \DRAM_mem_reg[7][4]  ( .D(n1962), .CK(CLK), .RN(n965), .Q(n3001) );
  DFFR_X1 \DRAM_mem_reg[7][3]  ( .D(n1961), .CK(CLK), .RN(n966), .Q(n3009) );
  DFFR_X1 \DRAM_mem_reg[7][2]  ( .D(n1960), .CK(CLK), .RN(n966), .Q(n3017) );
  DFFR_X1 \DRAM_mem_reg[7][1]  ( .D(n1959), .CK(CLK), .RN(n966), .Q(n3025) );
  DFFR_X1 \DRAM_mem_reg[7][0]  ( .D(n1958), .CK(CLK), .RN(n966), .Q(n3033) );
  DFFR_X1 \DRAM_mem_reg[8][31]  ( .D(n1957), .CK(CLK), .RN(n966), .Q(n325) );
  DFFR_X1 \DRAM_mem_reg[8][30]  ( .D(n1956), .CK(CLK), .RN(n966), .Q(n326) );
  DFFR_X1 \DRAM_mem_reg[8][29]  ( .D(n1955), .CK(CLK), .RN(n966), .Q(n327) );
  DFFR_X1 \DRAM_mem_reg[8][28]  ( .D(n1954), .CK(CLK), .RN(n966), .Q(n328) );
  DFFR_X1 \DRAM_mem_reg[8][27]  ( .D(n1953), .CK(CLK), .RN(n966), .Q(n329) );
  DFFR_X1 \DRAM_mem_reg[8][26]  ( .D(n1952), .CK(CLK), .RN(n966), .Q(n330) );
  DFFR_X1 \DRAM_mem_reg[8][25]  ( .D(n1951), .CK(CLK), .RN(n966), .Q(n331) );
  DFFR_X1 \DRAM_mem_reg[8][24]  ( .D(n1950), .CK(CLK), .RN(n966), .Q(n332) );
  DFFR_X1 \DRAM_mem_reg[8][23]  ( .D(n1949), .CK(CLK), .RN(n967), .Q(n333) );
  DFFR_X1 \DRAM_mem_reg[8][22]  ( .D(n1948), .CK(CLK), .RN(n967), .Q(n334) );
  DFFR_X1 \DRAM_mem_reg[8][21]  ( .D(n1947), .CK(CLK), .RN(n967), .Q(n335) );
  DFFR_X1 \DRAM_mem_reg[8][20]  ( .D(n1946), .CK(CLK), .RN(n967), .Q(n336) );
  DFFR_X1 \DRAM_mem_reg[8][19]  ( .D(n1945), .CK(CLK), .RN(n967), .Q(n337) );
  DFFR_X1 \DRAM_mem_reg[8][18]  ( .D(n1944), .CK(CLK), .RN(n967), .Q(n338) );
  DFFR_X1 \DRAM_mem_reg[8][17]  ( .D(n1943), .CK(CLK), .RN(n967), .Q(n339) );
  DFFR_X1 \DRAM_mem_reg[8][16]  ( .D(n1942), .CK(CLK), .RN(n967), .Q(n340) );
  DFFR_X1 \DRAM_mem_reg[8][15]  ( .D(n1941), .CK(CLK), .RN(n967), .Q(n841), 
        .QN(n3101) );
  DFFR_X1 \DRAM_mem_reg[8][14]  ( .D(n1940), .CK(CLK), .RN(n967), .Q(n24) );
  DFFR_X1 \DRAM_mem_reg[8][13]  ( .D(n1939), .CK(CLK), .RN(n967), .Q(n32) );
  DFFR_X1 \DRAM_mem_reg[8][12]  ( .D(n1938), .CK(CLK), .RN(n967), .Q(n40) );
  DFFR_X1 \DRAM_mem_reg[8][11]  ( .D(n1937), .CK(CLK), .RN(n968), .Q(n48) );
  DFFR_X1 \DRAM_mem_reg[8][10]  ( .D(n1936), .CK(CLK), .RN(n968), .Q(n56) );
  DFFR_X1 \DRAM_mem_reg[8][9]  ( .D(n1935), .CK(CLK), .RN(n968), .Q(n64) );
  DFFR_X1 \DRAM_mem_reg[8][8]  ( .D(n1934), .CK(CLK), .RN(n968), .Q(n72) );
  DFFR_X1 \DRAM_mem_reg[8][7]  ( .D(n1933), .CK(CLK), .RN(n968), .Q(n842), 
        .QN(n3102) );
  DFFR_X1 \DRAM_mem_reg[8][6]  ( .D(n1932), .CK(CLK), .RN(n968), .Q(n843), 
        .QN(n3103) );
  DFFR_X1 \DRAM_mem_reg[8][5]  ( .D(n1931), .CK(CLK), .RN(n968), .Q(n844), 
        .QN(n3104) );
  DFFR_X1 \DRAM_mem_reg[8][4]  ( .D(n1930), .CK(CLK), .RN(n968), .Q(n845), 
        .QN(n3105) );
  DFFR_X1 \DRAM_mem_reg[8][3]  ( .D(n1929), .CK(CLK), .RN(n968), .Q(n846), 
        .QN(n3106) );
  DFFR_X1 \DRAM_mem_reg[8][2]  ( .D(n1928), .CK(CLK), .RN(n968), .Q(n847), 
        .QN(n3107) );
  DFFR_X1 \DRAM_mem_reg[8][1]  ( .D(n1927), .CK(CLK), .RN(n968), .Q(n848), 
        .QN(n3108) );
  DFFR_X1 \DRAM_mem_reg[8][0]  ( .D(n1926), .CK(CLK), .RN(n968), .Q(n849), 
        .QN(n3109) );
  DFFR_X1 \DRAM_mem_reg[9][31]  ( .D(n1925), .CK(CLK), .RN(n969), .Q(n737), 
        .QN(n3110) );
  DFFR_X1 \DRAM_mem_reg[9][30]  ( .D(n1924), .CK(CLK), .RN(n969), .Q(n738), 
        .QN(n3111) );
  DFFR_X1 \DRAM_mem_reg[9][29]  ( .D(n1923), .CK(CLK), .RN(n969), .Q(n739), 
        .QN(n3112) );
  DFFR_X1 \DRAM_mem_reg[9][28]  ( .D(n1922), .CK(CLK), .RN(n969), .Q(n740), 
        .QN(n3113) );
  DFFR_X1 \DRAM_mem_reg[9][27]  ( .D(n1921), .CK(CLK), .RN(n969), .Q(n741), 
        .QN(n3114) );
  DFFR_X1 \DRAM_mem_reg[9][26]  ( .D(n1920), .CK(CLK), .RN(n969), .Q(n742), 
        .QN(n3115) );
  DFFR_X1 \DRAM_mem_reg[9][25]  ( .D(n1919), .CK(CLK), .RN(n969), .Q(n743), 
        .QN(n3116) );
  DFFR_X1 \DRAM_mem_reg[9][24]  ( .D(n1918), .CK(CLK), .RN(n969), .Q(n744), 
        .QN(n3117) );
  DFFR_X1 \DRAM_mem_reg[9][23]  ( .D(n1917), .CK(CLK), .RN(n969), .Q(n745), 
        .QN(n3118) );
  DFFR_X1 \DRAM_mem_reg[9][22]  ( .D(n1916), .CK(CLK), .RN(n969), .Q(n746), 
        .QN(n3119) );
  DFFR_X1 \DRAM_mem_reg[9][21]  ( .D(n1915), .CK(CLK), .RN(n969), .Q(n747), 
        .QN(n3120) );
  DFFR_X1 \DRAM_mem_reg[9][20]  ( .D(n1914), .CK(CLK), .RN(n969), .Q(n748), 
        .QN(n3121) );
  DFFR_X1 \DRAM_mem_reg[9][19]  ( .D(n1913), .CK(CLK), .RN(n970), .Q(n749), 
        .QN(n3122) );
  DFFR_X1 \DRAM_mem_reg[9][18]  ( .D(n1912), .CK(CLK), .RN(n970), .Q(n750), 
        .QN(n3123) );
  DFFR_X1 \DRAM_mem_reg[9][17]  ( .D(n1911), .CK(CLK), .RN(n970), .Q(n751), 
        .QN(n3124) );
  DFFR_X1 \DRAM_mem_reg[9][16]  ( .D(n1910), .CK(CLK), .RN(n970), .Q(n752), 
        .QN(n3125) );
  DFFR_X1 \DRAM_mem_reg[9][15]  ( .D(n1909), .CK(CLK), .RN(n970), .Q(n850), 
        .QN(n3126) );
  DFFR_X1 \DRAM_mem_reg[9][14]  ( .D(n1908), .CK(CLK), .RN(n970), .Q(n260) );
  DFFR_X1 \DRAM_mem_reg[9][13]  ( .D(n1907), .CK(CLK), .RN(n970), .Q(n268) );
  DFFR_X1 \DRAM_mem_reg[9][12]  ( .D(n1906), .CK(CLK), .RN(n970), .Q(n276) );
  DFFR_X1 \DRAM_mem_reg[9][11]  ( .D(n1905), .CK(CLK), .RN(n970), .Q(n284) );
  DFFR_X1 \DRAM_mem_reg[9][10]  ( .D(n1904), .CK(CLK), .RN(n970), .Q(n292) );
  DFFR_X1 \DRAM_mem_reg[9][9]  ( .D(n1903), .CK(CLK), .RN(n970), .Q(n300) );
  DFFR_X1 \DRAM_mem_reg[9][8]  ( .D(n1902), .CK(CLK), .RN(n970), .Q(n308) );
  DFFR_X1 \DRAM_mem_reg[9][7]  ( .D(n1901), .CK(CLK), .RN(n971), .Q(n753), 
        .QN(n3127) );
  DFFR_X1 \DRAM_mem_reg[9][6]  ( .D(n1900), .CK(CLK), .RN(n971), .Q(n754), 
        .QN(n3128) );
  DFFR_X1 \DRAM_mem_reg[9][5]  ( .D(n1899), .CK(CLK), .RN(n971), .Q(n755), 
        .QN(n3129) );
  DFFR_X1 \DRAM_mem_reg[9][4]  ( .D(n1898), .CK(CLK), .RN(n971), .Q(n756), 
        .QN(n3130) );
  DFFR_X1 \DRAM_mem_reg[9][3]  ( .D(n1897), .CK(CLK), .RN(n971), .Q(n757), 
        .QN(n3131) );
  DFFR_X1 \DRAM_mem_reg[9][2]  ( .D(n1896), .CK(CLK), .RN(n971), .Q(n758), 
        .QN(n3132) );
  DFFR_X1 \DRAM_mem_reg[9][1]  ( .D(n1895), .CK(CLK), .RN(n971), .Q(n759), 
        .QN(n3133) );
  DFFR_X1 \DRAM_mem_reg[9][0]  ( .D(n1894), .CK(CLK), .RN(n971), .Q(n760), 
        .QN(n3134) );
  DFFR_X1 \DRAM_mem_reg[10][31]  ( .D(n1893), .CK(CLK), .RN(n971), .Q(n89) );
  DFFR_X1 \DRAM_mem_reg[10][30]  ( .D(n1892), .CK(CLK), .RN(n971), .Q(n90) );
  DFFR_X1 \DRAM_mem_reg[10][29]  ( .D(n1891), .CK(CLK), .RN(n971), .Q(n91) );
  DFFR_X1 \DRAM_mem_reg[10][28]  ( .D(n1890), .CK(CLK), .RN(n971), .Q(n92) );
  DFFR_X1 \DRAM_mem_reg[10][27]  ( .D(n1889), .CK(CLK), .RN(n972), .Q(n93) );
  DFFR_X1 \DRAM_mem_reg[10][26]  ( .D(n1888), .CK(CLK), .RN(n972), .Q(n94) );
  DFFR_X1 \DRAM_mem_reg[10][25]  ( .D(n1887), .CK(CLK), .RN(n972), .Q(n95) );
  DFFR_X1 \DRAM_mem_reg[10][24]  ( .D(n1886), .CK(CLK), .RN(n972), .Q(n96) );
  DFFR_X1 \DRAM_mem_reg[10][23]  ( .D(n1885), .CK(CLK), .RN(n972), .Q(n97) );
  DFFR_X1 \DRAM_mem_reg[10][22]  ( .D(n1884), .CK(CLK), .RN(n972), .Q(n98) );
  DFFR_X1 \DRAM_mem_reg[10][21]  ( .D(n1883), .CK(CLK), .RN(n972), .Q(n99) );
  DFFR_X1 \DRAM_mem_reg[10][20]  ( .D(n1882), .CK(CLK), .RN(n972), .Q(n100) );
  DFFR_X1 \DRAM_mem_reg[10][19]  ( .D(n1881), .CK(CLK), .RN(n972), .Q(n101) );
  DFFR_X1 \DRAM_mem_reg[10][18]  ( .D(n1880), .CK(CLK), .RN(n972), .Q(n102) );
  DFFR_X1 \DRAM_mem_reg[10][17]  ( .D(n1879), .CK(CLK), .RN(n972), .Q(n103) );
  DFFR_X1 \DRAM_mem_reg[10][16]  ( .D(n1878), .CK(CLK), .RN(n972), .Q(n104) );
  DFFR_X1 \DRAM_mem_reg[10][15]  ( .D(n1877), .CK(CLK), .RN(n973), .Q(n851), 
        .QN(n3135) );
  DFFR_X1 \DRAM_mem_reg[10][14]  ( .D(n1876), .CK(CLK), .RN(n973), .Q(n473), 
        .QN(n3136) );
  DFFR_X1 \DRAM_mem_reg[10][13]  ( .D(n1875), .CK(CLK), .RN(n973), .Q(n474), 
        .QN(n3137) );
  DFFR_X1 \DRAM_mem_reg[10][12]  ( .D(n1874), .CK(CLK), .RN(n973), .Q(n475), 
        .QN(n3138) );
  DFFR_X1 \DRAM_mem_reg[10][11]  ( .D(n1873), .CK(CLK), .RN(n973), .Q(n476), 
        .QN(n3139) );
  DFFR_X1 \DRAM_mem_reg[10][10]  ( .D(n1872), .CK(CLK), .RN(n973), .Q(n477), 
        .QN(n3140) );
  DFFR_X1 \DRAM_mem_reg[10][9]  ( .D(n1871), .CK(CLK), .RN(n973), .Q(n478), 
        .QN(n3141) );
  DFFR_X1 \DRAM_mem_reg[10][8]  ( .D(n1870), .CK(CLK), .RN(n973), .Q(n479), 
        .QN(n3142) );
  DFFR_X1 \DRAM_mem_reg[10][7]  ( .D(n1869), .CK(CLK), .RN(n973), .Q(n365) );
  DFFR_X1 \DRAM_mem_reg[10][6]  ( .D(n1868), .CK(CLK), .RN(n973), .Q(n369) );
  DFFR_X1 \DRAM_mem_reg[10][5]  ( .D(n1867), .CK(CLK), .RN(n973), .Q(n373) );
  DFFR_X1 \DRAM_mem_reg[10][4]  ( .D(n1866), .CK(CLK), .RN(n973), .Q(n377) );
  DFFR_X1 \DRAM_mem_reg[10][3]  ( .D(n1865), .CK(CLK), .RN(n974), .Q(n381) );
  DFFR_X1 \DRAM_mem_reg[10][2]  ( .D(n1864), .CK(CLK), .RN(n974), .Q(n385) );
  DFFR_X1 \DRAM_mem_reg[10][1]  ( .D(n1863), .CK(CLK), .RN(n974), .Q(n389) );
  DFFR_X1 \DRAM_mem_reg[10][0]  ( .D(n1862), .CK(CLK), .RN(n974), .Q(n393) );
  DFFR_X1 \DRAM_mem_reg[11][31]  ( .D(n1861), .CK(CLK), .RN(n974), .Q(n852), 
        .QN(n3143) );
  DFFR_X1 \DRAM_mem_reg[11][30]  ( .D(n1860), .CK(CLK), .RN(n974), .Q(n853), 
        .QN(n3144) );
  DFFR_X1 \DRAM_mem_reg[11][29]  ( .D(n1859), .CK(CLK), .RN(n974), .Q(n854), 
        .QN(n3145) );
  DFFR_X1 \DRAM_mem_reg[11][28]  ( .D(n1858), .CK(CLK), .RN(n974), .Q(n855), 
        .QN(n3146) );
  DFFR_X1 \DRAM_mem_reg[11][27]  ( .D(n1857), .CK(CLK), .RN(n974), .Q(n856), 
        .QN(n3147) );
  DFFR_X1 \DRAM_mem_reg[11][26]  ( .D(n1856), .CK(CLK), .RN(n974), .Q(n857), 
        .QN(n3148) );
  DFFR_X1 \DRAM_mem_reg[11][25]  ( .D(n1855), .CK(CLK), .RN(n974), .Q(n858), 
        .QN(n3149) );
  DFFR_X1 \DRAM_mem_reg[11][24]  ( .D(n1854), .CK(CLK), .RN(n974), .Q(n859), 
        .QN(n3150) );
  DFFR_X1 \DRAM_mem_reg[11][23]  ( .D(n1853), .CK(CLK), .RN(n975), .Q(n860), 
        .QN(n3151) );
  DFFR_X1 \DRAM_mem_reg[11][22]  ( .D(n1852), .CK(CLK), .RN(n975), .Q(n861), 
        .QN(n3152) );
  DFFR_X1 \DRAM_mem_reg[11][21]  ( .D(n1851), .CK(CLK), .RN(n975), .Q(n862), 
        .QN(n3153) );
  DFFR_X1 \DRAM_mem_reg[11][20]  ( .D(n1850), .CK(CLK), .RN(n975), .Q(n863), 
        .QN(n3154) );
  DFFR_X1 \DRAM_mem_reg[11][19]  ( .D(n1849), .CK(CLK), .RN(n975), .Q(n864), 
        .QN(n3155) );
  DFFR_X1 \DRAM_mem_reg[11][18]  ( .D(n1848), .CK(CLK), .RN(n975), .Q(n865), 
        .QN(n3156) );
  DFFR_X1 \DRAM_mem_reg[11][17]  ( .D(n1847), .CK(CLK), .RN(n975), .Q(n866), 
        .QN(n3157) );
  DFFR_X1 \DRAM_mem_reg[11][16]  ( .D(n1846), .CK(CLK), .RN(n975), .Q(n867), 
        .QN(n3158) );
  DFFR_X1 \DRAM_mem_reg[11][15]  ( .D(n1845), .CK(CLK), .RN(n975), .Q(n868), 
        .QN(n3159) );
  DFFR_X1 \DRAM_mem_reg[11][14]  ( .D(n1844), .CK(CLK), .RN(n975), .Q(n597), 
        .QN(n3160) );
  DFFR_X1 \DRAM_mem_reg[11][13]  ( .D(n1843), .CK(CLK), .RN(n975), .Q(n598), 
        .QN(n3161) );
  DFFR_X1 \DRAM_mem_reg[11][12]  ( .D(n1842), .CK(CLK), .RN(n975), .Q(n599), 
        .QN(n3162) );
  DFFR_X1 \DRAM_mem_reg[11][11]  ( .D(n1841), .CK(CLK), .RN(n976), .Q(n600), 
        .QN(n3163) );
  DFFR_X1 \DRAM_mem_reg[11][10]  ( .D(n1840), .CK(CLK), .RN(n976), .Q(n601), 
        .QN(n3164) );
  DFFR_X1 \DRAM_mem_reg[11][9]  ( .D(n1839), .CK(CLK), .RN(n976), .Q(n602), 
        .QN(n3165) );
  DFFR_X1 \DRAM_mem_reg[11][8]  ( .D(n1838), .CK(CLK), .RN(n976), .Q(n603), 
        .QN(n3166) );
  DFFR_X1 \DRAM_mem_reg[11][7]  ( .D(n1837), .CK(CLK), .RN(n976), .Q(n129) );
  DFFR_X1 \DRAM_mem_reg[11][6]  ( .D(n1836), .CK(CLK), .RN(n976), .Q(n133) );
  DFFR_X1 \DRAM_mem_reg[11][5]  ( .D(n1835), .CK(CLK), .RN(n976), .Q(n137) );
  DFFR_X1 \DRAM_mem_reg[11][4]  ( .D(n1834), .CK(CLK), .RN(n976), .Q(n141) );
  DFFR_X1 \DRAM_mem_reg[11][3]  ( .D(n1833), .CK(CLK), .RN(n976), .Q(n145) );
  DFFR_X1 \DRAM_mem_reg[11][2]  ( .D(n1832), .CK(CLK), .RN(n976), .Q(n149) );
  DFFR_X1 \DRAM_mem_reg[11][1]  ( .D(n1831), .CK(CLK), .RN(n976), .Q(n153) );
  DFFR_X1 \DRAM_mem_reg[11][0]  ( .D(n1830), .CK(CLK), .RN(n976), .Q(n157) );
  DFFR_X1 \DRAM_mem_reg[12][31]  ( .D(n1829), .CK(CLK), .RN(n977), .Q(n105) );
  DFFR_X1 \DRAM_mem_reg[12][30]  ( .D(n1828), .CK(CLK), .RN(n977), .Q(n106) );
  DFFR_X1 \DRAM_mem_reg[12][29]  ( .D(n1827), .CK(CLK), .RN(n977), .Q(n107) );
  DFFR_X1 \DRAM_mem_reg[12][28]  ( .D(n1826), .CK(CLK), .RN(n977), .Q(n108) );
  DFFR_X1 \DRAM_mem_reg[12][27]  ( .D(n1825), .CK(CLK), .RN(n977), .Q(n109) );
  DFFR_X1 \DRAM_mem_reg[12][26]  ( .D(n1824), .CK(CLK), .RN(n977), .Q(n110) );
  DFFR_X1 \DRAM_mem_reg[12][25]  ( .D(n1823), .CK(CLK), .RN(n977), .Q(n111) );
  DFFR_X1 \DRAM_mem_reg[12][24]  ( .D(n1822), .CK(CLK), .RN(n977), .Q(n112) );
  DFFR_X1 \DRAM_mem_reg[12][23]  ( .D(n1821), .CK(CLK), .RN(n977), .Q(n113) );
  DFFR_X1 \DRAM_mem_reg[12][22]  ( .D(n1820), .CK(CLK), .RN(n977), .Q(n114) );
  DFFR_X1 \DRAM_mem_reg[12][21]  ( .D(n1819), .CK(CLK), .RN(n977), .Q(n115) );
  DFFR_X1 \DRAM_mem_reg[12][20]  ( .D(n1818), .CK(CLK), .RN(n977), .Q(n116) );
  DFFR_X1 \DRAM_mem_reg[12][19]  ( .D(n1817), .CK(CLK), .RN(n978), .Q(n117) );
  DFFR_X1 \DRAM_mem_reg[12][18]  ( .D(n1816), .CK(CLK), .RN(n978), .Q(n118) );
  DFFR_X1 \DRAM_mem_reg[12][17]  ( .D(n1815), .CK(CLK), .RN(n978), .Q(n119) );
  DFFR_X1 \DRAM_mem_reg[12][16]  ( .D(n1814), .CK(CLK), .RN(n978), .Q(n120) );
  DFFR_X1 \DRAM_mem_reg[12][15]  ( .D(n1813), .CK(CLK), .RN(n978), .Q(n761), 
        .QN(n3167) );
  DFFR_X1 \DRAM_mem_reg[12][14]  ( .D(n1812), .CK(CLK), .RN(n978), .Q(n23) );
  DFFR_X1 \DRAM_mem_reg[12][13]  ( .D(n1811), .CK(CLK), .RN(n978), .Q(n31) );
  DFFR_X1 \DRAM_mem_reg[12][12]  ( .D(n1810), .CK(CLK), .RN(n978), .Q(n39) );
  DFFR_X1 \DRAM_mem_reg[12][11]  ( .D(n1809), .CK(CLK), .RN(n978), .Q(n47) );
  DFFR_X1 \DRAM_mem_reg[12][10]  ( .D(n1808), .CK(CLK), .RN(n978), .Q(n55) );
  DFFR_X1 \DRAM_mem_reg[12][9]  ( .D(n1807), .CK(CLK), .RN(n978), .Q(n63) );
  DFFR_X1 \DRAM_mem_reg[12][8]  ( .D(n1806), .CK(CLK), .RN(n978), .Q(n71) );
  DFFR_X1 \DRAM_mem_reg[12][7]  ( .D(n1805), .CK(CLK), .RN(n979), .Q(n869), 
        .QN(n3168) );
  DFFR_X1 \DRAM_mem_reg[12][6]  ( .D(n1804), .CK(CLK), .RN(n979), .Q(n870), 
        .QN(n3169) );
  DFFR_X1 \DRAM_mem_reg[12][5]  ( .D(n1803), .CK(CLK), .RN(n979), .Q(n871), 
        .QN(n3170) );
  DFFR_X1 \DRAM_mem_reg[12][4]  ( .D(n1802), .CK(CLK), .RN(n979), .Q(n872), 
        .QN(n3171) );
  DFFR_X1 \DRAM_mem_reg[12][3]  ( .D(n1801), .CK(CLK), .RN(n979), .Q(n873), 
        .QN(n3172) );
  DFFR_X1 \DRAM_mem_reg[12][2]  ( .D(n1800), .CK(CLK), .RN(n979), .Q(n874), 
        .QN(n3173) );
  DFFR_X1 \DRAM_mem_reg[12][1]  ( .D(n1799), .CK(CLK), .RN(n979), .Q(n875), 
        .QN(n3174) );
  DFFR_X1 \DRAM_mem_reg[12][0]  ( .D(n1798), .CK(CLK), .RN(n979), .Q(n876), 
        .QN(n3175) );
  DFFR_X1 \DRAM_mem_reg[13][31]  ( .D(n1797), .CK(CLK), .RN(n979), .Q(n877), 
        .QN(n3176) );
  DFFR_X1 \DRAM_mem_reg[13][30]  ( .D(n1796), .CK(CLK), .RN(n979), .Q(n878), 
        .QN(n3177) );
  DFFR_X1 \DRAM_mem_reg[13][29]  ( .D(n1795), .CK(CLK), .RN(n979), .Q(n879), 
        .QN(n3178) );
  DFFR_X1 \DRAM_mem_reg[13][28]  ( .D(n1794), .CK(CLK), .RN(n979), .Q(n880), 
        .QN(n3179) );
  DFFR_X1 \DRAM_mem_reg[13][27]  ( .D(n1793), .CK(CLK), .RN(n980), .Q(n881), 
        .QN(n3180) );
  DFFR_X1 \DRAM_mem_reg[13][26]  ( .D(n1792), .CK(CLK), .RN(n980), .Q(n882), 
        .QN(n3181) );
  DFFR_X1 \DRAM_mem_reg[13][25]  ( .D(n1791), .CK(CLK), .RN(n980), .Q(n883), 
        .QN(n3182) );
  DFFR_X1 \DRAM_mem_reg[13][24]  ( .D(n1790), .CK(CLK), .RN(n980), .Q(n884), 
        .QN(n3183) );
  DFFR_X1 \DRAM_mem_reg[13][23]  ( .D(n1789), .CK(CLK), .RN(n980), .Q(n885), 
        .QN(n3184) );
  DFFR_X1 \DRAM_mem_reg[13][22]  ( .D(n1788), .CK(CLK), .RN(n980), .Q(n886), 
        .QN(n3185) );
  DFFR_X1 \DRAM_mem_reg[13][21]  ( .D(n1787), .CK(CLK), .RN(n980), .Q(n887), 
        .QN(n3186) );
  DFFR_X1 \DRAM_mem_reg[13][20]  ( .D(n1786), .CK(CLK), .RN(n980), .Q(n888), 
        .QN(n3187) );
  DFFR_X1 \DRAM_mem_reg[13][19]  ( .D(n1785), .CK(CLK), .RN(n980), .Q(n889), 
        .QN(n3188) );
  DFFR_X1 \DRAM_mem_reg[13][18]  ( .D(n1784), .CK(CLK), .RN(n980), .Q(n890), 
        .QN(n3189) );
  DFFR_X1 \DRAM_mem_reg[13][17]  ( .D(n1783), .CK(CLK), .RN(n980), .Q(n891), 
        .QN(n3190) );
  DFFR_X1 \DRAM_mem_reg[13][16]  ( .D(n1782), .CK(CLK), .RN(n980), .Q(n892), 
        .QN(n3191) );
  DFFR_X1 \DRAM_mem_reg[13][15]  ( .D(n1781), .CK(CLK), .RN(n981), .Q(n762), 
        .QN(n3192) );
  DFFR_X1 \DRAM_mem_reg[13][14]  ( .D(n1780), .CK(CLK), .RN(n981), .Q(n259) );
  DFFR_X1 \DRAM_mem_reg[13][13]  ( .D(n1779), .CK(CLK), .RN(n981), .Q(n267) );
  DFFR_X1 \DRAM_mem_reg[13][12]  ( .D(n1778), .CK(CLK), .RN(n981), .Q(n275) );
  DFFR_X1 \DRAM_mem_reg[13][11]  ( .D(n1777), .CK(CLK), .RN(n981), .Q(n283) );
  DFFR_X1 \DRAM_mem_reg[13][10]  ( .D(n1776), .CK(CLK), .RN(n981), .Q(n291) );
  DFFR_X1 \DRAM_mem_reg[13][9]  ( .D(n1775), .CK(CLK), .RN(n981), .Q(n299) );
  DFFR_X1 \DRAM_mem_reg[13][8]  ( .D(n1774), .CK(CLK), .RN(n981), .Q(n307) );
  DFFR_X1 \DRAM_mem_reg[13][7]  ( .D(n1773), .CK(CLK), .RN(n981), .Q(n763), 
        .QN(n3193) );
  DFFR_X1 \DRAM_mem_reg[13][6]  ( .D(n1772), .CK(CLK), .RN(n981), .Q(n764), 
        .QN(n3194) );
  DFFR_X1 \DRAM_mem_reg[13][5]  ( .D(n1771), .CK(CLK), .RN(n981), .Q(n765), 
        .QN(n3195) );
  DFFR_X1 \DRAM_mem_reg[13][4]  ( .D(n1770), .CK(CLK), .RN(n981), .Q(n766), 
        .QN(n3196) );
  DFFR_X1 \DRAM_mem_reg[13][3]  ( .D(n1769), .CK(CLK), .RN(n982), .Q(n767), 
        .QN(n3197) );
  DFFR_X1 \DRAM_mem_reg[13][2]  ( .D(n1768), .CK(CLK), .RN(n982), .Q(n768), 
        .QN(n3198) );
  DFFR_X1 \DRAM_mem_reg[13][1]  ( .D(n1767), .CK(CLK), .RN(n982), .Q(n769), 
        .QN(n3199) );
  DFFR_X1 \DRAM_mem_reg[13][0]  ( .D(n1766), .CK(CLK), .RN(n982), .Q(n770), 
        .QN(n3200) );
  DFFR_X1 \DRAM_mem_reg[14][31]  ( .D(n1765), .CK(CLK), .RN(n982), .Q(n893), 
        .QN(n3201) );
  DFFR_X1 \DRAM_mem_reg[14][30]  ( .D(n1764), .CK(CLK), .RN(n982), .Q(n894), 
        .QN(n3202) );
  DFFR_X1 \DRAM_mem_reg[14][29]  ( .D(n1763), .CK(CLK), .RN(n982), .Q(n895), 
        .QN(n3203) );
  DFFR_X1 \DRAM_mem_reg[14][28]  ( .D(n1762), .CK(CLK), .RN(n982), .Q(n896), 
        .QN(n3204) );
  DFFR_X1 \DRAM_mem_reg[14][27]  ( .D(n1761), .CK(CLK), .RN(n982), .Q(n897), 
        .QN(n3205) );
  DFFR_X1 \DRAM_mem_reg[14][26]  ( .D(n1760), .CK(CLK), .RN(n982), .Q(n898), 
        .QN(n3206) );
  DFFR_X1 \DRAM_mem_reg[14][25]  ( .D(n1759), .CK(CLK), .RN(n982), .Q(n899), 
        .QN(n3207) );
  DFFR_X1 \DRAM_mem_reg[14][24]  ( .D(n1758), .CK(CLK), .RN(n982), .Q(n900), 
        .QN(n3208) );
  DFFR_X1 \DRAM_mem_reg[14][23]  ( .D(n1757), .CK(CLK), .RN(n983), .Q(n901), 
        .QN(n3209) );
  DFFR_X1 \DRAM_mem_reg[14][22]  ( .D(n1756), .CK(CLK), .RN(n983), .Q(n902), 
        .QN(n3210) );
  DFFR_X1 \DRAM_mem_reg[14][21]  ( .D(n1755), .CK(CLK), .RN(n983), .Q(n903), 
        .QN(n3211) );
  DFFR_X1 \DRAM_mem_reg[14][20]  ( .D(n1754), .CK(CLK), .RN(n983), .Q(n904), 
        .QN(n3212) );
  DFFR_X1 \DRAM_mem_reg[14][19]  ( .D(n1753), .CK(CLK), .RN(n983), .Q(n905), 
        .QN(n3213) );
  DFFR_X1 \DRAM_mem_reg[14][18]  ( .D(n1752), .CK(CLK), .RN(n983), .Q(n906), 
        .QN(n3214) );
  DFFR_X1 \DRAM_mem_reg[14][17]  ( .D(n1751), .CK(CLK), .RN(n983), .Q(n907), 
        .QN(n3215) );
  DFFR_X1 \DRAM_mem_reg[14][16]  ( .D(n1750), .CK(CLK), .RN(n983), .Q(n908), 
        .QN(n3216) );
  DFFR_X1 \DRAM_mem_reg[14][15]  ( .D(n1749), .CK(CLK), .RN(n983), .Q(n771), 
        .QN(n3217) );
  DFFR_X1 \DRAM_mem_reg[14][14]  ( .D(n1748), .CK(CLK), .RN(n983), .Q(n480), 
        .QN(n3218) );
  DFFR_X1 \DRAM_mem_reg[14][13]  ( .D(n1747), .CK(CLK), .RN(n983), .Q(n481), 
        .QN(n3219) );
  DFFR_X1 \DRAM_mem_reg[14][12]  ( .D(n1746), .CK(CLK), .RN(n983), .Q(n482), 
        .QN(n3220) );
  DFFR_X1 \DRAM_mem_reg[14][11]  ( .D(n1745), .CK(CLK), .RN(n984), .Q(n483), 
        .QN(n3221) );
  DFFR_X1 \DRAM_mem_reg[14][10]  ( .D(n1744), .CK(CLK), .RN(n984), .Q(n484), 
        .QN(n3222) );
  DFFR_X1 \DRAM_mem_reg[14][9]  ( .D(n1743), .CK(CLK), .RN(n984), .Q(n485), 
        .QN(n3223) );
  DFFR_X1 \DRAM_mem_reg[14][8]  ( .D(n1742), .CK(CLK), .RN(n984), .Q(n486), 
        .QN(n3224) );
  DFFR_X1 \DRAM_mem_reg[14][7]  ( .D(n1741), .CK(CLK), .RN(n984), .Q(n366) );
  DFFR_X1 \DRAM_mem_reg[14][6]  ( .D(n1740), .CK(CLK), .RN(n984), .Q(n370) );
  DFFR_X1 \DRAM_mem_reg[14][5]  ( .D(n1739), .CK(CLK), .RN(n984), .Q(n374) );
  DFFR_X1 \DRAM_mem_reg[14][4]  ( .D(n1738), .CK(CLK), .RN(n984), .Q(n378) );
  DFFR_X1 \DRAM_mem_reg[14][3]  ( .D(n1737), .CK(CLK), .RN(n984), .Q(n382) );
  DFFR_X1 \DRAM_mem_reg[14][2]  ( .D(n1736), .CK(CLK), .RN(n984), .Q(n386) );
  DFFR_X1 \DRAM_mem_reg[14][1]  ( .D(n1735), .CK(CLK), .RN(n984), .Q(n390) );
  DFFR_X1 \DRAM_mem_reg[14][0]  ( .D(n1734), .CK(CLK), .RN(n984), .Q(n394) );
  DFFR_X1 \DRAM_mem_reg[15][31]  ( .D(n1733), .CK(CLK), .RN(n985), .Q(n772), 
        .QN(n3225) );
  DFFR_X1 \DRAM_mem_reg[15][30]  ( .D(n1732), .CK(CLK), .RN(n985), .Q(n773), 
        .QN(n3226) );
  DFFR_X1 \DRAM_mem_reg[15][29]  ( .D(n1731), .CK(CLK), .RN(n985), .Q(n774), 
        .QN(n3227) );
  DFFR_X1 \DRAM_mem_reg[15][28]  ( .D(n1730), .CK(CLK), .RN(n985), .Q(n775), 
        .QN(n3228) );
  DFFR_X1 \DRAM_mem_reg[15][27]  ( .D(n1729), .CK(CLK), .RN(n985), .Q(n776), 
        .QN(n3229) );
  DFFR_X1 \DRAM_mem_reg[15][26]  ( .D(n1728), .CK(CLK), .RN(n985), .Q(n777), 
        .QN(n3230) );
  DFFR_X1 \DRAM_mem_reg[15][25]  ( .D(n1727), .CK(CLK), .RN(n985), .Q(n778), 
        .QN(n3231) );
  DFFR_X1 \DRAM_mem_reg[15][24]  ( .D(n1726), .CK(CLK), .RN(n985), .Q(n779), 
        .QN(n3232) );
  DFFR_X1 \DRAM_mem_reg[15][23]  ( .D(n1725), .CK(CLK), .RN(n985), .Q(n780), 
        .QN(n3233) );
  DFFR_X1 \DRAM_mem_reg[15][22]  ( .D(n1724), .CK(CLK), .RN(n985), .Q(n781), 
        .QN(n3234) );
  DFFR_X1 \DRAM_mem_reg[15][21]  ( .D(n1723), .CK(CLK), .RN(n985), .Q(n782), 
        .QN(n3235) );
  DFFR_X1 \DRAM_mem_reg[15][20]  ( .D(n1722), .CK(CLK), .RN(n985), .Q(n783), 
        .QN(n3236) );
  DFFR_X1 \DRAM_mem_reg[15][19]  ( .D(n1721), .CK(CLK), .RN(n986), .Q(n784), 
        .QN(n3237) );
  DFFR_X1 \DRAM_mem_reg[15][18]  ( .D(n1720), .CK(CLK), .RN(n986), .Q(n785), 
        .QN(n3238) );
  DFFR_X1 \DRAM_mem_reg[15][17]  ( .D(n1719), .CK(CLK), .RN(n986), .Q(n786), 
        .QN(n3239) );
  DFFR_X1 \DRAM_mem_reg[15][16]  ( .D(n1718), .CK(CLK), .RN(n986), .Q(n787), 
        .QN(n3240) );
  DFFR_X1 \DRAM_mem_reg[15][15]  ( .D(n1717), .CK(CLK), .RN(n986), .Q(n788), 
        .QN(n3241) );
  DFFR_X1 \DRAM_mem_reg[15][14]  ( .D(n1716), .CK(CLK), .RN(n986), .Q(n604), 
        .QN(n3242) );
  DFFR_X1 \DRAM_mem_reg[15][13]  ( .D(n1715), .CK(CLK), .RN(n986), .Q(n605), 
        .QN(n3243) );
  DFFR_X1 \DRAM_mem_reg[15][12]  ( .D(n1714), .CK(CLK), .RN(n986), .Q(n606), 
        .QN(n3244) );
  DFFR_X1 \DRAM_mem_reg[15][11]  ( .D(n1713), .CK(CLK), .RN(n986), .Q(n607), 
        .QN(n3245) );
  DFFR_X1 \DRAM_mem_reg[15][10]  ( .D(n1712), .CK(CLK), .RN(n986), .Q(n608), 
        .QN(n3246) );
  DFFR_X1 \DRAM_mem_reg[15][9]  ( .D(n1711), .CK(CLK), .RN(n986), .Q(n609), 
        .QN(n3247) );
  DFFR_X1 \DRAM_mem_reg[15][8]  ( .D(n1710), .CK(CLK), .RN(n986), .Q(n610), 
        .QN(n3248) );
  DFFR_X1 \DRAM_mem_reg[15][7]  ( .D(n1709), .CK(CLK), .RN(n987), .Q(n130) );
  DFFR_X1 \DRAM_mem_reg[15][6]  ( .D(n1708), .CK(CLK), .RN(n987), .Q(n134) );
  DFFR_X1 \DRAM_mem_reg[15][5]  ( .D(n1707), .CK(CLK), .RN(n987), .Q(n138) );
  DFFR_X1 \DRAM_mem_reg[15][4]  ( .D(n1706), .CK(CLK), .RN(n987), .Q(n142) );
  DFFR_X1 \DRAM_mem_reg[15][3]  ( .D(n1705), .CK(CLK), .RN(n987), .Q(n146) );
  DFFR_X1 \DRAM_mem_reg[15][2]  ( .D(n1704), .CK(CLK), .RN(n987), .Q(n150) );
  DFFR_X1 \DRAM_mem_reg[15][1]  ( .D(n1703), .CK(CLK), .RN(n987), .Q(n154) );
  DFFR_X1 \DRAM_mem_reg[15][0]  ( .D(n1702), .CK(CLK), .RN(n987), .Q(n158) );
  DFFR_X1 \DRAM_mem_reg[16][31]  ( .D(n1701), .CK(CLK), .RN(n987), .Q(n611), 
        .QN(n3249) );
  DFFR_X1 \DRAM_mem_reg[16][30]  ( .D(n1700), .CK(CLK), .RN(n987), .Q(n612), 
        .QN(n3250) );
  DFFR_X1 \DRAM_mem_reg[16][29]  ( .D(n1699), .CK(CLK), .RN(n987), .Q(n613), 
        .QN(n3251) );
  DFFR_X1 \DRAM_mem_reg[16][28]  ( .D(n1698), .CK(CLK), .RN(n987), .Q(n614), 
        .QN(n3252) );
  DFFR_X1 \DRAM_mem_reg[16][27]  ( .D(n1697), .CK(CLK), .RN(n988), .Q(n615), 
        .QN(n3253) );
  DFFR_X1 \DRAM_mem_reg[16][26]  ( .D(n1696), .CK(CLK), .RN(n988), .Q(n616), 
        .QN(n3254) );
  DFFR_X1 \DRAM_mem_reg[16][25]  ( .D(n1695), .CK(CLK), .RN(n988), .Q(n617), 
        .QN(n3255) );
  DFFR_X1 \DRAM_mem_reg[16][24]  ( .D(n1694), .CK(CLK), .RN(n988), .Q(n618), 
        .QN(n3256) );
  DFFR_X1 \DRAM_mem_reg[16][23]  ( .D(n1693), .CK(CLK), .RN(n988), .Q(n619), 
        .QN(n3257) );
  DFFR_X1 \DRAM_mem_reg[16][22]  ( .D(n1692), .CK(CLK), .RN(n988), .Q(n620), 
        .QN(n3258) );
  DFFR_X1 \DRAM_mem_reg[16][21]  ( .D(n1691), .CK(CLK), .RN(n988), .Q(n621), 
        .QN(n3259) );
  DFFR_X1 \DRAM_mem_reg[16][20]  ( .D(n1690), .CK(CLK), .RN(n988), .Q(n622), 
        .QN(n3260) );
  DFFR_X1 \DRAM_mem_reg[16][19]  ( .D(n1689), .CK(CLK), .RN(n988), .Q(n623), 
        .QN(n3261) );
  DFFR_X1 \DRAM_mem_reg[16][18]  ( .D(n1688), .CK(CLK), .RN(n988), .Q(n624), 
        .QN(n3262) );
  DFFR_X1 \DRAM_mem_reg[16][17]  ( .D(n1687), .CK(CLK), .RN(n988), .Q(n625), 
        .QN(n3263) );
  DFFR_X1 \DRAM_mem_reg[16][16]  ( .D(n1686), .CK(CLK), .RN(n988), .Q(n626), 
        .QN(n3264) );
  DFFR_X1 \DRAM_mem_reg[16][15]  ( .D(n1685), .CK(CLK), .RN(n989), .Q(n125) );
  DFFR_X1 \DRAM_mem_reg[16][14]  ( .D(n1684), .CK(CLK), .RN(n989), .Q(n2936), 
        .QN(n429) );
  DFFR_X1 \DRAM_mem_reg[16][13]  ( .D(n1683), .CK(CLK), .RN(n989), .Q(n2942), 
        .QN(n433) );
  DFFR_X1 \DRAM_mem_reg[16][12]  ( .D(n1682), .CK(CLK), .RN(n989), .Q(n2948), 
        .QN(n437) );
  DFFR_X1 \DRAM_mem_reg[16][11]  ( .D(n1681), .CK(CLK), .RN(n989), .Q(n2954), 
        .QN(n441) );
  DFFR_X1 \DRAM_mem_reg[16][10]  ( .D(n1680), .CK(CLK), .RN(n989), .Q(n2960), 
        .QN(n445) );
  DFFR_X1 \DRAM_mem_reg[16][9]  ( .D(n1679), .CK(CLK), .RN(n989), .Q(n2966), 
        .QN(n449) );
  DFFR_X1 \DRAM_mem_reg[16][8]  ( .D(n1678), .CK(CLK), .RN(n989), .Q(n2972), 
        .QN(n453) );
  DFFR_X1 \DRAM_mem_reg[16][7]  ( .D(n1677), .CK(CLK), .RN(n989), .Q(n909), 
        .QN(n3265) );
  DFFR_X1 \DRAM_mem_reg[16][6]  ( .D(n1676), .CK(CLK), .RN(n989), .Q(n910), 
        .QN(n3266) );
  DFFR_X1 \DRAM_mem_reg[16][5]  ( .D(n1675), .CK(CLK), .RN(n989), .Q(n911), 
        .QN(n3267) );
  DFFR_X1 \DRAM_mem_reg[16][4]  ( .D(n1674), .CK(CLK), .RN(n989), .Q(n912), 
        .QN(n3268) );
  DFFR_X1 \DRAM_mem_reg[16][3]  ( .D(n1673), .CK(CLK), .RN(n990), .Q(n913), 
        .QN(n3269) );
  DFFR_X1 \DRAM_mem_reg[16][2]  ( .D(n1672), .CK(CLK), .RN(n990), .Q(n914), 
        .QN(n3270) );
  DFFR_X1 \DRAM_mem_reg[16][1]  ( .D(n1671), .CK(CLK), .RN(n990), .Q(n915), 
        .QN(n3271) );
  DFFR_X1 \DRAM_mem_reg[16][0]  ( .D(n1670), .CK(CLK), .RN(n990), .Q(n916), 
        .QN(n3272) );
  DFFR_X1 \DRAM_mem_reg[17][31]  ( .D(n1669), .CK(CLK), .RN(n990), .Q(n341) );
  DFFR_X1 \DRAM_mem_reg[17][30]  ( .D(n1668), .CK(CLK), .RN(n990), .Q(n342) );
  DFFR_X1 \DRAM_mem_reg[17][29]  ( .D(n1667), .CK(CLK), .RN(n990), .Q(n343) );
  DFFR_X1 \DRAM_mem_reg[17][28]  ( .D(n1666), .CK(CLK), .RN(n990), .Q(n344) );
  DFFR_X1 \DRAM_mem_reg[17][27]  ( .D(n1665), .CK(CLK), .RN(n990), .Q(n345) );
  DFFR_X1 \DRAM_mem_reg[17][26]  ( .D(n1664), .CK(CLK), .RN(n990), .Q(n346) );
  DFFR_X1 \DRAM_mem_reg[17][25]  ( .D(n1663), .CK(CLK), .RN(n990), .Q(n347) );
  DFFR_X1 \DRAM_mem_reg[17][24]  ( .D(n1662), .CK(CLK), .RN(n990), .Q(n348) );
  DFFR_X1 \DRAM_mem_reg[17][23]  ( .D(n1661), .CK(CLK), .RN(n991), .Q(n349) );
  DFFR_X1 \DRAM_mem_reg[17][22]  ( .D(n1660), .CK(CLK), .RN(n991), .Q(n350) );
  DFFR_X1 \DRAM_mem_reg[17][21]  ( .D(n1659), .CK(CLK), .RN(n991), .Q(n351) );
  DFFR_X1 \DRAM_mem_reg[17][20]  ( .D(n1658), .CK(CLK), .RN(n991), .Q(n352) );
  DFFR_X1 \DRAM_mem_reg[17][19]  ( .D(n1657), .CK(CLK), .RN(n991), .Q(n353) );
  DFFR_X1 \DRAM_mem_reg[17][18]  ( .D(n1656), .CK(CLK), .RN(n991), .Q(n354) );
  DFFR_X1 \DRAM_mem_reg[17][17]  ( .D(n1655), .CK(CLK), .RN(n991), .Q(n355) );
  DFFR_X1 \DRAM_mem_reg[17][16]  ( .D(n1654), .CK(CLK), .RN(n991), .Q(n356) );
  DFFR_X1 \DRAM_mem_reg[17][15]  ( .D(n1653), .CK(CLK), .RN(n991), .Q(n123) );
  DFFR_X1 \DRAM_mem_reg[17][14]  ( .D(n1652), .CK(CLK), .RN(n991), .Q(n2935), 
        .QN(n177) );
  DFFR_X1 \DRAM_mem_reg[17][13]  ( .D(n1651), .CK(CLK), .RN(n991), .Q(n2941), 
        .QN(n181) );
  DFFR_X1 \DRAM_mem_reg[17][12]  ( .D(n1650), .CK(CLK), .RN(n991), .Q(n2947), 
        .QN(n185) );
  DFFR_X1 \DRAM_mem_reg[17][11]  ( .D(n1649), .CK(CLK), .RN(n992), .Q(n2953), 
        .QN(n189) );
  DFFR_X1 \DRAM_mem_reg[17][10]  ( .D(n1648), .CK(CLK), .RN(n992), .Q(n2959), 
        .QN(n193) );
  DFFR_X1 \DRAM_mem_reg[17][9]  ( .D(n1647), .CK(CLK), .RN(n992), .Q(n2965), 
        .QN(n197) );
  DFFR_X1 \DRAM_mem_reg[17][8]  ( .D(n1646), .CK(CLK), .RN(n992), .Q(n2971), 
        .QN(n201) );
  DFFR_X1 \DRAM_mem_reg[17][7]  ( .D(n1645), .CK(CLK), .RN(n992), .Q(n789), 
        .QN(n3273) );
  DFFR_X1 \DRAM_mem_reg[17][6]  ( .D(n1644), .CK(CLK), .RN(n992), .Q(n790), 
        .QN(n3274) );
  DFFR_X1 \DRAM_mem_reg[17][5]  ( .D(n1643), .CK(CLK), .RN(n992), .Q(n791), 
        .QN(n3275) );
  DFFR_X1 \DRAM_mem_reg[17][4]  ( .D(n1642), .CK(CLK), .RN(n992), .Q(n792), 
        .QN(n3276) );
  DFFR_X1 \DRAM_mem_reg[17][3]  ( .D(n1641), .CK(CLK), .RN(n992), .Q(n793), 
        .QN(n3277) );
  DFFR_X1 \DRAM_mem_reg[17][2]  ( .D(n1640), .CK(CLK), .RN(n992), .Q(n794), 
        .QN(n3278) );
  DFFR_X1 \DRAM_mem_reg[17][1]  ( .D(n1639), .CK(CLK), .RN(n992), .Q(n795), 
        .QN(n3279) );
  DFFR_X1 \DRAM_mem_reg[17][0]  ( .D(n1638), .CK(CLK), .RN(n992), .Q(n796), 
        .QN(n3280) );
  DFFR_X1 \DRAM_mem_reg[18][31]  ( .D(n1637), .CK(CLK), .RN(n993), .Q(n487), 
        .QN(n3281) );
  DFFR_X1 \DRAM_mem_reg[18][30]  ( .D(n1636), .CK(CLK), .RN(n993), .Q(n488), 
        .QN(n3282) );
  DFFR_X1 \DRAM_mem_reg[18][29]  ( .D(n1635), .CK(CLK), .RN(n993), .Q(n489), 
        .QN(n3283) );
  DFFR_X1 \DRAM_mem_reg[18][28]  ( .D(n1634), .CK(CLK), .RN(n993), .Q(n490), 
        .QN(n3284) );
  DFFR_X1 \DRAM_mem_reg[18][27]  ( .D(n1633), .CK(CLK), .RN(n993), .Q(n491), 
        .QN(n3285) );
  DFFR_X1 \DRAM_mem_reg[18][26]  ( .D(n1632), .CK(CLK), .RN(n993), .Q(n492), 
        .QN(n3286) );
  DFFR_X1 \DRAM_mem_reg[18][25]  ( .D(n1631), .CK(CLK), .RN(n993), .Q(n493), 
        .QN(n3287) );
  DFFR_X1 \DRAM_mem_reg[18][24]  ( .D(n1630), .CK(CLK), .RN(n993), .Q(n494), 
        .QN(n3288) );
  DFFR_X1 \DRAM_mem_reg[18][23]  ( .D(n1629), .CK(CLK), .RN(n993), .Q(n495), 
        .QN(n3289) );
  DFFR_X1 \DRAM_mem_reg[18][22]  ( .D(n1628), .CK(CLK), .RN(n993), .Q(n496), 
        .QN(n3290) );
  DFFR_X1 \DRAM_mem_reg[18][21]  ( .D(n1627), .CK(CLK), .RN(n993), .Q(n497), 
        .QN(n3291) );
  DFFR_X1 \DRAM_mem_reg[18][20]  ( .D(n1626), .CK(CLK), .RN(n993), .Q(n498), 
        .QN(n3292) );
  DFFR_X1 \DRAM_mem_reg[18][19]  ( .D(n1625), .CK(CLK), .RN(n994), .Q(n499), 
        .QN(n3293) );
  DFFR_X1 \DRAM_mem_reg[18][18]  ( .D(n1624), .CK(CLK), .RN(n994), .Q(n500), 
        .QN(n3294) );
  DFFR_X1 \DRAM_mem_reg[18][17]  ( .D(n1623), .CK(CLK), .RN(n994), .Q(n501), 
        .QN(n3295) );
  DFFR_X1 \DRAM_mem_reg[18][16]  ( .D(n1622), .CK(CLK), .RN(n994), .Q(n502), 
        .QN(n3296) );
  DFFR_X1 \DRAM_mem_reg[18][15]  ( .D(n1621), .CK(CLK), .RN(n994), .Q(n121) );
  DFFR_X1 \DRAM_mem_reg[18][14]  ( .D(n1620), .CK(CLK), .RN(n994), .Q(n17) );
  DFFR_X1 \DRAM_mem_reg[18][13]  ( .D(n1619), .CK(CLK), .RN(n994), .Q(n25) );
  DFFR_X1 \DRAM_mem_reg[18][12]  ( .D(n1618), .CK(CLK), .RN(n994), .Q(n33) );
  DFFR_X1 \DRAM_mem_reg[18][11]  ( .D(n1617), .CK(CLK), .RN(n994), .Q(n41) );
  DFFR_X1 \DRAM_mem_reg[18][10]  ( .D(n1616), .CK(CLK), .RN(n994), .Q(n49) );
  DFFR_X1 \DRAM_mem_reg[18][9]  ( .D(n1615), .CK(CLK), .RN(n994), .Q(n57) );
  DFFR_X1 \DRAM_mem_reg[18][8]  ( .D(n1614), .CK(CLK), .RN(n994), .Q(n65) );
  DFFR_X1 \DRAM_mem_reg[18][7]  ( .D(n1613), .CK(CLK), .RN(n995), .Q(n2980) );
  DFFR_X1 \DRAM_mem_reg[18][6]  ( .D(n1612), .CK(CLK), .RN(n995), .Q(n2988) );
  DFFR_X1 \DRAM_mem_reg[18][5]  ( .D(n1611), .CK(CLK), .RN(n995), .Q(n2996) );
  DFFR_X1 \DRAM_mem_reg[18][4]  ( .D(n1610), .CK(CLK), .RN(n995), .Q(n3004) );
  DFFR_X1 \DRAM_mem_reg[18][3]  ( .D(n1609), .CK(CLK), .RN(n995), .Q(n3012) );
  DFFR_X1 \DRAM_mem_reg[18][2]  ( .D(n1608), .CK(CLK), .RN(n995), .Q(n3020) );
  DFFR_X1 \DRAM_mem_reg[18][1]  ( .D(n1607), .CK(CLK), .RN(n995), .Q(n3028) );
  DFFR_X1 \DRAM_mem_reg[18][0]  ( .D(n1606), .CK(CLK), .RN(n995), .Q(n3036) );
  DFFR_X1 \DRAM_mem_reg[19][31]  ( .D(n1605), .CK(CLK), .RN(n995), .Q(n627), 
        .QN(n3297) );
  DFFR_X1 \DRAM_mem_reg[19][30]  ( .D(n1604), .CK(CLK), .RN(n995), .Q(n628), 
        .QN(n3298) );
  DFFR_X1 \DRAM_mem_reg[19][29]  ( .D(n1603), .CK(CLK), .RN(n995), .Q(n629), 
        .QN(n3299) );
  DFFR_X1 \DRAM_mem_reg[19][28]  ( .D(n1602), .CK(CLK), .RN(n995), .Q(n630), 
        .QN(n3300) );
  DFFR_X1 \DRAM_mem_reg[19][27]  ( .D(n1601), .CK(CLK), .RN(n996), .Q(n631), 
        .QN(n3301) );
  DFFR_X1 \DRAM_mem_reg[19][26]  ( .D(n1600), .CK(CLK), .RN(n996), .Q(n632), 
        .QN(n3302) );
  DFFR_X1 \DRAM_mem_reg[19][25]  ( .D(n1599), .CK(CLK), .RN(n996), .Q(n633), 
        .QN(n3303) );
  DFFR_X1 \DRAM_mem_reg[19][24]  ( .D(n1598), .CK(CLK), .RN(n996), .Q(n634), 
        .QN(n3304) );
  DFFR_X1 \DRAM_mem_reg[19][23]  ( .D(n1597), .CK(CLK), .RN(n996), .Q(n635), 
        .QN(n3305) );
  DFFR_X1 \DRAM_mem_reg[19][22]  ( .D(n1596), .CK(CLK), .RN(n996), .Q(n636), 
        .QN(n3306) );
  DFFR_X1 \DRAM_mem_reg[19][21]  ( .D(n1595), .CK(CLK), .RN(n996), .Q(n637), 
        .QN(n3307) );
  DFFR_X1 \DRAM_mem_reg[19][20]  ( .D(n1594), .CK(CLK), .RN(n996), .Q(n638), 
        .QN(n3308) );
  DFFR_X1 \DRAM_mem_reg[19][19]  ( .D(n1593), .CK(CLK), .RN(n996), .Q(n639), 
        .QN(n3309) );
  DFFR_X1 \DRAM_mem_reg[19][18]  ( .D(n1592), .CK(CLK), .RN(n996), .Q(n640), 
        .QN(n3310) );
  DFFR_X1 \DRAM_mem_reg[19][17]  ( .D(n1591), .CK(CLK), .RN(n996), .Q(n641), 
        .QN(n3311) );
  DFFR_X1 \DRAM_mem_reg[19][16]  ( .D(n1590), .CK(CLK), .RN(n996), .Q(n642), 
        .QN(n3312) );
  DFFR_X1 \DRAM_mem_reg[19][15]  ( .D(n1589), .CK(CLK), .RN(n997), .Q(n127) );
  DFFR_X1 \DRAM_mem_reg[19][14]  ( .D(n1588), .CK(CLK), .RN(n997), .Q(n253) );
  DFFR_X1 \DRAM_mem_reg[19][13]  ( .D(n1587), .CK(CLK), .RN(n997), .Q(n261) );
  DFFR_X1 \DRAM_mem_reg[19][12]  ( .D(n1586), .CK(CLK), .RN(n997), .Q(n269) );
  DFFR_X1 \DRAM_mem_reg[19][11]  ( .D(n1585), .CK(CLK), .RN(n997), .Q(n277) );
  DFFR_X1 \DRAM_mem_reg[19][10]  ( .D(n1584), .CK(CLK), .RN(n997), .Q(n285) );
  DFFR_X1 \DRAM_mem_reg[19][9]  ( .D(n1583), .CK(CLK), .RN(n997), .Q(n293) );
  DFFR_X1 \DRAM_mem_reg[19][8]  ( .D(n1582), .CK(CLK), .RN(n997), .Q(n301) );
  DFFR_X1 \DRAM_mem_reg[19][7]  ( .D(n1581), .CK(CLK), .RN(n997), .Q(n2979) );
  DFFR_X1 \DRAM_mem_reg[19][6]  ( .D(n1580), .CK(CLK), .RN(n997), .Q(n2987) );
  DFFR_X1 \DRAM_mem_reg[19][5]  ( .D(n1579), .CK(CLK), .RN(n997), .Q(n2995) );
  DFFR_X1 \DRAM_mem_reg[19][4]  ( .D(n1578), .CK(CLK), .RN(n997), .Q(n3003) );
  DFFR_X1 \DRAM_mem_reg[19][3]  ( .D(n1577), .CK(CLK), .RN(n998), .Q(n3011) );
  DFFR_X1 \DRAM_mem_reg[19][2]  ( .D(n1576), .CK(CLK), .RN(n998), .Q(n3019) );
  DFFR_X1 \DRAM_mem_reg[19][1]  ( .D(n1575), .CK(CLK), .RN(n998), .Q(n3027) );
  DFFR_X1 \DRAM_mem_reg[19][0]  ( .D(n1574), .CK(CLK), .RN(n998), .Q(n3035) );
  DFFR_X1 \DRAM_mem_reg[20][31]  ( .D(n1573), .CK(CLK), .RN(n998), .Q(n643), 
        .QN(n3313) );
  DFFR_X1 \DRAM_mem_reg[20][30]  ( .D(n1572), .CK(CLK), .RN(n998), .Q(n644), 
        .QN(n3314) );
  DFFR_X1 \DRAM_mem_reg[20][29]  ( .D(n1571), .CK(CLK), .RN(n998), .Q(n645), 
        .QN(n3315) );
  DFFR_X1 \DRAM_mem_reg[20][28]  ( .D(n1570), .CK(CLK), .RN(n998), .Q(n646), 
        .QN(n3316) );
  DFFR_X1 \DRAM_mem_reg[20][27]  ( .D(n1569), .CK(CLK), .RN(n998), .Q(n647), 
        .QN(n3317) );
  DFFR_X1 \DRAM_mem_reg[20][26]  ( .D(n1568), .CK(CLK), .RN(n998), .Q(n648), 
        .QN(n3318) );
  DFFR_X1 \DRAM_mem_reg[20][25]  ( .D(n1567), .CK(CLK), .RN(n998), .Q(n649), 
        .QN(n3319) );
  DFFR_X1 \DRAM_mem_reg[20][24]  ( .D(n1566), .CK(CLK), .RN(n998), .Q(n650), 
        .QN(n3320) );
  DFFR_X1 \DRAM_mem_reg[20][23]  ( .D(n1565), .CK(CLK), .RN(n999), .Q(n651), 
        .QN(n3321) );
  DFFR_X1 \DRAM_mem_reg[20][22]  ( .D(n1564), .CK(CLK), .RN(n999), .Q(n652), 
        .QN(n3322) );
  DFFR_X1 \DRAM_mem_reg[20][21]  ( .D(n1563), .CK(CLK), .RN(n999), .Q(n653), 
        .QN(n3323) );
  DFFR_X1 \DRAM_mem_reg[20][20]  ( .D(n1562), .CK(CLK), .RN(n999), .Q(n654), 
        .QN(n3324) );
  DFFR_X1 \DRAM_mem_reg[20][19]  ( .D(n1561), .CK(CLK), .RN(n999), .Q(n655), 
        .QN(n3325) );
  DFFR_X1 \DRAM_mem_reg[20][18]  ( .D(n1560), .CK(CLK), .RN(n999), .Q(n656), 
        .QN(n3326) );
  DFFR_X1 \DRAM_mem_reg[20][17]  ( .D(n1559), .CK(CLK), .RN(n999), .Q(n657), 
        .QN(n3327) );
  DFFR_X1 \DRAM_mem_reg[20][16]  ( .D(n1558), .CK(CLK), .RN(n999), .Q(n658), 
        .QN(n3328) );
  DFFR_X1 \DRAM_mem_reg[20][15]  ( .D(n1557), .CK(CLK), .RN(n999), .Q(n361) );
  DFFR_X1 \DRAM_mem_reg[20][14]  ( .D(n1556), .CK(CLK), .RN(n999), .Q(n2934), 
        .QN(n430) );
  DFFR_X1 \DRAM_mem_reg[20][13]  ( .D(n1555), .CK(CLK), .RN(n999), .Q(n2940), 
        .QN(n434) );
  DFFR_X1 \DRAM_mem_reg[20][12]  ( .D(n1554), .CK(CLK), .RN(n999), .Q(n2946), 
        .QN(n438) );
  DFFR_X1 \DRAM_mem_reg[20][11]  ( .D(n1553), .CK(CLK), .RN(n1000), .Q(n2952), 
        .QN(n442) );
  DFFR_X1 \DRAM_mem_reg[20][10]  ( .D(n1552), .CK(CLK), .RN(n1000), .Q(n2958), 
        .QN(n446) );
  DFFR_X1 \DRAM_mem_reg[20][9]  ( .D(n1551), .CK(CLK), .RN(n1000), .Q(n2964), 
        .QN(n450) );
  DFFR_X1 \DRAM_mem_reg[20][8]  ( .D(n1550), .CK(CLK), .RN(n1000), .Q(n2970), 
        .QN(n454) );
  DFFR_X1 \DRAM_mem_reg[20][7]  ( .D(n1549), .CK(CLK), .RN(n1000), .Q(n917), 
        .QN(n3329) );
  DFFR_X1 \DRAM_mem_reg[20][6]  ( .D(n1548), .CK(CLK), .RN(n1000), .Q(n918), 
        .QN(n3330) );
  DFFR_X1 \DRAM_mem_reg[20][5]  ( .D(n1547), .CK(CLK), .RN(n1000), .Q(n919), 
        .QN(n3331) );
  DFFR_X1 \DRAM_mem_reg[20][4]  ( .D(n1546), .CK(CLK), .RN(n1000), .Q(n920), 
        .QN(n3332) );
  DFFR_X1 \DRAM_mem_reg[20][3]  ( .D(n1545), .CK(CLK), .RN(n1000), .Q(n921), 
        .QN(n3333) );
  DFFR_X1 \DRAM_mem_reg[20][2]  ( .D(n1544), .CK(CLK), .RN(n1000), .Q(n922), 
        .QN(n3334) );
  DFFR_X1 \DRAM_mem_reg[20][1]  ( .D(n1543), .CK(CLK), .RN(n1000), .Q(n923), 
        .QN(n3335) );
  DFFR_X1 \DRAM_mem_reg[20][0]  ( .D(n1542), .CK(CLK), .RN(n1000), .Q(n924), 
        .QN(n3336) );
  DFFR_X1 \DRAM_mem_reg[21][31]  ( .D(n1541), .CK(CLK), .RN(n1001), .Q(n503), 
        .QN(n3337) );
  DFFR_X1 \DRAM_mem_reg[21][30]  ( .D(n1540), .CK(CLK), .RN(n1001), .Q(n504), 
        .QN(n3338) );
  DFFR_X1 \DRAM_mem_reg[21][29]  ( .D(n1539), .CK(CLK), .RN(n1001), .Q(n505), 
        .QN(n3339) );
  DFFR_X1 \DRAM_mem_reg[21][28]  ( .D(n1538), .CK(CLK), .RN(n1001), .Q(n506), 
        .QN(n3340) );
  DFFR_X1 \DRAM_mem_reg[21][27]  ( .D(n1537), .CK(CLK), .RN(n1001), .Q(n507), 
        .QN(n3341) );
  DFFR_X1 \DRAM_mem_reg[21][26]  ( .D(n1536), .CK(CLK), .RN(n1001), .Q(n508), 
        .QN(n3342) );
  DFFR_X1 \DRAM_mem_reg[21][25]  ( .D(n1535), .CK(CLK), .RN(n1001), .Q(n509), 
        .QN(n3343) );
  DFFR_X1 \DRAM_mem_reg[21][24]  ( .D(n1534), .CK(CLK), .RN(n1001), .Q(n510), 
        .QN(n3344) );
  DFFR_X1 \DRAM_mem_reg[21][23]  ( .D(n1533), .CK(CLK), .RN(n1001), .Q(n511), 
        .QN(n3345) );
  DFFR_X1 \DRAM_mem_reg[21][22]  ( .D(n1532), .CK(CLK), .RN(n1001), .Q(n512), 
        .QN(n3346) );
  DFFR_X1 \DRAM_mem_reg[21][21]  ( .D(n1531), .CK(CLK), .RN(n1001), .Q(n513), 
        .QN(n3347) );
  DFFR_X1 \DRAM_mem_reg[21][20]  ( .D(n1530), .CK(CLK), .RN(n1001), .Q(n514), 
        .QN(n3348) );
  DFFR_X1 \DRAM_mem_reg[21][19]  ( .D(n1529), .CK(CLK), .RN(n1002), .Q(n515), 
        .QN(n3349) );
  DFFR_X1 \DRAM_mem_reg[21][18]  ( .D(n1528), .CK(CLK), .RN(n1002), .Q(n516), 
        .QN(n3350) );
  DFFR_X1 \DRAM_mem_reg[21][17]  ( .D(n1527), .CK(CLK), .RN(n1002), .Q(n517), 
        .QN(n3351) );
  DFFR_X1 \DRAM_mem_reg[21][16]  ( .D(n1526), .CK(CLK), .RN(n1002), .Q(n518), 
        .QN(n3352) );
  DFFR_X1 \DRAM_mem_reg[21][15]  ( .D(n1525), .CK(CLK), .RN(n1002), .Q(n359)
         );
  DFFR_X1 \DRAM_mem_reg[21][14]  ( .D(n1524), .CK(CLK), .RN(n1002), .Q(n2933), 
        .QN(n178) );
  DFFR_X1 \DRAM_mem_reg[21][13]  ( .D(n1523), .CK(CLK), .RN(n1002), .Q(n2939), 
        .QN(n182) );
  DFFR_X1 \DRAM_mem_reg[21][12]  ( .D(n1522), .CK(CLK), .RN(n1002), .Q(n2945), 
        .QN(n186) );
  DFFR_X1 \DRAM_mem_reg[21][11]  ( .D(n1521), .CK(CLK), .RN(n1002), .Q(n2951), 
        .QN(n190) );
  DFFR_X1 \DRAM_mem_reg[21][10]  ( .D(n1520), .CK(CLK), .RN(n1002), .Q(n2957), 
        .QN(n194) );
  DFFR_X1 \DRAM_mem_reg[21][9]  ( .D(n1519), .CK(CLK), .RN(n1002), .Q(n2963), 
        .QN(n198) );
  DFFR_X1 \DRAM_mem_reg[21][8]  ( .D(n1518), .CK(CLK), .RN(n1002), .Q(n2969), 
        .QN(n202) );
  DFFR_X1 \DRAM_mem_reg[21][7]  ( .D(n1517), .CK(CLK), .RN(n1003), .Q(n797), 
        .QN(n3353) );
  DFFR_X1 \DRAM_mem_reg[21][6]  ( .D(n1516), .CK(CLK), .RN(n1003), .Q(n798), 
        .QN(n3354) );
  DFFR_X1 \DRAM_mem_reg[21][5]  ( .D(n1515), .CK(CLK), .RN(n1003), .Q(n799), 
        .QN(n3355) );
  DFFR_X1 \DRAM_mem_reg[21][4]  ( .D(n1514), .CK(CLK), .RN(n1003), .Q(n800), 
        .QN(n3356) );
  DFFR_X1 \DRAM_mem_reg[21][3]  ( .D(n1513), .CK(CLK), .RN(n1003), .Q(n801), 
        .QN(n3357) );
  DFFR_X1 \DRAM_mem_reg[21][2]  ( .D(n1512), .CK(CLK), .RN(n1003), .Q(n802), 
        .QN(n3358) );
  DFFR_X1 \DRAM_mem_reg[21][1]  ( .D(n1511), .CK(CLK), .RN(n1003), .Q(n803), 
        .QN(n3359) );
  DFFR_X1 \DRAM_mem_reg[21][0]  ( .D(n1510), .CK(CLK), .RN(n1003), .Q(n804), 
        .QN(n3360) );
  DFFR_X1 \DRAM_mem_reg[22][31]  ( .D(n1509), .CK(CLK), .RN(n1003), .Q(n519), 
        .QN(n3361) );
  DFFR_X1 \DRAM_mem_reg[22][30]  ( .D(n1508), .CK(CLK), .RN(n1003), .Q(n520), 
        .QN(n3362) );
  DFFR_X1 \DRAM_mem_reg[22][29]  ( .D(n1507), .CK(CLK), .RN(n1003), .Q(n521), 
        .QN(n3363) );
  DFFR_X1 \DRAM_mem_reg[22][28]  ( .D(n1506), .CK(CLK), .RN(n1003), .Q(n522), 
        .QN(n3364) );
  DFFR_X1 \DRAM_mem_reg[22][27]  ( .D(n1505), .CK(CLK), .RN(n1004), .Q(n523), 
        .QN(n3365) );
  DFFR_X1 \DRAM_mem_reg[22][26]  ( .D(n1504), .CK(CLK), .RN(n1004), .Q(n524), 
        .QN(n3366) );
  DFFR_X1 \DRAM_mem_reg[22][25]  ( .D(n1503), .CK(CLK), .RN(n1004), .Q(n525), 
        .QN(n3367) );
  DFFR_X1 \DRAM_mem_reg[22][24]  ( .D(n1502), .CK(CLK), .RN(n1004), .Q(n526), 
        .QN(n3368) );
  DFFR_X1 \DRAM_mem_reg[22][23]  ( .D(n1501), .CK(CLK), .RN(n1004), .Q(n527), 
        .QN(n3369) );
  DFFR_X1 \DRAM_mem_reg[22][22]  ( .D(n1500), .CK(CLK), .RN(n1004), .Q(n528), 
        .QN(n3370) );
  DFFR_X1 \DRAM_mem_reg[22][21]  ( .D(n1499), .CK(CLK), .RN(n1004), .Q(n529), 
        .QN(n3371) );
  DFFR_X1 \DRAM_mem_reg[22][20]  ( .D(n1498), .CK(CLK), .RN(n1004), .Q(n530), 
        .QN(n3372) );
  DFFR_X1 \DRAM_mem_reg[22][19]  ( .D(n1497), .CK(CLK), .RN(n1004), .Q(n531), 
        .QN(n3373) );
  DFFR_X1 \DRAM_mem_reg[22][18]  ( .D(n1496), .CK(CLK), .RN(n1004), .Q(n532), 
        .QN(n3374) );
  DFFR_X1 \DRAM_mem_reg[22][17]  ( .D(n1495), .CK(CLK), .RN(n1004), .Q(n533), 
        .QN(n3375) );
  DFFR_X1 \DRAM_mem_reg[22][16]  ( .D(n1494), .CK(CLK), .RN(n1004), .Q(n534), 
        .QN(n3376) );
  DFFR_X1 \DRAM_mem_reg[22][15]  ( .D(n1493), .CK(CLK), .RN(n1005), .Q(n357)
         );
  DFFR_X1 \DRAM_mem_reg[22][14]  ( .D(n1492), .CK(CLK), .RN(n1005), .Q(n18) );
  DFFR_X1 \DRAM_mem_reg[22][13]  ( .D(n1491), .CK(CLK), .RN(n1005), .Q(n26) );
  DFFR_X1 \DRAM_mem_reg[22][12]  ( .D(n1490), .CK(CLK), .RN(n1005), .Q(n34) );
  DFFR_X1 \DRAM_mem_reg[22][11]  ( .D(n1489), .CK(CLK), .RN(n1005), .Q(n42) );
  DFFR_X1 \DRAM_mem_reg[22][10]  ( .D(n1488), .CK(CLK), .RN(n1005), .Q(n50) );
  DFFR_X1 \DRAM_mem_reg[22][9]  ( .D(n1487), .CK(CLK), .RN(n1005), .Q(n58) );
  DFFR_X1 \DRAM_mem_reg[22][8]  ( .D(n1486), .CK(CLK), .RN(n1005), .Q(n66) );
  DFFR_X1 \DRAM_mem_reg[22][7]  ( .D(n1485), .CK(CLK), .RN(n1005), .Q(n2982)
         );
  DFFR_X1 \DRAM_mem_reg[22][6]  ( .D(n1484), .CK(CLK), .RN(n1005), .Q(n2990)
         );
  DFFR_X1 \DRAM_mem_reg[22][5]  ( .D(n1483), .CK(CLK), .RN(n1005), .Q(n2998)
         );
  DFFR_X1 \DRAM_mem_reg[22][4]  ( .D(n1482), .CK(CLK), .RN(n1005), .Q(n3006)
         );
  DFFR_X1 \DRAM_mem_reg[22][3]  ( .D(n1481), .CK(CLK), .RN(n1006), .Q(n3014)
         );
  DFFR_X1 \DRAM_mem_reg[22][2]  ( .D(n1480), .CK(CLK), .RN(n1006), .Q(n3022)
         );
  DFFR_X1 \DRAM_mem_reg[22][1]  ( .D(n1479), .CK(CLK), .RN(n1006), .Q(n3030)
         );
  DFFR_X1 \DRAM_mem_reg[22][0]  ( .D(n1478), .CK(CLK), .RN(n1006), .Q(n3038)
         );
  DFFR_X1 \DRAM_mem_reg[23][31]  ( .D(n1477), .CK(CLK), .RN(n1006), .Q(n659), 
        .QN(n3377) );
  DFFR_X1 \DRAM_mem_reg[23][30]  ( .D(n1476), .CK(CLK), .RN(n1006), .Q(n660), 
        .QN(n3378) );
  DFFR_X1 \DRAM_mem_reg[23][29]  ( .D(n1475), .CK(CLK), .RN(n1006), .Q(n661), 
        .QN(n3379) );
  DFFR_X1 \DRAM_mem_reg[23][28]  ( .D(n1474), .CK(CLK), .RN(n1006), .Q(n662), 
        .QN(n3380) );
  DFFR_X1 \DRAM_mem_reg[23][27]  ( .D(n1473), .CK(CLK), .RN(n1006), .Q(n663), 
        .QN(n3381) );
  DFFR_X1 \DRAM_mem_reg[23][26]  ( .D(n1472), .CK(CLK), .RN(n1006), .Q(n664), 
        .QN(n3382) );
  DFFR_X1 \DRAM_mem_reg[23][25]  ( .D(n1471), .CK(CLK), .RN(n1006), .Q(n665), 
        .QN(n3383) );
  DFFR_X1 \DRAM_mem_reg[23][24]  ( .D(n1470), .CK(CLK), .RN(n1006), .Q(n666), 
        .QN(n3384) );
  DFFR_X1 \DRAM_mem_reg[23][23]  ( .D(n1469), .CK(CLK), .RN(n1007), .Q(n667), 
        .QN(n3385) );
  DFFR_X1 \DRAM_mem_reg[23][22]  ( .D(n1468), .CK(CLK), .RN(n1007), .Q(n668), 
        .QN(n3386) );
  DFFR_X1 \DRAM_mem_reg[23][21]  ( .D(n1467), .CK(CLK), .RN(n1007), .Q(n669), 
        .QN(n3387) );
  DFFR_X1 \DRAM_mem_reg[23][20]  ( .D(n1466), .CK(CLK), .RN(n1007), .Q(n670), 
        .QN(n3388) );
  DFFR_X1 \DRAM_mem_reg[23][19]  ( .D(n1465), .CK(CLK), .RN(n1007), .Q(n671), 
        .QN(n3389) );
  DFFR_X1 \DRAM_mem_reg[23][18]  ( .D(n1464), .CK(CLK), .RN(n1007), .Q(n672), 
        .QN(n3390) );
  DFFR_X1 \DRAM_mem_reg[23][17]  ( .D(n1463), .CK(CLK), .RN(n1007), .Q(n673), 
        .QN(n3391) );
  DFFR_X1 \DRAM_mem_reg[23][16]  ( .D(n1462), .CK(CLK), .RN(n1007), .Q(n674), 
        .QN(n3392) );
  DFFR_X1 \DRAM_mem_reg[23][15]  ( .D(n1461), .CK(CLK), .RN(n1007), .Q(n363)
         );
  DFFR_X1 \DRAM_mem_reg[23][14]  ( .D(n1460), .CK(CLK), .RN(n1007), .Q(n254)
         );
  DFFR_X1 \DRAM_mem_reg[23][13]  ( .D(n1459), .CK(CLK), .RN(n1007), .Q(n262)
         );
  DFFR_X1 \DRAM_mem_reg[23][12]  ( .D(n1458), .CK(CLK), .RN(n1007), .Q(n270)
         );
  DFFR_X1 \DRAM_mem_reg[23][11]  ( .D(n1457), .CK(CLK), .RN(n1008), .Q(n278)
         );
  DFFR_X1 \DRAM_mem_reg[23][10]  ( .D(n1456), .CK(CLK), .RN(n1008), .Q(n286)
         );
  DFFR_X1 \DRAM_mem_reg[23][9]  ( .D(n1455), .CK(CLK), .RN(n1008), .Q(n294) );
  DFFR_X1 \DRAM_mem_reg[23][8]  ( .D(n1454), .CK(CLK), .RN(n1008), .Q(n302) );
  DFFR_X1 \DRAM_mem_reg[23][7]  ( .D(n1453), .CK(CLK), .RN(n1008), .Q(n2981)
         );
  DFFR_X1 \DRAM_mem_reg[23][6]  ( .D(n1452), .CK(CLK), .RN(n1008), .Q(n2989)
         );
  DFFR_X1 \DRAM_mem_reg[23][5]  ( .D(n1451), .CK(CLK), .RN(n1008), .Q(n2997)
         );
  DFFR_X1 \DRAM_mem_reg[23][4]  ( .D(n1450), .CK(CLK), .RN(n1008), .Q(n3005)
         );
  DFFR_X1 \DRAM_mem_reg[23][3]  ( .D(n1449), .CK(CLK), .RN(n1008), .Q(n3013)
         );
  DFFR_X1 \DRAM_mem_reg[23][2]  ( .D(n1448), .CK(CLK), .RN(n1008), .Q(n3021)
         );
  DFFR_X1 \DRAM_mem_reg[23][1]  ( .D(n1447), .CK(CLK), .RN(n1008), .Q(n3029)
         );
  DFFR_X1 \DRAM_mem_reg[23][0]  ( .D(n1446), .CK(CLK), .RN(n1008), .Q(n3037)
         );
  DFFR_X1 \DRAM_mem_reg[24][31]  ( .D(n1445), .CK(CLK), .RN(n1009), .Q(n675), 
        .QN(n3393) );
  DFFR_X1 \DRAM_mem_reg[24][30]  ( .D(n1444), .CK(CLK), .RN(n1009), .Q(n676), 
        .QN(n3394) );
  DFFR_X1 \DRAM_mem_reg[24][29]  ( .D(n1443), .CK(CLK), .RN(n1009), .Q(n677), 
        .QN(n3395) );
  DFFR_X1 \DRAM_mem_reg[24][28]  ( .D(n1442), .CK(CLK), .RN(n1009), .Q(n678), 
        .QN(n3396) );
  DFFR_X1 \DRAM_mem_reg[24][27]  ( .D(n1441), .CK(CLK), .RN(n1009), .Q(n679), 
        .QN(n3397) );
  DFFR_X1 \DRAM_mem_reg[24][26]  ( .D(n1440), .CK(CLK), .RN(n1009), .Q(n680), 
        .QN(n3398) );
  DFFR_X1 \DRAM_mem_reg[24][25]  ( .D(n1439), .CK(CLK), .RN(n1009), .Q(n681), 
        .QN(n3399) );
  DFFR_X1 \DRAM_mem_reg[24][24]  ( .D(n1438), .CK(CLK), .RN(n1009), .Q(n682), 
        .QN(n3400) );
  DFFR_X1 \DRAM_mem_reg[24][23]  ( .D(n1437), .CK(CLK), .RN(n1009), .Q(n683), 
        .QN(n3401) );
  DFFR_X1 \DRAM_mem_reg[24][22]  ( .D(n1436), .CK(CLK), .RN(n1009), .Q(n684), 
        .QN(n3402) );
  DFFR_X1 \DRAM_mem_reg[24][21]  ( .D(n1435), .CK(CLK), .RN(n1009), .Q(n685), 
        .QN(n3403) );
  DFFR_X1 \DRAM_mem_reg[24][20]  ( .D(n1434), .CK(CLK), .RN(n1009), .Q(n686), 
        .QN(n3404) );
  DFFR_X1 \DRAM_mem_reg[24][19]  ( .D(n1433), .CK(CLK), .RN(n1010), .Q(n687), 
        .QN(n3405) );
  DFFR_X1 \DRAM_mem_reg[24][18]  ( .D(n1432), .CK(CLK), .RN(n1010), .Q(n688), 
        .QN(n3406) );
  DFFR_X1 \DRAM_mem_reg[24][17]  ( .D(n1431), .CK(CLK), .RN(n1010), .Q(n689), 
        .QN(n3407) );
  DFFR_X1 \DRAM_mem_reg[24][16]  ( .D(n1430), .CK(CLK), .RN(n1010), .Q(n690), 
        .QN(n3408) );
  DFFR_X1 \DRAM_mem_reg[24][15]  ( .D(n1429), .CK(CLK), .RN(n1010), .Q(n925), 
        .QN(n3409) );
  DFFR_X1 \DRAM_mem_reg[24][14]  ( .D(n1428), .CK(CLK), .RN(n1010), .Q(n20) );
  DFFR_X1 \DRAM_mem_reg[24][13]  ( .D(n1427), .CK(CLK), .RN(n1010), .Q(n28) );
  DFFR_X1 \DRAM_mem_reg[24][12]  ( .D(n1426), .CK(CLK), .RN(n1010), .Q(n36) );
  DFFR_X1 \DRAM_mem_reg[24][11]  ( .D(n1425), .CK(CLK), .RN(n1010), .Q(n44) );
  DFFR_X1 \DRAM_mem_reg[24][10]  ( .D(n1424), .CK(CLK), .RN(n1010), .Q(n52) );
  DFFR_X1 \DRAM_mem_reg[24][9]  ( .D(n1423), .CK(CLK), .RN(n1010), .Q(n60) );
  DFFR_X1 \DRAM_mem_reg[24][8]  ( .D(n1422), .CK(CLK), .RN(n1010), .Q(n68) );
  DFFR_X1 \DRAM_mem_reg[24][7]  ( .D(n1421), .CK(CLK), .RN(n1011), .Q(n926), 
        .QN(n3410) );
  DFFR_X1 \DRAM_mem_reg[24][6]  ( .D(n1420), .CK(CLK), .RN(n1011), .Q(n927), 
        .QN(n3411) );
  DFFR_X1 \DRAM_mem_reg[24][5]  ( .D(n1419), .CK(CLK), .RN(n1011), .Q(n928), 
        .QN(n3412) );
  DFFR_X1 \DRAM_mem_reg[24][4]  ( .D(n1418), .CK(CLK), .RN(n1011), .Q(n929), 
        .QN(n3413) );
  DFFR_X1 \DRAM_mem_reg[24][3]  ( .D(n1417), .CK(CLK), .RN(n1011), .Q(n930), 
        .QN(n3414) );
  DFFR_X1 \DRAM_mem_reg[24][2]  ( .D(n1416), .CK(CLK), .RN(n1011), .Q(n931), 
        .QN(n3415) );
  DFFR_X1 \DRAM_mem_reg[24][1]  ( .D(n1415), .CK(CLK), .RN(n1011), .Q(n932), 
        .QN(n3416) );
  DFFR_X1 \DRAM_mem_reg[24][0]  ( .D(n1414), .CK(CLK), .RN(n1011), .Q(n933), 
        .QN(n3417) );
  DFFR_X1 \DRAM_mem_reg[25][31]  ( .D(n1413), .CK(CLK), .RN(n1011), .Q(n535), 
        .QN(n3418) );
  DFFR_X1 \DRAM_mem_reg[25][30]  ( .D(n1412), .CK(CLK), .RN(n1011), .Q(n536), 
        .QN(n3419) );
  DFFR_X1 \DRAM_mem_reg[25][29]  ( .D(n1411), .CK(CLK), .RN(n1011), .Q(n537), 
        .QN(n3420) );
  DFFR_X1 \DRAM_mem_reg[25][28]  ( .D(n1410), .CK(CLK), .RN(n1011), .Q(n538), 
        .QN(n3421) );
  DFFR_X1 \DRAM_mem_reg[25][27]  ( .D(n1409), .CK(CLK), .RN(n1012), .Q(n539), 
        .QN(n3422) );
  DFFR_X1 \DRAM_mem_reg[25][26]  ( .D(n1408), .CK(CLK), .RN(n1012), .Q(n540), 
        .QN(n3423) );
  DFFR_X1 \DRAM_mem_reg[25][25]  ( .D(n1407), .CK(CLK), .RN(n1012), .Q(n541), 
        .QN(n3424) );
  DFFR_X1 \DRAM_mem_reg[25][24]  ( .D(n1406), .CK(CLK), .RN(n1012), .Q(n542), 
        .QN(n3425) );
  DFFR_X1 \DRAM_mem_reg[25][23]  ( .D(n1405), .CK(CLK), .RN(n1012), .Q(n543), 
        .QN(n3426) );
  DFFR_X1 \DRAM_mem_reg[25][22]  ( .D(n1404), .CK(CLK), .RN(n1012), .Q(n544), 
        .QN(n3427) );
  DFFR_X1 \DRAM_mem_reg[25][21]  ( .D(n1403), .CK(CLK), .RN(n1012), .Q(n545), 
        .QN(n3428) );
  DFFR_X1 \DRAM_mem_reg[25][20]  ( .D(n1402), .CK(CLK), .RN(n1012), .Q(n546), 
        .QN(n3429) );
  DFFR_X1 \DRAM_mem_reg[25][19]  ( .D(n1401), .CK(CLK), .RN(n1012), .Q(n547), 
        .QN(n3430) );
  DFFR_X1 \DRAM_mem_reg[25][18]  ( .D(n1400), .CK(CLK), .RN(n1012), .Q(n548), 
        .QN(n3431) );
  DFFR_X1 \DRAM_mem_reg[25][17]  ( .D(n1399), .CK(CLK), .RN(n1012), .Q(n549), 
        .QN(n3432) );
  DFFR_X1 \DRAM_mem_reg[25][16]  ( .D(n1398), .CK(CLK), .RN(n1012), .Q(n550), 
        .QN(n3433) );
  DFFR_X1 \DRAM_mem_reg[25][15]  ( .D(n1397), .CK(CLK), .RN(n1013), .Q(n934), 
        .QN(n3434) );
  DFFR_X1 \DRAM_mem_reg[25][14]  ( .D(n1396), .CK(CLK), .RN(n1013), .Q(n256)
         );
  DFFR_X1 \DRAM_mem_reg[25][13]  ( .D(n1395), .CK(CLK), .RN(n1013), .Q(n264)
         );
  DFFR_X1 \DRAM_mem_reg[25][12]  ( .D(n1394), .CK(CLK), .RN(n1013), .Q(n272)
         );
  DFFR_X1 \DRAM_mem_reg[25][11]  ( .D(n1393), .CK(CLK), .RN(n1013), .Q(n280)
         );
  DFFR_X1 \DRAM_mem_reg[25][10]  ( .D(n1392), .CK(CLK), .RN(n1013), .Q(n288)
         );
  DFFR_X1 \DRAM_mem_reg[25][9]  ( .D(n1391), .CK(CLK), .RN(n1013), .Q(n296) );
  DFFR_X1 \DRAM_mem_reg[25][8]  ( .D(n1390), .CK(CLK), .RN(n1013), .Q(n304) );
  DFFR_X1 \DRAM_mem_reg[25][7]  ( .D(n1389), .CK(CLK), .RN(n1013), .Q(n805), 
        .QN(n3435) );
  DFFR_X1 \DRAM_mem_reg[25][6]  ( .D(n1388), .CK(CLK), .RN(n1013), .Q(n806), 
        .QN(n3436) );
  DFFR_X1 \DRAM_mem_reg[25][5]  ( .D(n1387), .CK(CLK), .RN(n1013), .Q(n807), 
        .QN(n3437) );
  DFFR_X1 \DRAM_mem_reg[25][4]  ( .D(n1386), .CK(CLK), .RN(n1013), .Q(n808), 
        .QN(n3438) );
  DFFR_X1 \DRAM_mem_reg[25][3]  ( .D(n1385), .CK(CLK), .RN(n1014), .Q(n809), 
        .QN(n3439) );
  DFFR_X1 \DRAM_mem_reg[25][2]  ( .D(n1384), .CK(CLK), .RN(n1014), .Q(n810), 
        .QN(n3440) );
  DFFR_X1 \DRAM_mem_reg[25][1]  ( .D(n1383), .CK(CLK), .RN(n1014), .Q(n811), 
        .QN(n3441) );
  DFFR_X1 \DRAM_mem_reg[25][0]  ( .D(n1382), .CK(CLK), .RN(n1014), .Q(n812), 
        .QN(n3442) );
  DFFR_X1 \DRAM_mem_reg[26][31]  ( .D(n1381), .CK(CLK), .RN(n1014), .Q(n551), 
        .QN(n3443) );
  DFFR_X1 \DRAM_mem_reg[26][30]  ( .D(n1380), .CK(CLK), .RN(n1014), .Q(n552), 
        .QN(n3444) );
  DFFR_X1 \DRAM_mem_reg[26][29]  ( .D(n1379), .CK(CLK), .RN(n1014), .Q(n553), 
        .QN(n3445) );
  DFFR_X1 \DRAM_mem_reg[26][28]  ( .D(n1378), .CK(CLK), .RN(n1014), .Q(n554), 
        .QN(n3446) );
  DFFR_X1 \DRAM_mem_reg[26][27]  ( .D(n1377), .CK(CLK), .RN(n1014), .Q(n555), 
        .QN(n3447) );
  DFFR_X1 \DRAM_mem_reg[26][26]  ( .D(n1376), .CK(CLK), .RN(n1014), .Q(n556), 
        .QN(n3448) );
  DFFR_X1 \DRAM_mem_reg[26][25]  ( .D(n1375), .CK(CLK), .RN(n1014), .Q(n557), 
        .QN(n3449) );
  DFFR_X1 \DRAM_mem_reg[26][24]  ( .D(n1374), .CK(CLK), .RN(n1014), .Q(n558), 
        .QN(n3450) );
  DFFR_X1 \DRAM_mem_reg[26][23]  ( .D(n1373), .CK(CLK), .RN(n1015), .Q(n559), 
        .QN(n3451) );
  DFFR_X1 \DRAM_mem_reg[26][22]  ( .D(n1372), .CK(CLK), .RN(n1015), .Q(n560), 
        .QN(n3452) );
  DFFR_X1 \DRAM_mem_reg[26][21]  ( .D(n1371), .CK(CLK), .RN(n1015), .Q(n561), 
        .QN(n3453) );
  DFFR_X1 \DRAM_mem_reg[26][20]  ( .D(n1370), .CK(CLK), .RN(n1015), .Q(n562), 
        .QN(n3454) );
  DFFR_X1 \DRAM_mem_reg[26][19]  ( .D(n1369), .CK(CLK), .RN(n1015), .Q(n563), 
        .QN(n3455) );
  DFFR_X1 \DRAM_mem_reg[26][18]  ( .D(n1368), .CK(CLK), .RN(n1015), .Q(n564), 
        .QN(n3456) );
  DFFR_X1 \DRAM_mem_reg[26][17]  ( .D(n1367), .CK(CLK), .RN(n1015), .Q(n565), 
        .QN(n3457) );
  DFFR_X1 \DRAM_mem_reg[26][16]  ( .D(n1366), .CK(CLK), .RN(n1015), .Q(n566), 
        .QN(n3458) );
  DFFR_X1 \DRAM_mem_reg[26][15]  ( .D(n1365), .CK(CLK), .RN(n1015), .Q(n935), 
        .QN(n3459) );
  DFFR_X1 \DRAM_mem_reg[26][14]  ( .D(n1364), .CK(CLK), .RN(n1015), .Q(n567), 
        .QN(n3460) );
  DFFR_X1 \DRAM_mem_reg[26][13]  ( .D(n1363), .CK(CLK), .RN(n1015), .Q(n568), 
        .QN(n3461) );
  DFFR_X1 \DRAM_mem_reg[26][12]  ( .D(n1362), .CK(CLK), .RN(n1015), .Q(n569), 
        .QN(n3462) );
  DFFR_X1 \DRAM_mem_reg[26][11]  ( .D(n1361), .CK(CLK), .RN(n1016), .Q(n570), 
        .QN(n3463) );
  DFFR_X1 \DRAM_mem_reg[26][10]  ( .D(n1360), .CK(CLK), .RN(n1016), .Q(n571), 
        .QN(n3464) );
  DFFR_X1 \DRAM_mem_reg[26][9]  ( .D(n1359), .CK(CLK), .RN(n1016), .Q(n572), 
        .QN(n3465) );
  DFFR_X1 \DRAM_mem_reg[26][8]  ( .D(n1358), .CK(CLK), .RN(n1016), .Q(n573), 
        .QN(n3466) );
  DFFR_X1 \DRAM_mem_reg[26][7]  ( .D(n1357), .CK(CLK), .RN(n1016), .Q(n367) );
  DFFR_X1 \DRAM_mem_reg[26][6]  ( .D(n1356), .CK(CLK), .RN(n1016), .Q(n371) );
  DFFR_X1 \DRAM_mem_reg[26][5]  ( .D(n1355), .CK(CLK), .RN(n1016), .Q(n375) );
  DFFR_X1 \DRAM_mem_reg[26][4]  ( .D(n1354), .CK(CLK), .RN(n1016), .Q(n379) );
  DFFR_X1 \DRAM_mem_reg[26][3]  ( .D(n1353), .CK(CLK), .RN(n1016), .Q(n383) );
  DFFR_X1 \DRAM_mem_reg[26][2]  ( .D(n1352), .CK(CLK), .RN(n1016), .Q(n387) );
  DFFR_X1 \DRAM_mem_reg[26][1]  ( .D(n1351), .CK(CLK), .RN(n1016), .Q(n391) );
  DFFR_X1 \DRAM_mem_reg[26][0]  ( .D(n1350), .CK(CLK), .RN(n1016), .Q(n395) );
  DFFR_X1 \DRAM_mem_reg[27][31]  ( .D(n1349), .CK(CLK), .RN(n1017), .Q(n221)
         );
  DFFR_X1 \DRAM_mem_reg[27][30]  ( .D(n1348), .CK(CLK), .RN(n1017), .Q(n222)
         );
  DFFR_X1 \DRAM_mem_reg[27][29]  ( .D(n1347), .CK(CLK), .RN(n1017), .Q(n223)
         );
  DFFR_X1 \DRAM_mem_reg[27][28]  ( .D(n1346), .CK(CLK), .RN(n1017), .Q(n224)
         );
  DFFR_X1 \DRAM_mem_reg[27][27]  ( .D(n1345), .CK(CLK), .RN(n1017), .Q(n225)
         );
  DFFR_X1 \DRAM_mem_reg[27][26]  ( .D(n1344), .CK(CLK), .RN(n1017), .Q(n226)
         );
  DFFR_X1 \DRAM_mem_reg[27][25]  ( .D(n1343), .CK(CLK), .RN(n1017), .Q(n227)
         );
  DFFR_X1 \DRAM_mem_reg[27][24]  ( .D(n1342), .CK(CLK), .RN(n1017), .Q(n228)
         );
  DFFR_X1 \DRAM_mem_reg[27][23]  ( .D(n1341), .CK(CLK), .RN(n1017), .Q(n229)
         );
  DFFR_X1 \DRAM_mem_reg[27][22]  ( .D(n1340), .CK(CLK), .RN(n1017), .Q(n230)
         );
  DFFR_X1 \DRAM_mem_reg[27][21]  ( .D(n1339), .CK(CLK), .RN(n1017), .Q(n231)
         );
  DFFR_X1 \DRAM_mem_reg[27][20]  ( .D(n1338), .CK(CLK), .RN(n1017), .Q(n232)
         );
  DFFR_X1 \DRAM_mem_reg[27][19]  ( .D(n1337), .CK(CLK), .RN(n1018), .Q(n233)
         );
  DFFR_X1 \DRAM_mem_reg[27][18]  ( .D(n1336), .CK(CLK), .RN(n1018), .Q(n234)
         );
  DFFR_X1 \DRAM_mem_reg[27][17]  ( .D(n1335), .CK(CLK), .RN(n1018), .Q(n235)
         );
  DFFR_X1 \DRAM_mem_reg[27][16]  ( .D(n1334), .CK(CLK), .RN(n1018), .Q(n236)
         );
  DFFR_X1 \DRAM_mem_reg[27][15]  ( .D(n1333), .CK(CLK), .RN(n1018), .Q(n936), 
        .QN(n3467) );
  DFFR_X1 \DRAM_mem_reg[27][14]  ( .D(n1332), .CK(CLK), .RN(n1018), .Q(n691), 
        .QN(n3468) );
  DFFR_X1 \DRAM_mem_reg[27][13]  ( .D(n1331), .CK(CLK), .RN(n1018), .Q(n692), 
        .QN(n3469) );
  DFFR_X1 \DRAM_mem_reg[27][12]  ( .D(n1330), .CK(CLK), .RN(n1018), .Q(n693), 
        .QN(n3470) );
  DFFR_X1 \DRAM_mem_reg[27][11]  ( .D(n1329), .CK(CLK), .RN(n1018), .Q(n694), 
        .QN(n3471) );
  DFFR_X1 \DRAM_mem_reg[27][10]  ( .D(n1328), .CK(CLK), .RN(n1018), .Q(n695), 
        .QN(n3472) );
  DFFR_X1 \DRAM_mem_reg[27][9]  ( .D(n1327), .CK(CLK), .RN(n1018), .Q(n696), 
        .QN(n3473) );
  DFFR_X1 \DRAM_mem_reg[27][8]  ( .D(n1326), .CK(CLK), .RN(n1018), .Q(n697), 
        .QN(n3474) );
  DFFR_X1 \DRAM_mem_reg[27][7]  ( .D(n1325), .CK(CLK), .RN(n1019), .Q(n131) );
  DFFR_X1 \DRAM_mem_reg[27][6]  ( .D(n1324), .CK(CLK), .RN(n1019), .Q(n135) );
  DFFR_X1 \DRAM_mem_reg[27][5]  ( .D(n1323), .CK(CLK), .RN(n1019), .Q(n139) );
  DFFR_X1 \DRAM_mem_reg[27][4]  ( .D(n1322), .CK(CLK), .RN(n1019), .Q(n143) );
  DFFR_X1 \DRAM_mem_reg[27][3]  ( .D(n1321), .CK(CLK), .RN(n1019), .Q(n147) );
  DFFR_X1 \DRAM_mem_reg[27][2]  ( .D(n1320), .CK(CLK), .RN(n1019), .Q(n151) );
  DFFR_X1 \DRAM_mem_reg[27][1]  ( .D(n1319), .CK(CLK), .RN(n1019), .Q(n155) );
  DFFR_X1 \DRAM_mem_reg[27][0]  ( .D(n1318), .CK(CLK), .RN(n1019), .Q(n159) );
  DFFR_X1 \DRAM_mem_reg[28][31]  ( .D(n1317), .CK(CLK), .RN(n1019), .Q(n237)
         );
  DFFR_X1 \DRAM_mem_reg[28][30]  ( .D(n1316), .CK(CLK), .RN(n1019), .Q(n238)
         );
  DFFR_X1 \DRAM_mem_reg[28][29]  ( .D(n1315), .CK(CLK), .RN(n1019), .Q(n239)
         );
  DFFR_X1 \DRAM_mem_reg[28][28]  ( .D(n1314), .CK(CLK), .RN(n1019), .Q(n240)
         );
  DFFR_X1 \DRAM_mem_reg[28][27]  ( .D(n1313), .CK(CLK), .RN(n1020), .Q(n241)
         );
  DFFR_X1 \DRAM_mem_reg[28][26]  ( .D(n1312), .CK(CLK), .RN(n1020), .Q(n242)
         );
  DFFR_X1 \DRAM_mem_reg[28][25]  ( .D(n1311), .CK(CLK), .RN(n1020), .Q(n243)
         );
  DFFR_X1 \DRAM_mem_reg[28][24]  ( .D(n1310), .CK(CLK), .RN(n1020), .Q(n244)
         );
  DFFR_X1 \DRAM_mem_reg[28][23]  ( .D(n1309), .CK(CLK), .RN(n1020), .Q(n245)
         );
  DFFR_X1 \DRAM_mem_reg[28][22]  ( .D(n1308), .CK(CLK), .RN(n1020), .Q(n246)
         );
  DFFR_X1 \DRAM_mem_reg[28][21]  ( .D(n1307), .CK(CLK), .RN(n1020), .Q(n247)
         );
  DFFR_X1 \DRAM_mem_reg[28][20]  ( .D(n1306), .CK(CLK), .RN(n1020), .Q(n248)
         );
  DFFR_X1 \DRAM_mem_reg[28][19]  ( .D(n1305), .CK(CLK), .RN(n1020), .Q(n249)
         );
  DFFR_X1 \DRAM_mem_reg[28][18]  ( .D(n1304), .CK(CLK), .RN(n1020), .Q(n250)
         );
  DFFR_X1 \DRAM_mem_reg[28][17]  ( .D(n1303), .CK(CLK), .RN(n1020), .Q(n251)
         );
  DFFR_X1 \DRAM_mem_reg[28][16]  ( .D(n1302), .CK(CLK), .RN(n1020), .Q(n252)
         );
  DFFR_X1 \DRAM_mem_reg[28][15]  ( .D(n1301), .CK(CLK), .RN(n1021), .Q(n813), 
        .QN(n3475) );
  DFFR_X1 \DRAM_mem_reg[28][14]  ( .D(n1300), .CK(CLK), .RN(n1021), .Q(n19) );
  DFFR_X1 \DRAM_mem_reg[28][13]  ( .D(n1299), .CK(CLK), .RN(n1021), .Q(n27) );
  DFFR_X1 \DRAM_mem_reg[28][12]  ( .D(n1298), .CK(CLK), .RN(n1021), .Q(n35) );
  DFFR_X1 \DRAM_mem_reg[28][11]  ( .D(n1297), .CK(CLK), .RN(n1021), .Q(n43) );
  DFFR_X1 \DRAM_mem_reg[28][10]  ( .D(n1296), .CK(CLK), .RN(n1021), .Q(n51) );
  DFFR_X1 \DRAM_mem_reg[28][9]  ( .D(n1295), .CK(CLK), .RN(n1021), .Q(n59) );
  DFFR_X1 \DRAM_mem_reg[28][8]  ( .D(n1294), .CK(CLK), .RN(n1021), .Q(n67) );
  DFFR_X1 \DRAM_mem_reg[28][7]  ( .D(n1293), .CK(CLK), .RN(n1021), .Q(n937), 
        .QN(n3476) );
  DFFR_X1 \DRAM_mem_reg[28][6]  ( .D(n1292), .CK(CLK), .RN(n1021), .Q(n938), 
        .QN(n3477) );
  DFFR_X1 \DRAM_mem_reg[28][5]  ( .D(n1291), .CK(CLK), .RN(n1021), .Q(n939), 
        .QN(n3478) );
  DFFR_X1 \DRAM_mem_reg[28][4]  ( .D(n1290), .CK(CLK), .RN(n1021), .Q(n940), 
        .QN(n3479) );
  DFFR_X1 \DRAM_mem_reg[28][3]  ( .D(n1289), .CK(CLK), .RN(n1022), .Q(n941), 
        .QN(n3480) );
  DFFR_X1 \DRAM_mem_reg[28][2]  ( .D(n1288), .CK(CLK), .RN(n1022), .Q(n942), 
        .QN(n3481) );
  DFFR_X1 \DRAM_mem_reg[28][1]  ( .D(n1287), .CK(CLK), .RN(n1022), .Q(n943), 
        .QN(n3482) );
  DFFR_X1 \DRAM_mem_reg[28][0]  ( .D(n1286), .CK(CLK), .RN(n1022), .Q(n944), 
        .QN(n3483) );
  DFFR_X1 \DRAM_mem_reg[29][31]  ( .D(n1285), .CK(CLK), .RN(n1022), .Q(n574), 
        .QN(n3484) );
  DFFR_X1 \DRAM_mem_reg[29][30]  ( .D(n1284), .CK(CLK), .RN(n1022), .Q(n575), 
        .QN(n3485) );
  DFFR_X1 \DRAM_mem_reg[29][29]  ( .D(n1283), .CK(CLK), .RN(n1022), .Q(n576), 
        .QN(n3486) );
  DFFR_X1 \DRAM_mem_reg[29][28]  ( .D(n1282), .CK(CLK), .RN(n1022), .Q(n577), 
        .QN(n3487) );
  DFFR_X1 \DRAM_mem_reg[29][27]  ( .D(n1281), .CK(CLK), .RN(n1022), .Q(n578), 
        .QN(n3488) );
  DFFR_X1 \DRAM_mem_reg[29][26]  ( .D(n1280), .CK(CLK), .RN(n1022), .Q(n579), 
        .QN(n3489) );
  DFFR_X1 \DRAM_mem_reg[29][25]  ( .D(n1279), .CK(CLK), .RN(n1022), .Q(n580), 
        .QN(n3490) );
  DFFR_X1 \DRAM_mem_reg[29][24]  ( .D(n1278), .CK(CLK), .RN(n1022), .Q(n581), 
        .QN(n3491) );
  DFFR_X1 \DRAM_mem_reg[29][23]  ( .D(n1277), .CK(CLK), .RN(n1023), .Q(n582), 
        .QN(n3492) );
  DFFR_X1 \DRAM_mem_reg[29][22]  ( .D(n1276), .CK(CLK), .RN(n1023), .Q(n583), 
        .QN(n3493) );
  DFFR_X1 \DRAM_mem_reg[29][21]  ( .D(n1275), .CK(CLK), .RN(n1023), .Q(n584), 
        .QN(n3494) );
  DFFR_X1 \DRAM_mem_reg[29][20]  ( .D(n1274), .CK(CLK), .RN(n1023), .Q(n585), 
        .QN(n3495) );
  DFFR_X1 \DRAM_mem_reg[29][19]  ( .D(n1273), .CK(CLK), .RN(n1023), .Q(n586), 
        .QN(n3496) );
  DFFR_X1 \DRAM_mem_reg[29][18]  ( .D(n1272), .CK(CLK), .RN(n1023), .Q(n587), 
        .QN(n3497) );
  DFFR_X1 \DRAM_mem_reg[29][17]  ( .D(n1271), .CK(CLK), .RN(n1023), .Q(n588), 
        .QN(n3498) );
  DFFR_X1 \DRAM_mem_reg[29][16]  ( .D(n1270), .CK(CLK), .RN(n1023), .Q(n589), 
        .QN(n3499) );
  DFFR_X1 \DRAM_mem_reg[29][15]  ( .D(n1269), .CK(CLK), .RN(n1023), .Q(n814), 
        .QN(n3500) );
  DFFR_X1 \DRAM_mem_reg[29][14]  ( .D(n1268), .CK(CLK), .RN(n1023), .Q(n255)
         );
  DFFR_X1 \DRAM_mem_reg[29][13]  ( .D(n1267), .CK(CLK), .RN(n1023), .Q(n263)
         );
  DFFR_X1 \DRAM_mem_reg[29][12]  ( .D(n1266), .CK(CLK), .RN(n1023), .Q(n271)
         );
  DFFR_X1 \DRAM_mem_reg[29][11]  ( .D(n1265), .CK(CLK), .RN(n1024), .Q(n279)
         );
  DFFR_X1 \DRAM_mem_reg[29][10]  ( .D(n1264), .CK(CLK), .RN(n1024), .Q(n287)
         );
  DFFR_X1 \DRAM_mem_reg[29][9]  ( .D(n1263), .CK(CLK), .RN(n1024), .Q(n295) );
  DFFR_X1 \DRAM_mem_reg[29][8]  ( .D(n1262), .CK(CLK), .RN(n1024), .Q(n303) );
  DFFR_X1 \DRAM_mem_reg[29][7]  ( .D(n1261), .CK(CLK), .RN(n1024), .Q(n815), 
        .QN(n3501) );
  DFFR_X1 \DRAM_mem_reg[29][6]  ( .D(n1260), .CK(CLK), .RN(n1024), .Q(n816), 
        .QN(n3502) );
  DFFR_X1 \DRAM_mem_reg[29][5]  ( .D(n1259), .CK(CLK), .RN(n1024), .Q(n817), 
        .QN(n3503) );
  DFFR_X1 \DRAM_mem_reg[29][4]  ( .D(n1258), .CK(CLK), .RN(n1024), .Q(n818), 
        .QN(n3504) );
  DFFR_X1 \DRAM_mem_reg[29][3]  ( .D(n1257), .CK(CLK), .RN(n1024), .Q(n819), 
        .QN(n3505) );
  DFFR_X1 \DRAM_mem_reg[29][2]  ( .D(n1256), .CK(CLK), .RN(n1024), .Q(n820), 
        .QN(n3506) );
  DFFR_X1 \DRAM_mem_reg[29][1]  ( .D(n1255), .CK(CLK), .RN(n1024), .Q(n821), 
        .QN(n3507) );
  DFFR_X1 \DRAM_mem_reg[29][0]  ( .D(n1254), .CK(CLK), .RN(n1024), .Q(n822), 
        .QN(n3508) );
  DFFR_X1 \DRAM_mem_reg[30][31]  ( .D(n1253), .CK(CLK), .RN(n1025), .Q(n1) );
  DFFR_X1 \DRAM_mem_reg[30][30]  ( .D(n1252), .CK(CLK), .RN(n1025), .Q(n2) );
  DFFR_X1 \DRAM_mem_reg[30][29]  ( .D(n1251), .CK(CLK), .RN(n1025), .Q(n3) );
  DFFR_X1 \DRAM_mem_reg[30][28]  ( .D(n1250), .CK(CLK), .RN(n1025), .Q(n4) );
  DFFR_X1 \DRAM_mem_reg[30][27]  ( .D(n1249), .CK(CLK), .RN(n1025), .Q(n5) );
  DFFR_X1 \DRAM_mem_reg[30][26]  ( .D(n1248), .CK(CLK), .RN(n1025), .Q(n6) );
  DFFR_X1 \DRAM_mem_reg[30][25]  ( .D(n1247), .CK(CLK), .RN(n1025), .Q(n7) );
  DFFR_X1 \DRAM_mem_reg[30][24]  ( .D(n1246), .CK(CLK), .RN(n1025), .Q(n8) );
  DFFR_X1 \DRAM_mem_reg[30][23]  ( .D(n1245), .CK(CLK), .RN(n1025), .Q(n9) );
  DFFR_X1 \DRAM_mem_reg[30][22]  ( .D(n1244), .CK(CLK), .RN(n1025), .Q(n10) );
  DFFR_X1 \DRAM_mem_reg[30][21]  ( .D(n1243), .CK(CLK), .RN(n1025), .Q(n11) );
  DFFR_X1 \DRAM_mem_reg[30][20]  ( .D(n1242), .CK(CLK), .RN(n1025), .Q(n12) );
  DFFR_X1 \DRAM_mem_reg[30][19]  ( .D(n1241), .CK(CLK), .RN(n1026), .Q(n13) );
  DFFR_X1 \DRAM_mem_reg[30][18]  ( .D(n1240), .CK(CLK), .RN(n1026), .Q(n14) );
  DFFR_X1 \DRAM_mem_reg[30][17]  ( .D(n1239), .CK(CLK), .RN(n1026), .Q(n15) );
  DFFR_X1 \DRAM_mem_reg[30][16]  ( .D(n1238), .CK(CLK), .RN(n1026), .Q(n16) );
  DFFR_X1 \DRAM_mem_reg[30][15]  ( .D(n1237), .CK(CLK), .RN(n1026), .Q(n823), 
        .QN(n3509) );
  DFFR_X1 \DRAM_mem_reg[30][14]  ( .D(n1236), .CK(CLK), .RN(n1026), .Q(n590), 
        .QN(n3510) );
  DFFR_X1 \DRAM_mem_reg[30][13]  ( .D(n1235), .CK(CLK), .RN(n1026), .Q(n591), 
        .QN(n3511) );
  DFFR_X1 \DRAM_mem_reg[30][12]  ( .D(n1234), .CK(CLK), .RN(n1026), .Q(n592), 
        .QN(n3512) );
  DFFR_X1 \DRAM_mem_reg[30][11]  ( .D(n1233), .CK(CLK), .RN(n1026), .Q(n593), 
        .QN(n3513) );
  DFFR_X1 \DRAM_mem_reg[30][10]  ( .D(n1232), .CK(CLK), .RN(n1026), .Q(n594), 
        .QN(n3514) );
  DFFR_X1 \DRAM_mem_reg[30][9]  ( .D(n1231), .CK(CLK), .RN(n1026), .Q(n595), 
        .QN(n3515) );
  DFFR_X1 \DRAM_mem_reg[30][8]  ( .D(n1230), .CK(CLK), .RN(n1026), .Q(n596), 
        .QN(n3516) );
  DFFR_X1 \DRAM_mem_reg[30][7]  ( .D(n1229), .CK(CLK), .RN(n1027), .Q(n368) );
  DFFR_X1 \DRAM_mem_reg[30][6]  ( .D(n1228), .CK(CLK), .RN(n1027), .Q(n372) );
  DFFR_X1 \DRAM_mem_reg[30][5]  ( .D(n1227), .CK(CLK), .RN(n1027), .Q(n376) );
  DFFR_X1 \DRAM_mem_reg[30][4]  ( .D(n1226), .CK(CLK), .RN(n1027), .Q(n380) );
  DFFR_X1 \DRAM_mem_reg[30][3]  ( .D(n1225), .CK(CLK), .RN(n1027), .Q(n384) );
  DFFR_X1 \DRAM_mem_reg[30][2]  ( .D(n1224), .CK(CLK), .RN(n1027), .Q(n388) );
  DFFR_X1 \DRAM_mem_reg[30][1]  ( .D(n1223), .CK(CLK), .RN(n1027), .Q(n392) );
  DFFR_X1 \DRAM_mem_reg[30][0]  ( .D(n1222), .CK(CLK), .RN(n1027), .Q(n396) );
  DFFR_X1 \DRAM_mem_reg[31][31]  ( .D(n1221), .CK(CLK), .RN(n1027), .Q(n698), 
        .QN(n3517) );
  DFFR_X1 \DRAM_mem_reg[31][30]  ( .D(n1220), .CK(CLK), .RN(n1027), .Q(n699), 
        .QN(n3518) );
  DFFR_X1 \DRAM_mem_reg[31][29]  ( .D(n1219), .CK(CLK), .RN(n1027), .Q(n700), 
        .QN(n3519) );
  DFFR_X1 \DRAM_mem_reg[31][28]  ( .D(n1218), .CK(CLK), .RN(n1027), .Q(n701), 
        .QN(n3520) );
  DFFR_X1 \DRAM_mem_reg[31][27]  ( .D(n1217), .CK(CLK), .RN(n1028), .Q(n702), 
        .QN(n3521) );
  DFFR_X1 \DRAM_mem_reg[31][26]  ( .D(n1216), .CK(CLK), .RN(n1028), .Q(n703), 
        .QN(n3522) );
  DFFR_X1 \DRAM_mem_reg[31][25]  ( .D(n1215), .CK(CLK), .RN(n1028), .Q(n704), 
        .QN(n3523) );
  DFFR_X1 \DRAM_mem_reg[31][24]  ( .D(n1214), .CK(CLK), .RN(n1028), .Q(n705), 
        .QN(n3524) );
  DFFR_X1 \DRAM_mem_reg[31][23]  ( .D(n1213), .CK(CLK), .RN(n1028), .Q(n706), 
        .QN(n3525) );
  DFFR_X1 \DRAM_mem_reg[31][22]  ( .D(n1212), .CK(CLK), .RN(n1028), .Q(n707), 
        .QN(n3526) );
  DFFR_X1 \DRAM_mem_reg[31][21]  ( .D(n1211), .CK(CLK), .RN(n1028), .Q(n708), 
        .QN(n3527) );
  DFFR_X1 \DRAM_mem_reg[31][20]  ( .D(n1210), .CK(CLK), .RN(n1028), .Q(n709), 
        .QN(n3528) );
  DFFR_X1 \DRAM_mem_reg[31][19]  ( .D(n1209), .CK(CLK), .RN(n1028), .Q(n710), 
        .QN(n3529) );
  DFFR_X1 \DRAM_mem_reg[31][18]  ( .D(n1208), .CK(CLK), .RN(n1028), .Q(n711), 
        .QN(n3530) );
  DFFR_X1 \DRAM_mem_reg[31][17]  ( .D(n1207), .CK(CLK), .RN(n1028), .Q(n712), 
        .QN(n3531) );
  DFFR_X1 \DRAM_mem_reg[31][16]  ( .D(n1206), .CK(CLK), .RN(n1028), .Q(n713), 
        .QN(n3532) );
  DFFR_X1 \DRAM_mem_reg[31][15]  ( .D(n1205), .CK(CLK), .RN(n1029), .Q(n824), 
        .QN(n3533) );
  DFFR_X1 \DRAM_mem_reg[31][14]  ( .D(n1204), .CK(CLK), .RN(n1029), .Q(n714), 
        .QN(n3534) );
  DFFR_X1 \DRAM_mem_reg[31][13]  ( .D(n1203), .CK(CLK), .RN(n1029), .Q(n715), 
        .QN(n3535) );
  DFFR_X1 \DRAM_mem_reg[31][12]  ( .D(n1202), .CK(CLK), .RN(n1029), .Q(n716), 
        .QN(n3536) );
  DFFR_X1 \DRAM_mem_reg[31][11]  ( .D(n1201), .CK(CLK), .RN(n1029), .Q(n717), 
        .QN(n3537) );
  DFFR_X1 \DRAM_mem_reg[31][10]  ( .D(n1200), .CK(CLK), .RN(n1029), .Q(n718), 
        .QN(n3538) );
  DFFR_X1 \DRAM_mem_reg[31][9]  ( .D(n1199), .CK(CLK), .RN(n1029), .Q(n719), 
        .QN(n3539) );
  DFFR_X1 \DRAM_mem_reg[31][8]  ( .D(n1198), .CK(CLK), .RN(n1029), .Q(n720), 
        .QN(n3540) );
  DFFR_X1 \DRAM_mem_reg[31][7]  ( .D(n1197), .CK(CLK), .RN(n1029), .Q(n132) );
  DFFR_X1 \DRAM_mem_reg[31][6]  ( .D(n1196), .CK(CLK), .RN(n1029), .Q(n136) );
  DFFR_X1 \DRAM_mem_reg[31][5]  ( .D(n1195), .CK(CLK), .RN(n1029), .Q(n140) );
  DFFR_X1 \DRAM_mem_reg[31][4]  ( .D(n1194), .CK(CLK), .RN(n1029), .Q(n144) );
  DFFR_X1 \DRAM_mem_reg[31][3]  ( .D(n1193), .CK(CLK), .RN(n1030), .Q(n148) );
  DFFR_X1 \DRAM_mem_reg[31][2]  ( .D(n1192), .CK(CLK), .RN(n1030), .Q(n152) );
  DFFR_X1 \DRAM_mem_reg[31][1]  ( .D(n1191), .CK(CLK), .RN(n1030), .Q(n156) );
  DFFR_X1 \DRAM_mem_reg[31][0]  ( .D(n1190), .CK(CLK), .RN(n1030), .Q(n160) );
  AND2_X2 U8141 ( .A1(n2464), .A2(n2403), .ZN(n2465) );
  AND2_X2 U8142 ( .A1(n2458), .A2(n2411), .ZN(n2461) );
  AND2_X2 U8143 ( .A1(n2464), .A2(n2410), .ZN(n2466) );
  AND2_X2 U8144 ( .A1(n2471), .A2(n2409), .ZN(n2470) );
  AND2_X2 U8145 ( .A1(n2458), .A2(n2403), .ZN(n2459) );
  AND2_X2 U8146 ( .A1(n2464), .A2(n2411), .ZN(n2467) );
  AND2_X2 U8147 ( .A1(n2477), .A2(n2409), .ZN(n2476) );
  AND2_X2 U8148 ( .A1(n2482), .A2(n2410), .ZN(n2484) );
  AND2_X2 U8149 ( .A1(n2482), .A2(n2403), .ZN(n2483) );
  AND2_X2 U8150 ( .A1(n2487), .A2(n2411), .ZN(n2490) );
  AND2_X2 U8151 ( .A1(n2471), .A2(n2410), .ZN(n2473) );
  AND2_X2 U8152 ( .A1(n2445), .A2(n2409), .ZN(n2413) );
  AND2_X2 U8153 ( .A1(n2487), .A2(n2403), .ZN(n2488) );
  AND2_X2 U8154 ( .A1(n2471), .A2(n2411), .ZN(n2474) );
  AND2_X2 U8155 ( .A1(n2477), .A2(n2410), .ZN(n2479) );
  AND2_X2 U8156 ( .A1(n2452), .A2(n2409), .ZN(n2451) );
  AND2_X2 U8157 ( .A1(n2477), .A2(n2411), .ZN(n2480) );
  AND2_X2 U8158 ( .A1(n2458), .A2(n2409), .ZN(n2457) );
  AND2_X2 U8159 ( .A1(n2452), .A2(n2403), .ZN(n2453) );
  AND2_X2 U8160 ( .A1(n2445), .A2(n2410), .ZN(n2447) );
  AND2_X2 U8161 ( .A1(n2487), .A2(n2409), .ZN(n2486) );
  AND2_X2 U8162 ( .A1(n2445), .A2(n2403), .ZN(n2446) );
  AND2_X2 U8163 ( .A1(n2482), .A2(n2411), .ZN(n2485) );
  AND2_X2 U8164 ( .A1(n2452), .A2(n2410), .ZN(n2454) );
  OAI21_X2 U8165 ( .B1(n2405), .B2(n2406), .A(n2407), .ZN(n1094) );
  AND2_X2 U8166 ( .A1(n2482), .A2(n2409), .ZN(n2481) );
  AND2_X2 U8167 ( .A1(n2477), .A2(n2403), .ZN(n2478) );
  AND2_X2 U8168 ( .A1(n2464), .A2(n2409), .ZN(n2463) );
  NOR2_X2 U8169 ( .A1(Addr[0]), .A2(Addr[1]), .ZN(n2409) );
  AND2_X2 U8170 ( .A1(n2458), .A2(n2410), .ZN(n2460) );
  AND2_X2 U8171 ( .A1(n2471), .A2(n2403), .ZN(n2472) );
  NOR2_X2 U8172 ( .A1(n2884), .A2(Addr[1]), .ZN(n2403) );
  AND2_X2 U8173 ( .A1(n2487), .A2(n2410), .ZN(n2489) );
  NOR2_X2 U8174 ( .A1(n2883), .A2(Addr[0]), .ZN(n2410) );
  AND2_X2 U8175 ( .A1(n2445), .A2(n2411), .ZN(n2448) );
  AND2_X2 U8176 ( .A1(n2452), .A2(n2411), .ZN(n2455) );
  NOR2_X2 U8177 ( .A1(n2884), .A2(n2883), .ZN(n2411) );
  BUF_X1 U8178 ( .A(n13687), .Z(n1031) );
  BUF_X1 U8179 ( .A(n13687), .Z(n1032) );
  BUF_X1 U8180 ( .A(n13687), .Z(n1033) );
  BUF_X1 U8181 ( .A(n13687), .Z(n1034) );
  BUF_X1 U8182 ( .A(n13687), .Z(n1035) );
  BUF_X1 U8183 ( .A(n13687), .Z(n1036) );
  BUF_X1 U8184 ( .A(n13687), .Z(n1037) );
  BUF_X1 U8185 ( .A(n13687), .Z(n1038) );
  BUF_X1 U8186 ( .A(n13687), .Z(n1039) );
  BUF_X1 U8187 ( .A(n13687), .Z(n1040) );
  BUF_X1 U8188 ( .A(n13687), .Z(n1041) );
  BUF_X1 U8189 ( .A(n13687), .Z(n1042) );
  BUF_X1 U8190 ( .A(n13687), .Z(n1043) );
  BUF_X1 U8191 ( .A(n13687), .Z(n1044) );
  BUF_X1 U8192 ( .A(n13687), .Z(n1045) );
  CLKBUF_X1 U8193 ( .A(n1045), .Z(n945) );
  CLKBUF_X1 U8194 ( .A(n1045), .Z(n946) );
  CLKBUF_X1 U8195 ( .A(n1044), .Z(n947) );
  CLKBUF_X1 U8196 ( .A(n1044), .Z(n948) );
  CLKBUF_X1 U8197 ( .A(n1044), .Z(n949) );
  CLKBUF_X1 U8198 ( .A(n1044), .Z(n950) );
  CLKBUF_X1 U8199 ( .A(n1044), .Z(n951) );
  CLKBUF_X1 U8200 ( .A(n1044), .Z(n952) );
  CLKBUF_X1 U8201 ( .A(n1043), .Z(n953) );
  CLKBUF_X1 U8202 ( .A(n1043), .Z(n954) );
  CLKBUF_X1 U8203 ( .A(n1043), .Z(n955) );
  CLKBUF_X1 U8204 ( .A(n1043), .Z(n956) );
  CLKBUF_X1 U8205 ( .A(n1043), .Z(n957) );
  CLKBUF_X1 U8206 ( .A(n1043), .Z(n958) );
  CLKBUF_X1 U8207 ( .A(n1042), .Z(n959) );
  CLKBUF_X1 U8208 ( .A(n1042), .Z(n960) );
  CLKBUF_X1 U8209 ( .A(n1042), .Z(n961) );
  CLKBUF_X1 U8210 ( .A(n1042), .Z(n962) );
  CLKBUF_X1 U8211 ( .A(n1042), .Z(n963) );
  CLKBUF_X1 U8212 ( .A(n1042), .Z(n964) );
  CLKBUF_X1 U8213 ( .A(n1041), .Z(n965) );
  CLKBUF_X1 U8214 ( .A(n1041), .Z(n966) );
  CLKBUF_X1 U8215 ( .A(n1041), .Z(n967) );
  CLKBUF_X1 U8216 ( .A(n1041), .Z(n968) );
  CLKBUF_X1 U8217 ( .A(n1041), .Z(n969) );
  CLKBUF_X1 U8218 ( .A(n1041), .Z(n970) );
  CLKBUF_X1 U8219 ( .A(n1040), .Z(n971) );
  CLKBUF_X1 U8220 ( .A(n1040), .Z(n972) );
  CLKBUF_X1 U8221 ( .A(n1040), .Z(n973) );
  CLKBUF_X1 U8222 ( .A(n1040), .Z(n974) );
  CLKBUF_X1 U8223 ( .A(n1040), .Z(n975) );
  CLKBUF_X1 U8224 ( .A(n1040), .Z(n976) );
  CLKBUF_X1 U8225 ( .A(n1039), .Z(n977) );
  CLKBUF_X1 U8226 ( .A(n1039), .Z(n978) );
  CLKBUF_X1 U8227 ( .A(n1039), .Z(n979) );
  CLKBUF_X1 U8228 ( .A(n1039), .Z(n980) );
  CLKBUF_X1 U8229 ( .A(n1039), .Z(n981) );
  CLKBUF_X1 U8230 ( .A(n1039), .Z(n982) );
  CLKBUF_X1 U8231 ( .A(n1038), .Z(n983) );
  CLKBUF_X1 U8232 ( .A(n1038), .Z(n984) );
  CLKBUF_X1 U8233 ( .A(n1038), .Z(n985) );
  CLKBUF_X1 U8234 ( .A(n1038), .Z(n986) );
  CLKBUF_X1 U8235 ( .A(n1038), .Z(n987) );
  CLKBUF_X1 U8236 ( .A(n1038), .Z(n988) );
  CLKBUF_X1 U8237 ( .A(n1037), .Z(n989) );
  CLKBUF_X1 U8238 ( .A(n1037), .Z(n990) );
  CLKBUF_X1 U8239 ( .A(n1037), .Z(n991) );
  CLKBUF_X1 U8240 ( .A(n1037), .Z(n992) );
  CLKBUF_X1 U8241 ( .A(n1037), .Z(n993) );
  CLKBUF_X1 U8242 ( .A(n1037), .Z(n994) );
  CLKBUF_X1 U8243 ( .A(n1036), .Z(n995) );
  CLKBUF_X1 U8244 ( .A(n1036), .Z(n996) );
  CLKBUF_X1 U8245 ( .A(n1036), .Z(n997) );
  CLKBUF_X1 U8246 ( .A(n1036), .Z(n998) );
  CLKBUF_X1 U8247 ( .A(n1036), .Z(n999) );
  CLKBUF_X1 U8248 ( .A(n1036), .Z(n1000) );
  CLKBUF_X1 U8249 ( .A(n1035), .Z(n1001) );
  CLKBUF_X1 U8250 ( .A(n1035), .Z(n1002) );
  CLKBUF_X1 U8251 ( .A(n1035), .Z(n1003) );
  CLKBUF_X1 U8252 ( .A(n1035), .Z(n1004) );
  CLKBUF_X1 U8253 ( .A(n1035), .Z(n1005) );
  CLKBUF_X1 U8254 ( .A(n1035), .Z(n1006) );
  CLKBUF_X1 U8255 ( .A(n1034), .Z(n1007) );
  CLKBUF_X1 U8256 ( .A(n1034), .Z(n1008) );
  CLKBUF_X1 U8257 ( .A(n1034), .Z(n1009) );
  CLKBUF_X1 U8258 ( .A(n1034), .Z(n1010) );
  CLKBUF_X1 U8259 ( .A(n1034), .Z(n1011) );
  CLKBUF_X1 U8260 ( .A(n1034), .Z(n1012) );
  CLKBUF_X1 U8261 ( .A(n1033), .Z(n1013) );
  CLKBUF_X1 U8262 ( .A(n1033), .Z(n1014) );
  CLKBUF_X1 U8263 ( .A(n1033), .Z(n1015) );
  CLKBUF_X1 U8264 ( .A(n1033), .Z(n1016) );
  CLKBUF_X1 U8265 ( .A(n1033), .Z(n1017) );
  CLKBUF_X1 U8266 ( .A(n1033), .Z(n1018) );
  CLKBUF_X1 U8267 ( .A(n1032), .Z(n1019) );
  CLKBUF_X1 U8268 ( .A(n1032), .Z(n1020) );
  CLKBUF_X1 U8269 ( .A(n1032), .Z(n1021) );
  CLKBUF_X1 U8270 ( .A(n1032), .Z(n1022) );
  CLKBUF_X1 U8271 ( .A(n1032), .Z(n1023) );
  CLKBUF_X1 U8272 ( .A(n1032), .Z(n1024) );
  CLKBUF_X1 U8273 ( .A(n1031), .Z(n1025) );
  CLKBUF_X1 U8274 ( .A(n1031), .Z(n1026) );
  CLKBUF_X1 U8275 ( .A(n1031), .Z(n1027) );
  CLKBUF_X1 U8276 ( .A(n1031), .Z(n1028) );
  CLKBUF_X1 U8277 ( .A(n1031), .Z(n1029) );
  CLKBUF_X1 U8278 ( .A(n1031), .Z(n1030) );
  NAND4_X1 U8279 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n7404)
         );
  NOR4_X1 U8280 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049)
         );
  OAI221_X1 U8281 ( .B1(n3110), .B2(n1054), .C1(n3143), .C2(n1055), .A(n1056), 
        .ZN(n1053) );
  AOI22_X1 U8282 ( .A1(n1057), .A2(n89), .B1(n1058), .B2(n341), .ZN(n1056) );
  OAI221_X1 U8283 ( .B1(n3225), .B2(n1059), .C1(n3176), .C2(n1060), .A(n1061), 
        .ZN(n1052) );
  AOI22_X1 U8284 ( .A1(n1062), .A2(n105), .B1(n1063), .B2(n325), .ZN(n1061) );
  OAI221_X1 U8285 ( .B1(n1064), .B2(n413), .C1(n3201), .C2(n1065), .A(n1066), 
        .ZN(n1051) );
  AOI22_X1 U8286 ( .A1(n1067), .A2(n73), .B1(n1068), .B2(n309), .ZN(n1066) );
  OAI221_X1 U8287 ( .B1(n1069), .B2(n205), .C1(n1070), .C2(n457), .A(n1071), 
        .ZN(n1050) );
  AOI222_X1 U8288 ( .A1(n2901), .A2(n1072), .B1(n1073), .B2(n161), .C1(n1074), 
        .C2(n397), .ZN(n1071) );
  NOR4_X1 U8289 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1048)
         );
  OAI22_X1 U8290 ( .A1(n3484), .A2(n1079), .B1(n3377), .B2(n1080), .ZN(n1078)
         );
  OAI22_X1 U8291 ( .A1(n3361), .A2(n1081), .B1(n3313), .B2(n1082), .ZN(n1077)
         );
  OAI22_X1 U8292 ( .A1(n3337), .A2(n1083), .B1(n3297), .B2(n1084), .ZN(n1076)
         );
  OAI22_X1 U8293 ( .A1(n3281), .A2(n1085), .B1(n3249), .B2(n1086), .ZN(n1075)
         );
  AOI221_X1 U8294 ( .B1(n1087), .B2(n237), .C1(n1088), .C2(n1), .A(n1089), 
        .ZN(n1047) );
  OAI22_X1 U8295 ( .A1(n3418), .A2(n1090), .B1(n3517), .B2(n1091), .ZN(n1089)
         );
  AOI211_X1 U8296 ( .C1(n1092), .C2(n221), .A(n1093), .B(n1094), .ZN(n1046) );
  OAI22_X1 U8297 ( .A1(n3443), .A2(n1095), .B1(n3393), .B2(n1096), .ZN(n1093)
         );
  NAND4_X1 U8298 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n7403)
         );
  NOR4_X1 U8299 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100)
         );
  OAI221_X1 U8300 ( .B1(n3111), .B2(n1054), .C1(n3144), .C2(n1055), .A(n1105), 
        .ZN(n1104) );
  AOI22_X1 U8301 ( .A1(n1057), .A2(n90), .B1(n1058), .B2(n342), .ZN(n1105) );
  OAI221_X1 U8302 ( .B1(n3226), .B2(n1059), .C1(n3177), .C2(n1060), .A(n1106), 
        .ZN(n1103) );
  AOI22_X1 U8303 ( .A1(n1062), .A2(n106), .B1(n1063), .B2(n326), .ZN(n1106) );
  OAI221_X1 U8304 ( .B1(n1064), .B2(n414), .C1(n3202), .C2(n1065), .A(n1107), 
        .ZN(n1102) );
  AOI22_X1 U8305 ( .A1(n1067), .A2(n74), .B1(n1068), .B2(n310), .ZN(n1107) );
  OAI221_X1 U8306 ( .B1(n1069), .B2(n206), .C1(n1070), .C2(n458), .A(n1108), 
        .ZN(n1101) );
  AOI222_X1 U8307 ( .A1(n2902), .A2(n1072), .B1(n1073), .B2(n162), .C1(n1074), 
        .C2(n398), .ZN(n1108) );
  NOR4_X1 U8308 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1099)
         );
  OAI22_X1 U8309 ( .A1(n3485), .A2(n1079), .B1(n3378), .B2(n1080), .ZN(n1112)
         );
  OAI22_X1 U8310 ( .A1(n3362), .A2(n1081), .B1(n3314), .B2(n1082), .ZN(n1111)
         );
  OAI22_X1 U8311 ( .A1(n3338), .A2(n1083), .B1(n3298), .B2(n1084), .ZN(n1110)
         );
  OAI22_X1 U8312 ( .A1(n3282), .A2(n1085), .B1(n3250), .B2(n1086), .ZN(n1109)
         );
  AOI221_X1 U8313 ( .B1(n1087), .B2(n238), .C1(n1088), .C2(n2), .A(n1113), 
        .ZN(n1098) );
  OAI22_X1 U8314 ( .A1(n3419), .A2(n1090), .B1(n3518), .B2(n1091), .ZN(n1113)
         );
  AOI211_X1 U8315 ( .C1(n1092), .C2(n222), .A(n1114), .B(n1094), .ZN(n1097) );
  OAI22_X1 U8316 ( .A1(n3444), .A2(n1095), .B1(n3394), .B2(n1096), .ZN(n1114)
         );
  NAND4_X1 U8317 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n7402)
         );
  NOR4_X1 U8318 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118)
         );
  OAI221_X1 U8319 ( .B1(n3112), .B2(n1054), .C1(n3145), .C2(n1055), .A(n1123), 
        .ZN(n1122) );
  AOI22_X1 U8320 ( .A1(n1057), .A2(n91), .B1(n1058), .B2(n343), .ZN(n1123) );
  OAI221_X1 U8321 ( .B1(n3227), .B2(n1059), .C1(n3178), .C2(n1060), .A(n1124), 
        .ZN(n1121) );
  AOI22_X1 U8322 ( .A1(n1062), .A2(n107), .B1(n1063), .B2(n327), .ZN(n1124) );
  OAI221_X1 U8323 ( .B1(n1064), .B2(n415), .C1(n3203), .C2(n1065), .A(n1125), 
        .ZN(n1120) );
  AOI22_X1 U8324 ( .A1(n1067), .A2(n75), .B1(n1068), .B2(n311), .ZN(n1125) );
  OAI221_X1 U8325 ( .B1(n1069), .B2(n207), .C1(n1070), .C2(n459), .A(n1126), 
        .ZN(n1119) );
  AOI222_X1 U8326 ( .A1(n2903), .A2(n1072), .B1(n1073), .B2(n163), .C1(n1074), 
        .C2(n399), .ZN(n1126) );
  NOR4_X1 U8327 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1117)
         );
  OAI22_X1 U8328 ( .A1(n3486), .A2(n1079), .B1(n3379), .B2(n1080), .ZN(n1130)
         );
  OAI22_X1 U8329 ( .A1(n3363), .A2(n1081), .B1(n3315), .B2(n1082), .ZN(n1129)
         );
  OAI22_X1 U8330 ( .A1(n3339), .A2(n1083), .B1(n3299), .B2(n1084), .ZN(n1128)
         );
  OAI22_X1 U8331 ( .A1(n3283), .A2(n1085), .B1(n3251), .B2(n1086), .ZN(n1127)
         );
  AOI221_X1 U8332 ( .B1(n1087), .B2(n239), .C1(n1088), .C2(n3), .A(n1131), 
        .ZN(n1116) );
  OAI22_X1 U8333 ( .A1(n3420), .A2(n1090), .B1(n3519), .B2(n1091), .ZN(n1131)
         );
  AOI211_X1 U8334 ( .C1(n1092), .C2(n223), .A(n1132), .B(n1094), .ZN(n1115) );
  OAI22_X1 U8335 ( .A1(n3445), .A2(n1095), .B1(n3395), .B2(n1096), .ZN(n1132)
         );
  NAND4_X1 U8336 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n7401)
         );
  NOR4_X1 U8337 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136)
         );
  OAI221_X1 U8338 ( .B1(n3113), .B2(n1054), .C1(n3146), .C2(n1055), .A(n1141), 
        .ZN(n1140) );
  AOI22_X1 U8339 ( .A1(n1057), .A2(n92), .B1(n1058), .B2(n344), .ZN(n1141) );
  OAI221_X1 U8340 ( .B1(n3228), .B2(n1059), .C1(n3179), .C2(n1060), .A(n1142), 
        .ZN(n1139) );
  AOI22_X1 U8341 ( .A1(n1062), .A2(n108), .B1(n1063), .B2(n328), .ZN(n1142) );
  OAI221_X1 U8342 ( .B1(n1064), .B2(n416), .C1(n3204), .C2(n1065), .A(n1143), 
        .ZN(n1138) );
  AOI22_X1 U8343 ( .A1(n1067), .A2(n76), .B1(n1068), .B2(n312), .ZN(n1143) );
  OAI221_X1 U8344 ( .B1(n1069), .B2(n208), .C1(n1070), .C2(n460), .A(n1144), 
        .ZN(n1137) );
  AOI222_X1 U8345 ( .A1(n2904), .A2(n1072), .B1(n1073), .B2(n164), .C1(n1074), 
        .C2(n400), .ZN(n1144) );
  NOR4_X1 U8346 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1135)
         );
  OAI22_X1 U8347 ( .A1(n3487), .A2(n1079), .B1(n3380), .B2(n1080), .ZN(n1148)
         );
  OAI22_X1 U8348 ( .A1(n3364), .A2(n1081), .B1(n3316), .B2(n1082), .ZN(n1147)
         );
  OAI22_X1 U8349 ( .A1(n3340), .A2(n1083), .B1(n3300), .B2(n1084), .ZN(n1146)
         );
  OAI22_X1 U8350 ( .A1(n3284), .A2(n1085), .B1(n3252), .B2(n1086), .ZN(n1145)
         );
  AOI221_X1 U8351 ( .B1(n1087), .B2(n240), .C1(n1088), .C2(n4), .A(n1149), 
        .ZN(n1134) );
  OAI22_X1 U8352 ( .A1(n3421), .A2(n1090), .B1(n3520), .B2(n1091), .ZN(n1149)
         );
  AOI211_X1 U8353 ( .C1(n1092), .C2(n224), .A(n1150), .B(n1094), .ZN(n1133) );
  OAI22_X1 U8354 ( .A1(n3446), .A2(n1095), .B1(n3396), .B2(n1096), .ZN(n1150)
         );
  NAND4_X1 U8355 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n7400)
         );
  NOR4_X1 U8356 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154)
         );
  OAI221_X1 U8357 ( .B1(n3114), .B2(n1054), .C1(n3147), .C2(n1055), .A(n1159), 
        .ZN(n1158) );
  AOI22_X1 U8358 ( .A1(n1057), .A2(n93), .B1(n1058), .B2(n345), .ZN(n1159) );
  OAI221_X1 U8359 ( .B1(n3229), .B2(n1059), .C1(n3180), .C2(n1060), .A(n1160), 
        .ZN(n1157) );
  AOI22_X1 U8360 ( .A1(n1062), .A2(n109), .B1(n1063), .B2(n329), .ZN(n1160) );
  OAI221_X1 U8361 ( .B1(n1064), .B2(n417), .C1(n3205), .C2(n1065), .A(n1161), 
        .ZN(n1156) );
  AOI22_X1 U8362 ( .A1(n1067), .A2(n77), .B1(n1068), .B2(n313), .ZN(n1161) );
  OAI221_X1 U8363 ( .B1(n1069), .B2(n209), .C1(n1070), .C2(n461), .A(n1162), 
        .ZN(n1155) );
  AOI222_X1 U8364 ( .A1(n2905), .A2(n1072), .B1(n1073), .B2(n165), .C1(n1074), 
        .C2(n401), .ZN(n1162) );
  NOR4_X1 U8365 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1153)
         );
  OAI22_X1 U8366 ( .A1(n3488), .A2(n1079), .B1(n3381), .B2(n1080), .ZN(n1166)
         );
  OAI22_X1 U8367 ( .A1(n3365), .A2(n1081), .B1(n3317), .B2(n1082), .ZN(n1165)
         );
  OAI22_X1 U8368 ( .A1(n3341), .A2(n1083), .B1(n3301), .B2(n1084), .ZN(n1164)
         );
  OAI22_X1 U8369 ( .A1(n3285), .A2(n1085), .B1(n3253), .B2(n1086), .ZN(n1163)
         );
  AOI221_X1 U8370 ( .B1(n1087), .B2(n241), .C1(n1088), .C2(n5), .A(n1167), 
        .ZN(n1152) );
  OAI22_X1 U8371 ( .A1(n3422), .A2(n1090), .B1(n3521), .B2(n1091), .ZN(n1167)
         );
  AOI211_X1 U8372 ( .C1(n1092), .C2(n225), .A(n1168), .B(n1094), .ZN(n1151) );
  OAI22_X1 U8373 ( .A1(n3447), .A2(n1095), .B1(n3397), .B2(n1096), .ZN(n1168)
         );
  NAND4_X1 U8374 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n7399)
         );
  NOR4_X1 U8375 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172)
         );
  OAI221_X1 U8376 ( .B1(n3115), .B2(n1054), .C1(n3148), .C2(n1055), .A(n1177), 
        .ZN(n1176) );
  AOI22_X1 U8377 ( .A1(n1057), .A2(n94), .B1(n1058), .B2(n346), .ZN(n1177) );
  OAI221_X1 U8378 ( .B1(n3230), .B2(n1059), .C1(n3181), .C2(n1060), .A(n1178), 
        .ZN(n1175) );
  AOI22_X1 U8379 ( .A1(n1062), .A2(n110), .B1(n1063), .B2(n330), .ZN(n1178) );
  OAI221_X1 U8380 ( .B1(n1064), .B2(n418), .C1(n3206), .C2(n1065), .A(n1179), 
        .ZN(n1174) );
  AOI22_X1 U8381 ( .A1(n1067), .A2(n78), .B1(n1068), .B2(n314), .ZN(n1179) );
  OAI221_X1 U8382 ( .B1(n1069), .B2(n210), .C1(n1070), .C2(n462), .A(n1180), 
        .ZN(n1173) );
  AOI222_X1 U8383 ( .A1(n2906), .A2(n1072), .B1(n1073), .B2(n166), .C1(n1074), 
        .C2(n402), .ZN(n1180) );
  NOR4_X1 U8384 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1171)
         );
  OAI22_X1 U8385 ( .A1(n3489), .A2(n1079), .B1(n3382), .B2(n1080), .ZN(n1184)
         );
  OAI22_X1 U8386 ( .A1(n3366), .A2(n1081), .B1(n3318), .B2(n1082), .ZN(n1183)
         );
  OAI22_X1 U8387 ( .A1(n3342), .A2(n1083), .B1(n3302), .B2(n1084), .ZN(n1182)
         );
  OAI22_X1 U8388 ( .A1(n3286), .A2(n1085), .B1(n3254), .B2(n1086), .ZN(n1181)
         );
  AOI221_X1 U8389 ( .B1(n1087), .B2(n242), .C1(n1088), .C2(n6), .A(n1185), 
        .ZN(n1170) );
  OAI22_X1 U8390 ( .A1(n3423), .A2(n1090), .B1(n3522), .B2(n1091), .ZN(n1185)
         );
  AOI211_X1 U8391 ( .C1(n1092), .C2(n226), .A(n1186), .B(n1094), .ZN(n1169) );
  OAI22_X1 U8392 ( .A1(n3448), .A2(n1095), .B1(n3398), .B2(n1096), .ZN(n1186)
         );
  NAND4_X1 U8393 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n2214), .ZN(n7398)
         );
  NOR4_X1 U8394 ( .A1(n2215), .A2(n2216), .A3(n2217), .A4(n2218), .ZN(n2214)
         );
  OAI221_X1 U8395 ( .B1(n3116), .B2(n1054), .C1(n3149), .C2(n1055), .A(n2219), 
        .ZN(n2218) );
  AOI22_X1 U8396 ( .A1(n1057), .A2(n95), .B1(n1058), .B2(n347), .ZN(n2219) );
  OAI221_X1 U8397 ( .B1(n3231), .B2(n1059), .C1(n3182), .C2(n1060), .A(n2220), 
        .ZN(n2217) );
  AOI22_X1 U8398 ( .A1(n1062), .A2(n111), .B1(n1063), .B2(n331), .ZN(n2220) );
  OAI221_X1 U8399 ( .B1(n1064), .B2(n419), .C1(n3207), .C2(n1065), .A(n2221), 
        .ZN(n2216) );
  AOI22_X1 U8400 ( .A1(n1067), .A2(n79), .B1(n1068), .B2(n315), .ZN(n2221) );
  OAI221_X1 U8401 ( .B1(n1069), .B2(n211), .C1(n1070), .C2(n463), .A(n2222), 
        .ZN(n2215) );
  AOI222_X1 U8402 ( .A1(n2907), .A2(n1072), .B1(n1073), .B2(n167), .C1(n1074), 
        .C2(n403), .ZN(n2222) );
  NOR4_X1 U8403 ( .A1(n2223), .A2(n2224), .A3(n2225), .A4(n2226), .ZN(n1189)
         );
  OAI22_X1 U8404 ( .A1(n3490), .A2(n1079), .B1(n3383), .B2(n1080), .ZN(n2226)
         );
  OAI22_X1 U8405 ( .A1(n3367), .A2(n1081), .B1(n3319), .B2(n1082), .ZN(n2225)
         );
  OAI22_X1 U8406 ( .A1(n3343), .A2(n1083), .B1(n3303), .B2(n1084), .ZN(n2224)
         );
  OAI22_X1 U8407 ( .A1(n3287), .A2(n1085), .B1(n3255), .B2(n1086), .ZN(n2223)
         );
  AOI221_X1 U8408 ( .B1(n1087), .B2(n243), .C1(n1088), .C2(n7), .A(n2227), 
        .ZN(n1188) );
  OAI22_X1 U8409 ( .A1(n3424), .A2(n1090), .B1(n3523), .B2(n1091), .ZN(n2227)
         );
  AOI211_X1 U8410 ( .C1(n1092), .C2(n227), .A(n2228), .B(n1094), .ZN(n1187) );
  OAI22_X1 U8411 ( .A1(n3449), .A2(n1095), .B1(n3399), .B2(n1096), .ZN(n2228)
         );
  NAND4_X1 U8412 ( .A1(n2229), .A2(n2230), .A3(n2231), .A4(n2232), .ZN(n7397)
         );
  NOR4_X1 U8413 ( .A1(n2233), .A2(n2234), .A3(n2235), .A4(n2236), .ZN(n2232)
         );
  OAI221_X1 U8414 ( .B1(n3117), .B2(n1054), .C1(n3150), .C2(n1055), .A(n2237), 
        .ZN(n2236) );
  AOI22_X1 U8415 ( .A1(n1057), .A2(n96), .B1(n1058), .B2(n348), .ZN(n2237) );
  OAI221_X1 U8416 ( .B1(n3232), .B2(n1059), .C1(n3183), .C2(n1060), .A(n2238), 
        .ZN(n2235) );
  AOI22_X1 U8417 ( .A1(n1062), .A2(n112), .B1(n1063), .B2(n332), .ZN(n2238) );
  OAI221_X1 U8418 ( .B1(n1064), .B2(n420), .C1(n3208), .C2(n1065), .A(n2239), 
        .ZN(n2234) );
  AOI22_X1 U8419 ( .A1(n1067), .A2(n80), .B1(n1068), .B2(n316), .ZN(n2239) );
  OAI221_X1 U8420 ( .B1(n1069), .B2(n212), .C1(n1070), .C2(n464), .A(n2240), 
        .ZN(n2233) );
  AOI222_X1 U8421 ( .A1(n2908), .A2(n1072), .B1(n1073), .B2(n168), .C1(n1074), 
        .C2(n404), .ZN(n2240) );
  NOR4_X1 U8422 ( .A1(n2241), .A2(n2242), .A3(n2243), .A4(n2244), .ZN(n2231)
         );
  OAI22_X1 U8423 ( .A1(n3491), .A2(n1079), .B1(n3384), .B2(n1080), .ZN(n2244)
         );
  OAI22_X1 U8424 ( .A1(n3368), .A2(n1081), .B1(n3320), .B2(n1082), .ZN(n2243)
         );
  OAI22_X1 U8425 ( .A1(n3344), .A2(n1083), .B1(n3304), .B2(n1084), .ZN(n2242)
         );
  OAI22_X1 U8426 ( .A1(n3288), .A2(n1085), .B1(n3256), .B2(n1086), .ZN(n2241)
         );
  AOI221_X1 U8427 ( .B1(n1087), .B2(n244), .C1(n1088), .C2(n8), .A(n2245), 
        .ZN(n2230) );
  OAI22_X1 U8428 ( .A1(n3425), .A2(n1090), .B1(n3524), .B2(n1091), .ZN(n2245)
         );
  AOI211_X1 U8429 ( .C1(n1092), .C2(n228), .A(n2246), .B(n1094), .ZN(n2229) );
  OAI22_X1 U8430 ( .A1(n3450), .A2(n1095), .B1(n3400), .B2(n1096), .ZN(n2246)
         );
  NAND4_X1 U8431 ( .A1(n2247), .A2(n2248), .A3(n2249), .A4(n2250), .ZN(n7396)
         );
  NOR4_X1 U8432 ( .A1(n2251), .A2(n2252), .A3(n2253), .A4(n2254), .ZN(n2250)
         );
  OAI221_X1 U8433 ( .B1(n3118), .B2(n1054), .C1(n3151), .C2(n1055), .A(n2255), 
        .ZN(n2254) );
  AOI22_X1 U8434 ( .A1(n1057), .A2(n97), .B1(n1058), .B2(n349), .ZN(n2255) );
  OAI221_X1 U8435 ( .B1(n3233), .B2(n1059), .C1(n3184), .C2(n1060), .A(n2256), 
        .ZN(n2253) );
  AOI22_X1 U8436 ( .A1(n1062), .A2(n113), .B1(n1063), .B2(n333), .ZN(n2256) );
  OAI221_X1 U8437 ( .B1(n1064), .B2(n421), .C1(n3209), .C2(n1065), .A(n2257), 
        .ZN(n2252) );
  AOI22_X1 U8438 ( .A1(n1067), .A2(n81), .B1(n1068), .B2(n317), .ZN(n2257) );
  OAI221_X1 U8439 ( .B1(n1069), .B2(n213), .C1(n1070), .C2(n465), .A(n2258), 
        .ZN(n2251) );
  AOI222_X1 U8440 ( .A1(n2909), .A2(n1072), .B1(n1073), .B2(n169), .C1(n1074), 
        .C2(n405), .ZN(n2258) );
  NOR4_X1 U8441 ( .A1(n2259), .A2(n2260), .A3(n2261), .A4(n2262), .ZN(n2249)
         );
  OAI22_X1 U8442 ( .A1(n3492), .A2(n1079), .B1(n3385), .B2(n1080), .ZN(n2262)
         );
  OAI22_X1 U8443 ( .A1(n3369), .A2(n1081), .B1(n3321), .B2(n1082), .ZN(n2261)
         );
  OAI22_X1 U8444 ( .A1(n3345), .A2(n1083), .B1(n3305), .B2(n1084), .ZN(n2260)
         );
  OAI22_X1 U8445 ( .A1(n3289), .A2(n1085), .B1(n3257), .B2(n1086), .ZN(n2259)
         );
  AOI221_X1 U8446 ( .B1(n1087), .B2(n245), .C1(n1088), .C2(n9), .A(n2263), 
        .ZN(n2248) );
  OAI22_X1 U8447 ( .A1(n3426), .A2(n1090), .B1(n3525), .B2(n1091), .ZN(n2263)
         );
  AOI211_X1 U8448 ( .C1(n1092), .C2(n229), .A(n2264), .B(n1094), .ZN(n2247) );
  OAI22_X1 U8449 ( .A1(n3451), .A2(n1095), .B1(n3401), .B2(n1096), .ZN(n2264)
         );
  NAND4_X1 U8450 ( .A1(n2265), .A2(n2266), .A3(n2267), .A4(n2268), .ZN(n7395)
         );
  NOR4_X1 U8451 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2268)
         );
  OAI221_X1 U8452 ( .B1(n3119), .B2(n1054), .C1(n3152), .C2(n1055), .A(n2273), 
        .ZN(n2272) );
  AOI22_X1 U8453 ( .A1(n1057), .A2(n98), .B1(n1058), .B2(n350), .ZN(n2273) );
  OAI221_X1 U8454 ( .B1(n3234), .B2(n1059), .C1(n3185), .C2(n1060), .A(n2274), 
        .ZN(n2271) );
  AOI22_X1 U8455 ( .A1(n1062), .A2(n114), .B1(n1063), .B2(n334), .ZN(n2274) );
  OAI221_X1 U8456 ( .B1(n1064), .B2(n422), .C1(n3210), .C2(n1065), .A(n2275), 
        .ZN(n2270) );
  AOI22_X1 U8457 ( .A1(n1067), .A2(n82), .B1(n1068), .B2(n318), .ZN(n2275) );
  OAI221_X1 U8458 ( .B1(n1069), .B2(n214), .C1(n1070), .C2(n466), .A(n2276), 
        .ZN(n2269) );
  AOI222_X1 U8459 ( .A1(n2910), .A2(n1072), .B1(n1073), .B2(n170), .C1(n1074), 
        .C2(n406), .ZN(n2276) );
  NOR4_X1 U8460 ( .A1(n2277), .A2(n2278), .A3(n2279), .A4(n2280), .ZN(n2267)
         );
  OAI22_X1 U8461 ( .A1(n3493), .A2(n1079), .B1(n3386), .B2(n1080), .ZN(n2280)
         );
  OAI22_X1 U8462 ( .A1(n3370), .A2(n1081), .B1(n3322), .B2(n1082), .ZN(n2279)
         );
  OAI22_X1 U8463 ( .A1(n3346), .A2(n1083), .B1(n3306), .B2(n1084), .ZN(n2278)
         );
  OAI22_X1 U8464 ( .A1(n3290), .A2(n1085), .B1(n3258), .B2(n1086), .ZN(n2277)
         );
  AOI221_X1 U8465 ( .B1(n1087), .B2(n246), .C1(n1088), .C2(n10), .A(n2281), 
        .ZN(n2266) );
  OAI22_X1 U8466 ( .A1(n3427), .A2(n1090), .B1(n3526), .B2(n1091), .ZN(n2281)
         );
  AOI211_X1 U8467 ( .C1(n1092), .C2(n230), .A(n2282), .B(n1094), .ZN(n2265) );
  OAI22_X1 U8468 ( .A1(n3452), .A2(n1095), .B1(n3402), .B2(n1096), .ZN(n2282)
         );
  NAND4_X1 U8469 ( .A1(n2283), .A2(n2284), .A3(n2285), .A4(n2286), .ZN(n7394)
         );
  NOR4_X1 U8470 ( .A1(n2287), .A2(n2288), .A3(n2289), .A4(n2290), .ZN(n2286)
         );
  OAI221_X1 U8471 ( .B1(n3120), .B2(n1054), .C1(n3153), .C2(n1055), .A(n2291), 
        .ZN(n2290) );
  AOI22_X1 U8472 ( .A1(n1057), .A2(n99), .B1(n1058), .B2(n351), .ZN(n2291) );
  OAI221_X1 U8473 ( .B1(n3235), .B2(n1059), .C1(n3186), .C2(n1060), .A(n2292), 
        .ZN(n2289) );
  AOI22_X1 U8474 ( .A1(n1062), .A2(n115), .B1(n1063), .B2(n335), .ZN(n2292) );
  OAI221_X1 U8475 ( .B1(n1064), .B2(n423), .C1(n3211), .C2(n1065), .A(n2293), 
        .ZN(n2288) );
  AOI22_X1 U8476 ( .A1(n1067), .A2(n83), .B1(n1068), .B2(n319), .ZN(n2293) );
  OAI221_X1 U8477 ( .B1(n1069), .B2(n215), .C1(n1070), .C2(n467), .A(n2294), 
        .ZN(n2287) );
  AOI222_X1 U8478 ( .A1(n2911), .A2(n1072), .B1(n1073), .B2(n171), .C1(n1074), 
        .C2(n407), .ZN(n2294) );
  NOR4_X1 U8479 ( .A1(n2295), .A2(n2296), .A3(n2297), .A4(n2298), .ZN(n2285)
         );
  OAI22_X1 U8480 ( .A1(n3494), .A2(n1079), .B1(n3387), .B2(n1080), .ZN(n2298)
         );
  OAI22_X1 U8481 ( .A1(n3371), .A2(n1081), .B1(n3323), .B2(n1082), .ZN(n2297)
         );
  OAI22_X1 U8482 ( .A1(n3347), .A2(n1083), .B1(n3307), .B2(n1084), .ZN(n2296)
         );
  OAI22_X1 U8483 ( .A1(n3291), .A2(n1085), .B1(n3259), .B2(n1086), .ZN(n2295)
         );
  AOI221_X1 U8484 ( .B1(n1087), .B2(n247), .C1(n1088), .C2(n11), .A(n2299), 
        .ZN(n2284) );
  OAI22_X1 U8485 ( .A1(n3428), .A2(n1090), .B1(n3527), .B2(n1091), .ZN(n2299)
         );
  AOI211_X1 U8486 ( .C1(n1092), .C2(n231), .A(n2300), .B(n1094), .ZN(n2283) );
  OAI22_X1 U8487 ( .A1(n3453), .A2(n1095), .B1(n3403), .B2(n1096), .ZN(n2300)
         );
  NAND4_X1 U8488 ( .A1(n2301), .A2(n2302), .A3(n2303), .A4(n2304), .ZN(n7393)
         );
  NOR4_X1 U8489 ( .A1(n2305), .A2(n2306), .A3(n2307), .A4(n2308), .ZN(n2304)
         );
  OAI221_X1 U8490 ( .B1(n3121), .B2(n1054), .C1(n3154), .C2(n1055), .A(n2309), 
        .ZN(n2308) );
  AOI22_X1 U8491 ( .A1(n1057), .A2(n100), .B1(n1058), .B2(n352), .ZN(n2309) );
  OAI221_X1 U8492 ( .B1(n3236), .B2(n1059), .C1(n3187), .C2(n1060), .A(n2310), 
        .ZN(n2307) );
  AOI22_X1 U8493 ( .A1(n1062), .A2(n116), .B1(n1063), .B2(n336), .ZN(n2310) );
  OAI221_X1 U8494 ( .B1(n1064), .B2(n424), .C1(n3212), .C2(n1065), .A(n2311), 
        .ZN(n2306) );
  AOI22_X1 U8495 ( .A1(n1067), .A2(n84), .B1(n1068), .B2(n320), .ZN(n2311) );
  OAI221_X1 U8496 ( .B1(n1069), .B2(n216), .C1(n1070), .C2(n468), .A(n2312), 
        .ZN(n2305) );
  AOI222_X1 U8497 ( .A1(n2912), .A2(n1072), .B1(n1073), .B2(n172), .C1(n1074), 
        .C2(n408), .ZN(n2312) );
  NOR4_X1 U8498 ( .A1(n2313), .A2(n2314), .A3(n2315), .A4(n2316), .ZN(n2303)
         );
  OAI22_X1 U8499 ( .A1(n3495), .A2(n1079), .B1(n3388), .B2(n1080), .ZN(n2316)
         );
  OAI22_X1 U8500 ( .A1(n3372), .A2(n1081), .B1(n3324), .B2(n1082), .ZN(n2315)
         );
  OAI22_X1 U8501 ( .A1(n3348), .A2(n1083), .B1(n3308), .B2(n1084), .ZN(n2314)
         );
  OAI22_X1 U8502 ( .A1(n3292), .A2(n1085), .B1(n3260), .B2(n1086), .ZN(n2313)
         );
  AOI221_X1 U8503 ( .B1(n1087), .B2(n248), .C1(n1088), .C2(n12), .A(n2317), 
        .ZN(n2302) );
  OAI22_X1 U8504 ( .A1(n3429), .A2(n1090), .B1(n3528), .B2(n1091), .ZN(n2317)
         );
  AOI211_X1 U8505 ( .C1(n1092), .C2(n232), .A(n2318), .B(n1094), .ZN(n2301) );
  OAI22_X1 U8506 ( .A1(n3454), .A2(n1095), .B1(n3404), .B2(n1096), .ZN(n2318)
         );
  NAND4_X1 U8507 ( .A1(n2319), .A2(n2320), .A3(n2321), .A4(n2322), .ZN(n7392)
         );
  NOR4_X1 U8508 ( .A1(n2323), .A2(n2324), .A3(n2325), .A4(n2326), .ZN(n2322)
         );
  OAI221_X1 U8509 ( .B1(n3122), .B2(n1054), .C1(n3155), .C2(n1055), .A(n2327), 
        .ZN(n2326) );
  AOI22_X1 U8510 ( .A1(n1057), .A2(n101), .B1(n1058), .B2(n353), .ZN(n2327) );
  OAI221_X1 U8511 ( .B1(n3237), .B2(n1059), .C1(n3188), .C2(n1060), .A(n2328), 
        .ZN(n2325) );
  AOI22_X1 U8512 ( .A1(n1062), .A2(n117), .B1(n1063), .B2(n337), .ZN(n2328) );
  OAI221_X1 U8513 ( .B1(n1064), .B2(n425), .C1(n3213), .C2(n1065), .A(n2329), 
        .ZN(n2324) );
  AOI22_X1 U8514 ( .A1(n1067), .A2(n85), .B1(n1068), .B2(n321), .ZN(n2329) );
  OAI221_X1 U8515 ( .B1(n1069), .B2(n217), .C1(n1070), .C2(n469), .A(n2330), 
        .ZN(n2323) );
  AOI222_X1 U8516 ( .A1(n2913), .A2(n1072), .B1(n1073), .B2(n173), .C1(n1074), 
        .C2(n409), .ZN(n2330) );
  NOR4_X1 U8517 ( .A1(n2331), .A2(n2332), .A3(n2333), .A4(n2334), .ZN(n2321)
         );
  OAI22_X1 U8518 ( .A1(n3496), .A2(n1079), .B1(n3389), .B2(n1080), .ZN(n2334)
         );
  OAI22_X1 U8519 ( .A1(n3373), .A2(n1081), .B1(n3325), .B2(n1082), .ZN(n2333)
         );
  OAI22_X1 U8520 ( .A1(n3349), .A2(n1083), .B1(n3309), .B2(n1084), .ZN(n2332)
         );
  OAI22_X1 U8521 ( .A1(n3293), .A2(n1085), .B1(n3261), .B2(n1086), .ZN(n2331)
         );
  AOI221_X1 U8522 ( .B1(n1087), .B2(n249), .C1(n1088), .C2(n13), .A(n2335), 
        .ZN(n2320) );
  OAI22_X1 U8523 ( .A1(n3430), .A2(n1090), .B1(n3529), .B2(n1091), .ZN(n2335)
         );
  AOI211_X1 U8524 ( .C1(n1092), .C2(n233), .A(n2336), .B(n1094), .ZN(n2319) );
  OAI22_X1 U8525 ( .A1(n3455), .A2(n1095), .B1(n3405), .B2(n1096), .ZN(n2336)
         );
  NAND4_X1 U8526 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n7391)
         );
  NOR4_X1 U8527 ( .A1(n2341), .A2(n2342), .A3(n2343), .A4(n2344), .ZN(n2340)
         );
  OAI221_X1 U8528 ( .B1(n3123), .B2(n1054), .C1(n3156), .C2(n1055), .A(n2345), 
        .ZN(n2344) );
  AOI22_X1 U8529 ( .A1(n1057), .A2(n102), .B1(n1058), .B2(n354), .ZN(n2345) );
  OAI221_X1 U8530 ( .B1(n3238), .B2(n1059), .C1(n3189), .C2(n1060), .A(n2346), 
        .ZN(n2343) );
  AOI22_X1 U8531 ( .A1(n1062), .A2(n118), .B1(n1063), .B2(n338), .ZN(n2346) );
  OAI221_X1 U8532 ( .B1(n1064), .B2(n426), .C1(n3214), .C2(n1065), .A(n2347), 
        .ZN(n2342) );
  AOI22_X1 U8533 ( .A1(n1067), .A2(n86), .B1(n1068), .B2(n322), .ZN(n2347) );
  OAI221_X1 U8534 ( .B1(n1069), .B2(n218), .C1(n1070), .C2(n470), .A(n2348), 
        .ZN(n2341) );
  AOI222_X1 U8535 ( .A1(n2914), .A2(n1072), .B1(n1073), .B2(n174), .C1(n1074), 
        .C2(n410), .ZN(n2348) );
  NOR4_X1 U8536 ( .A1(n2349), .A2(n2350), .A3(n2351), .A4(n2352), .ZN(n2339)
         );
  OAI22_X1 U8537 ( .A1(n3497), .A2(n1079), .B1(n3390), .B2(n1080), .ZN(n2352)
         );
  OAI22_X1 U8538 ( .A1(n3374), .A2(n1081), .B1(n3326), .B2(n1082), .ZN(n2351)
         );
  OAI22_X1 U8539 ( .A1(n3350), .A2(n1083), .B1(n3310), .B2(n1084), .ZN(n2350)
         );
  OAI22_X1 U8540 ( .A1(n3294), .A2(n1085), .B1(n3262), .B2(n1086), .ZN(n2349)
         );
  AOI221_X1 U8541 ( .B1(n1087), .B2(n250), .C1(n1088), .C2(n14), .A(n2353), 
        .ZN(n2338) );
  OAI22_X1 U8542 ( .A1(n3431), .A2(n1090), .B1(n3530), .B2(n1091), .ZN(n2353)
         );
  AOI211_X1 U8543 ( .C1(n1092), .C2(n234), .A(n2354), .B(n1094), .ZN(n2337) );
  OAI22_X1 U8544 ( .A1(n3456), .A2(n1095), .B1(n3406), .B2(n1096), .ZN(n2354)
         );
  NAND4_X1 U8545 ( .A1(n2355), .A2(n2356), .A3(n2357), .A4(n2358), .ZN(n7390)
         );
  NOR4_X1 U8546 ( .A1(n2359), .A2(n2360), .A3(n2361), .A4(n2362), .ZN(n2358)
         );
  OAI221_X1 U8547 ( .B1(n3124), .B2(n1054), .C1(n3157), .C2(n1055), .A(n2363), 
        .ZN(n2362) );
  AOI22_X1 U8548 ( .A1(n1057), .A2(n103), .B1(n1058), .B2(n355), .ZN(n2363) );
  OAI221_X1 U8549 ( .B1(n3239), .B2(n1059), .C1(n3190), .C2(n1060), .A(n2364), 
        .ZN(n2361) );
  AOI22_X1 U8550 ( .A1(n1062), .A2(n119), .B1(n1063), .B2(n339), .ZN(n2364) );
  OAI221_X1 U8551 ( .B1(n1064), .B2(n427), .C1(n3215), .C2(n1065), .A(n2365), 
        .ZN(n2360) );
  AOI22_X1 U8552 ( .A1(n1067), .A2(n87), .B1(n1068), .B2(n323), .ZN(n2365) );
  OAI221_X1 U8553 ( .B1(n1069), .B2(n219), .C1(n1070), .C2(n471), .A(n2366), 
        .ZN(n2359) );
  AOI222_X1 U8554 ( .A1(n2915), .A2(n1072), .B1(n1073), .B2(n175), .C1(n1074), 
        .C2(n411), .ZN(n2366) );
  NOR4_X1 U8555 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(n2357)
         );
  OAI22_X1 U8556 ( .A1(n3498), .A2(n1079), .B1(n3391), .B2(n1080), .ZN(n2370)
         );
  OAI22_X1 U8557 ( .A1(n3375), .A2(n1081), .B1(n3327), .B2(n1082), .ZN(n2369)
         );
  OAI22_X1 U8558 ( .A1(n3351), .A2(n1083), .B1(n3311), .B2(n1084), .ZN(n2368)
         );
  OAI22_X1 U8559 ( .A1(n3295), .A2(n1085), .B1(n3263), .B2(n1086), .ZN(n2367)
         );
  AOI221_X1 U8560 ( .B1(n1087), .B2(n251), .C1(n1088), .C2(n15), .A(n2371), 
        .ZN(n2356) );
  OAI22_X1 U8561 ( .A1(n3432), .A2(n1090), .B1(n3531), .B2(n1091), .ZN(n2371)
         );
  AOI211_X1 U8562 ( .C1(n1092), .C2(n235), .A(n2372), .B(n1094), .ZN(n2355) );
  OAI22_X1 U8563 ( .A1(n3457), .A2(n1095), .B1(n3407), .B2(n1096), .ZN(n2372)
         );
  NAND4_X1 U8564 ( .A1(n2373), .A2(n2374), .A3(n2375), .A4(n2376), .ZN(n7389)
         );
  NOR4_X1 U8565 ( .A1(n2377), .A2(n2378), .A3(n2379), .A4(n2380), .ZN(n2376)
         );
  OAI221_X1 U8566 ( .B1(n3125), .B2(n1054), .C1(n3158), .C2(n1055), .A(n2381), 
        .ZN(n2380) );
  AOI22_X1 U8567 ( .A1(n1057), .A2(n104), .B1(n1058), .B2(n356), .ZN(n2381) );
  AND2_X1 U8568 ( .A1(n2382), .A2(n2383), .ZN(n1058) );
  AND2_X1 U8569 ( .A1(n2384), .A2(n2385), .ZN(n1057) );
  NAND2_X1 U8570 ( .A1(n2386), .A2(n2385), .ZN(n1055) );
  NAND2_X1 U8571 ( .A1(n2382), .A2(n2385), .ZN(n1054) );
  OAI221_X1 U8572 ( .B1(n3240), .B2(n1059), .C1(n3191), .C2(n1060), .A(n2387), 
        .ZN(n2379) );
  AOI22_X1 U8573 ( .A1(n1062), .A2(n120), .B1(n1063), .B2(n340), .ZN(n2387) );
  AND2_X1 U8574 ( .A1(n2388), .A2(n2385), .ZN(n1063) );
  AND2_X1 U8575 ( .A1(n2388), .A2(n2389), .ZN(n1062) );
  NAND2_X1 U8576 ( .A1(n2382), .A2(n2389), .ZN(n1060) );
  NAND2_X1 U8577 ( .A1(n2386), .A2(n2389), .ZN(n1059) );
  OAI221_X1 U8578 ( .B1(n1064), .B2(n428), .C1(n3216), .C2(n1065), .A(n2390), 
        .ZN(n2378) );
  AOI22_X1 U8579 ( .A1(n1067), .A2(n88), .B1(n1068), .B2(n324), .ZN(n2390) );
  AND2_X1 U8580 ( .A1(n2384), .A2(n2391), .ZN(n1068) );
  AND2_X1 U8581 ( .A1(n2388), .A2(n2391), .ZN(n1067) );
  NAND2_X1 U8582 ( .A1(n2384), .A2(n2389), .ZN(n1065) );
  NAND2_X1 U8583 ( .A1(n2386), .A2(n2391), .ZN(n1064) );
  OAI221_X1 U8584 ( .B1(n1069), .B2(n220), .C1(n1070), .C2(n472), .A(n2392), 
        .ZN(n2377) );
  AOI222_X1 U8585 ( .A1(n2916), .A2(n1072), .B1(n1073), .B2(n176), .C1(n1074), 
        .C2(n412), .ZN(n2392) );
  AND2_X1 U8586 ( .A1(n2382), .A2(n2391), .ZN(n1074) );
  AND2_X1 U8587 ( .A1(n2386), .A2(n2393), .ZN(n1073) );
  AND2_X1 U8588 ( .A1(n2384), .A2(n2393), .ZN(n1072) );
  NAND2_X1 U8589 ( .A1(n2388), .A2(n2393), .ZN(n1070) );
  NAND2_X1 U8590 ( .A1(n2382), .A2(n2393), .ZN(n1069) );
  NOR4_X1 U8591 ( .A1(n2394), .A2(n2395), .A3(n2396), .A4(n2397), .ZN(n2375)
         );
  OAI22_X1 U8592 ( .A1(n3499), .A2(n1079), .B1(n3392), .B2(n1080), .ZN(n2397)
         );
  NAND2_X1 U8593 ( .A1(n2386), .A2(n2398), .ZN(n1080) );
  NAND2_X1 U8594 ( .A1(n2382), .A2(n2399), .ZN(n1079) );
  OAI22_X1 U8595 ( .A1(n3376), .A2(n1081), .B1(n3328), .B2(n1082), .ZN(n2396)
         );
  NAND2_X1 U8596 ( .A1(n2388), .A2(n2398), .ZN(n1082) );
  NAND2_X1 U8597 ( .A1(n2384), .A2(n2398), .ZN(n1081) );
  OAI22_X1 U8598 ( .A1(n3352), .A2(n1083), .B1(n3312), .B2(n1084), .ZN(n2395)
         );
  NAND2_X1 U8599 ( .A1(n2386), .A2(n2383), .ZN(n1084) );
  NAND2_X1 U8600 ( .A1(n2382), .A2(n2398), .ZN(n1083) );
  OAI22_X1 U8601 ( .A1(n3296), .A2(n1085), .B1(n3264), .B2(n1086), .ZN(n2394)
         );
  NAND2_X1 U8602 ( .A1(n2388), .A2(n2383), .ZN(n1086) );
  NAND2_X1 U8603 ( .A1(n2384), .A2(n2383), .ZN(n1085) );
  AOI221_X1 U8604 ( .B1(n1087), .B2(n252), .C1(n1088), .C2(n16), .A(n2400), 
        .ZN(n2374) );
  OAI22_X1 U8605 ( .A1(n3433), .A2(n1090), .B1(n3532), .B2(n1091), .ZN(n2400)
         );
  NAND2_X1 U8606 ( .A1(n2386), .A2(n2399), .ZN(n1091) );
  NAND2_X1 U8607 ( .A1(n2382), .A2(n2401), .ZN(n1090) );
  AND2_X1 U8608 ( .A1(n2402), .A2(n2403), .ZN(n2382) );
  AND2_X1 U8609 ( .A1(n2384), .A2(n2399), .ZN(n1088) );
  AND2_X1 U8610 ( .A1(n2388), .A2(n2399), .ZN(n1087) );
  AOI211_X1 U8611 ( .C1(n1092), .C2(n236), .A(n2404), .B(n1094), .ZN(n2373) );
  INV_X1 U8612 ( .A(n2408), .ZN(n2406) );
  OAI22_X1 U8613 ( .A1(n3458), .A2(n1095), .B1(n3408), .B2(n1096), .ZN(n2404)
         );
  NAND2_X1 U8614 ( .A1(n2388), .A2(n2401), .ZN(n1096) );
  AND2_X1 U8615 ( .A1(n2402), .A2(n2409), .ZN(n2388) );
  NAND2_X1 U8616 ( .A1(n2384), .A2(n2401), .ZN(n1095) );
  AND2_X1 U8617 ( .A1(n2402), .A2(n2410), .ZN(n2384) );
  AND2_X1 U8618 ( .A1(n2386), .A2(n2401), .ZN(n1092) );
  AND2_X1 U8619 ( .A1(n2402), .A2(n2411), .ZN(n2386) );
  MUX2_X1 U8620 ( .A(n3039), .B(n2412), .S(n2413), .Z(n2213) );
  MUX2_X1 U8621 ( .A(n3040), .B(n2414), .S(n2413), .Z(n2212) );
  MUX2_X1 U8622 ( .A(n3041), .B(n2415), .S(n2413), .Z(n2211) );
  MUX2_X1 U8623 ( .A(n3042), .B(n2416), .S(n2413), .Z(n2210) );
  MUX2_X1 U8624 ( .A(n3043), .B(n2417), .S(n2413), .Z(n2209) );
  MUX2_X1 U8625 ( .A(n3044), .B(n2418), .S(n2413), .Z(n2208) );
  MUX2_X1 U8626 ( .A(n3045), .B(n2419), .S(n2413), .Z(n2207) );
  MUX2_X1 U8627 ( .A(n3046), .B(n2420), .S(n2413), .Z(n2206) );
  MUX2_X1 U8628 ( .A(n3047), .B(n2421), .S(n2413), .Z(n2205) );
  MUX2_X1 U8629 ( .A(n3048), .B(n2422), .S(n2413), .Z(n2204) );
  MUX2_X1 U8630 ( .A(n3049), .B(n2423), .S(n2413), .Z(n2203) );
  MUX2_X1 U8631 ( .A(n3050), .B(n2424), .S(n2413), .Z(n2202) );
  MUX2_X1 U8632 ( .A(n3051), .B(n2425), .S(n2413), .Z(n2201) );
  MUX2_X1 U8633 ( .A(n3052), .B(n2426), .S(n2413), .Z(n2200) );
  MUX2_X1 U8634 ( .A(n3053), .B(n2427), .S(n2413), .Z(n2199) );
  MUX2_X1 U8635 ( .A(n3054), .B(n2428), .S(n2413), .Z(n2198) );
  MUX2_X1 U8636 ( .A(n126), .B(n2429), .S(n2413), .Z(n2197) );
  MUX2_X1 U8637 ( .A(n3055), .B(n2430), .S(n2413), .Z(n2196) );
  MUX2_X1 U8638 ( .A(n3056), .B(n2431), .S(n2413), .Z(n2195) );
  MUX2_X1 U8639 ( .A(n3057), .B(n2432), .S(n2413), .Z(n2194) );
  MUX2_X1 U8640 ( .A(n3058), .B(n2433), .S(n2413), .Z(n2193) );
  MUX2_X1 U8641 ( .A(n3059), .B(n2434), .S(n2413), .Z(n2192) );
  MUX2_X1 U8642 ( .A(n3060), .B(n2435), .S(n2413), .Z(n2191) );
  MUX2_X1 U8643 ( .A(n3061), .B(n2436), .S(n2413), .Z(n2190) );
  MUX2_X1 U8644 ( .A(n825), .B(n2437), .S(n2413), .Z(n2189) );
  MUX2_X1 U8645 ( .A(n826), .B(n2438), .S(n2413), .Z(n2188) );
  MUX2_X1 U8646 ( .A(n827), .B(n2439), .S(n2413), .Z(n2187) );
  MUX2_X1 U8647 ( .A(n828), .B(n2440), .S(n2413), .Z(n2186) );
  MUX2_X1 U8648 ( .A(n829), .B(n2441), .S(n2413), .Z(n2185) );
  MUX2_X1 U8649 ( .A(n830), .B(n2442), .S(n2413), .Z(n2184) );
  MUX2_X1 U8650 ( .A(n831), .B(n2443), .S(n2413), .Z(n2183) );
  MUX2_X1 U8651 ( .A(n832), .B(n2444), .S(n2413), .Z(n2182) );
  MUX2_X1 U8652 ( .A(n2885), .B(n2412), .S(n2446), .Z(n2181) );
  MUX2_X1 U8653 ( .A(n2886), .B(n2414), .S(n2446), .Z(n2180) );
  MUX2_X1 U8654 ( .A(n2887), .B(n2415), .S(n2446), .Z(n2179) );
  MUX2_X1 U8655 ( .A(n2888), .B(n2416), .S(n2446), .Z(n2178) );
  MUX2_X1 U8656 ( .A(n2889), .B(n2417), .S(n2446), .Z(n2177) );
  MUX2_X1 U8657 ( .A(n2890), .B(n2418), .S(n2446), .Z(n2176) );
  MUX2_X1 U8658 ( .A(n2891), .B(n2419), .S(n2446), .Z(n2175) );
  MUX2_X1 U8659 ( .A(n2892), .B(n2420), .S(n2446), .Z(n2174) );
  MUX2_X1 U8660 ( .A(n2893), .B(n2421), .S(n2446), .Z(n2173) );
  MUX2_X1 U8661 ( .A(n2894), .B(n2422), .S(n2446), .Z(n2172) );
  MUX2_X1 U8662 ( .A(n2895), .B(n2423), .S(n2446), .Z(n2171) );
  MUX2_X1 U8663 ( .A(n2896), .B(n2424), .S(n2446), .Z(n2170) );
  MUX2_X1 U8664 ( .A(n2897), .B(n2425), .S(n2446), .Z(n2169) );
  MUX2_X1 U8665 ( .A(n2898), .B(n2426), .S(n2446), .Z(n2168) );
  MUX2_X1 U8666 ( .A(n2899), .B(n2427), .S(n2446), .Z(n2167) );
  MUX2_X1 U8667 ( .A(n2900), .B(n2428), .S(n2446), .Z(n2166) );
  MUX2_X1 U8668 ( .A(n124), .B(n2429), .S(n2446), .Z(n2165) );
  MUX2_X1 U8669 ( .A(n3070), .B(n2430), .S(n2446), .Z(n2164) );
  MUX2_X1 U8670 ( .A(n3071), .B(n2431), .S(n2446), .Z(n2163) );
  MUX2_X1 U8671 ( .A(n3072), .B(n2432), .S(n2446), .Z(n2162) );
  MUX2_X1 U8672 ( .A(n3073), .B(n2433), .S(n2446), .Z(n2161) );
  MUX2_X1 U8673 ( .A(n3074), .B(n2434), .S(n2446), .Z(n2160) );
  MUX2_X1 U8674 ( .A(n3075), .B(n2435), .S(n2446), .Z(n2159) );
  MUX2_X1 U8675 ( .A(n3076), .B(n2436), .S(n2446), .Z(n2158) );
  MUX2_X1 U8676 ( .A(n721), .B(n2437), .S(n2446), .Z(n2157) );
  MUX2_X1 U8677 ( .A(n722), .B(n2438), .S(n2446), .Z(n2156) );
  MUX2_X1 U8678 ( .A(n723), .B(n2439), .S(n2446), .Z(n2155) );
  MUX2_X1 U8679 ( .A(n724), .B(n2440), .S(n2446), .Z(n2154) );
  MUX2_X1 U8680 ( .A(n725), .B(n2441), .S(n2446), .Z(n2153) );
  MUX2_X1 U8681 ( .A(n726), .B(n2442), .S(n2446), .Z(n2152) );
  MUX2_X1 U8682 ( .A(n727), .B(n2443), .S(n2446), .Z(n2151) );
  MUX2_X1 U8683 ( .A(n728), .B(n2444), .S(n2446), .Z(n2150) );
  MUX2_X1 U8684 ( .A(n2901), .B(n2412), .S(n2447), .Z(n2149) );
  MUX2_X1 U8685 ( .A(n2902), .B(n2414), .S(n2447), .Z(n2148) );
  MUX2_X1 U8686 ( .A(n2903), .B(n2415), .S(n2447), .Z(n2147) );
  MUX2_X1 U8687 ( .A(n2904), .B(n2416), .S(n2447), .Z(n2146) );
  MUX2_X1 U8688 ( .A(n2905), .B(n2417), .S(n2447), .Z(n2145) );
  MUX2_X1 U8689 ( .A(n2906), .B(n2418), .S(n2447), .Z(n2144) );
  MUX2_X1 U8690 ( .A(n2907), .B(n2419), .S(n2447), .Z(n2143) );
  MUX2_X1 U8691 ( .A(n2908), .B(n2420), .S(n2447), .Z(n2142) );
  MUX2_X1 U8692 ( .A(n2909), .B(n2421), .S(n2447), .Z(n2141) );
  MUX2_X1 U8693 ( .A(n2910), .B(n2422), .S(n2447), .Z(n2140) );
  MUX2_X1 U8694 ( .A(n2911), .B(n2423), .S(n2447), .Z(n2139) );
  MUX2_X1 U8695 ( .A(n2912), .B(n2424), .S(n2447), .Z(n2138) );
  MUX2_X1 U8696 ( .A(n2913), .B(n2425), .S(n2447), .Z(n2137) );
  MUX2_X1 U8697 ( .A(n2914), .B(n2426), .S(n2447), .Z(n2136) );
  MUX2_X1 U8698 ( .A(n2915), .B(n2427), .S(n2447), .Z(n2135) );
  MUX2_X1 U8699 ( .A(n2916), .B(n2428), .S(n2447), .Z(n2134) );
  MUX2_X1 U8700 ( .A(n122), .B(n2429), .S(n2447), .Z(n2133) );
  MUX2_X1 U8701 ( .A(n21), .B(n2430), .S(n2447), .Z(n2132) );
  MUX2_X1 U8702 ( .A(n29), .B(n2431), .S(n2447), .Z(n2131) );
  MUX2_X1 U8703 ( .A(n37), .B(n2432), .S(n2447), .Z(n2130) );
  MUX2_X1 U8704 ( .A(n45), .B(n2433), .S(n2447), .Z(n2129) );
  MUX2_X1 U8705 ( .A(n53), .B(n2434), .S(n2447), .Z(n2128) );
  MUX2_X1 U8706 ( .A(n61), .B(n2435), .S(n2447), .Z(n2127) );
  MUX2_X1 U8707 ( .A(n69), .B(n2436), .S(n2447), .Z(n2126) );
  MUX2_X1 U8708 ( .A(n2976), .B(n2437), .S(n2447), .Z(n2125) );
  MUX2_X1 U8709 ( .A(n2984), .B(n2438), .S(n2447), .Z(n2124) );
  MUX2_X1 U8710 ( .A(n2992), .B(n2439), .S(n2447), .Z(n2123) );
  MUX2_X1 U8711 ( .A(n3000), .B(n2440), .S(n2447), .Z(n2122) );
  MUX2_X1 U8712 ( .A(n3008), .B(n2441), .S(n2447), .Z(n2121) );
  MUX2_X1 U8713 ( .A(n3016), .B(n2442), .S(n2447), .Z(n2120) );
  MUX2_X1 U8714 ( .A(n3024), .B(n2443), .S(n2447), .Z(n2119) );
  MUX2_X1 U8715 ( .A(n3032), .B(n2444), .S(n2447), .Z(n2118) );
  MUX2_X1 U8716 ( .A(n161), .B(n2412), .S(n2448), .Z(n2117) );
  MUX2_X1 U8717 ( .A(n162), .B(n2414), .S(n2448), .Z(n2116) );
  MUX2_X1 U8718 ( .A(n163), .B(n2415), .S(n2448), .Z(n2115) );
  MUX2_X1 U8719 ( .A(n164), .B(n2416), .S(n2448), .Z(n2114) );
  MUX2_X1 U8720 ( .A(n165), .B(n2417), .S(n2448), .Z(n2113) );
  MUX2_X1 U8721 ( .A(n166), .B(n2418), .S(n2448), .Z(n2112) );
  MUX2_X1 U8722 ( .A(n167), .B(n2419), .S(n2448), .Z(n2111) );
  MUX2_X1 U8723 ( .A(n168), .B(n2420), .S(n2448), .Z(n2110) );
  MUX2_X1 U8724 ( .A(n169), .B(n2421), .S(n2448), .Z(n2109) );
  MUX2_X1 U8725 ( .A(n170), .B(n2422), .S(n2448), .Z(n2108) );
  MUX2_X1 U8726 ( .A(n171), .B(n2423), .S(n2448), .Z(n2107) );
  MUX2_X1 U8727 ( .A(n172), .B(n2424), .S(n2448), .Z(n2106) );
  MUX2_X1 U8728 ( .A(n173), .B(n2425), .S(n2448), .Z(n2105) );
  MUX2_X1 U8729 ( .A(n174), .B(n2426), .S(n2448), .Z(n2104) );
  MUX2_X1 U8730 ( .A(n175), .B(n2427), .S(n2448), .Z(n2103) );
  MUX2_X1 U8731 ( .A(n176), .B(n2428), .S(n2448), .Z(n2102) );
  MUX2_X1 U8732 ( .A(n128), .B(n2429), .S(n2448), .Z(n2101) );
  MUX2_X1 U8733 ( .A(n257), .B(n2430), .S(n2448), .Z(n2100) );
  MUX2_X1 U8734 ( .A(n265), .B(n2431), .S(n2448), .Z(n2099) );
  MUX2_X1 U8735 ( .A(n273), .B(n2432), .S(n2448), .Z(n2098) );
  MUX2_X1 U8736 ( .A(n281), .B(n2433), .S(n2448), .Z(n2097) );
  MUX2_X1 U8737 ( .A(n289), .B(n2434), .S(n2448), .Z(n2096) );
  MUX2_X1 U8738 ( .A(n297), .B(n2435), .S(n2448), .Z(n2095) );
  MUX2_X1 U8739 ( .A(n305), .B(n2436), .S(n2448), .Z(n2094) );
  MUX2_X1 U8740 ( .A(n2975), .B(n2437), .S(n2448), .Z(n2093) );
  MUX2_X1 U8741 ( .A(n2983), .B(n2438), .S(n2448), .Z(n2092) );
  MUX2_X1 U8742 ( .A(n2991), .B(n2439), .S(n2448), .Z(n2091) );
  MUX2_X1 U8743 ( .A(n2999), .B(n2440), .S(n2448), .Z(n2090) );
  MUX2_X1 U8744 ( .A(n3007), .B(n2441), .S(n2448), .Z(n2089) );
  MUX2_X1 U8745 ( .A(n3015), .B(n2442), .S(n2448), .Z(n2088) );
  MUX2_X1 U8746 ( .A(n3023), .B(n2443), .S(n2448), .Z(n2087) );
  MUX2_X1 U8747 ( .A(n3031), .B(n2444), .S(n2448), .Z(n2086) );
  AND2_X1 U8748 ( .A1(n2449), .A2(n2450), .ZN(n2445) );
  MUX2_X1 U8749 ( .A(n73), .B(n2412), .S(n2451), .Z(n2085) );
  MUX2_X1 U8750 ( .A(n74), .B(n2414), .S(n2451), .Z(n2084) );
  MUX2_X1 U8751 ( .A(n75), .B(n2415), .S(n2451), .Z(n2083) );
  MUX2_X1 U8752 ( .A(n76), .B(n2416), .S(n2451), .Z(n2082) );
  MUX2_X1 U8753 ( .A(n77), .B(n2417), .S(n2451), .Z(n2081) );
  MUX2_X1 U8754 ( .A(n78), .B(n2418), .S(n2451), .Z(n2080) );
  MUX2_X1 U8755 ( .A(n79), .B(n2419), .S(n2451), .Z(n2079) );
  MUX2_X1 U8756 ( .A(n80), .B(n2420), .S(n2451), .Z(n2078) );
  MUX2_X1 U8757 ( .A(n81), .B(n2421), .S(n2451), .Z(n2077) );
  MUX2_X1 U8758 ( .A(n82), .B(n2422), .S(n2451), .Z(n2076) );
  MUX2_X1 U8759 ( .A(n83), .B(n2423), .S(n2451), .Z(n2075) );
  MUX2_X1 U8760 ( .A(n84), .B(n2424), .S(n2451), .Z(n2074) );
  MUX2_X1 U8761 ( .A(n85), .B(n2425), .S(n2451), .Z(n2073) );
  MUX2_X1 U8762 ( .A(n86), .B(n2426), .S(n2451), .Z(n2072) );
  MUX2_X1 U8763 ( .A(n87), .B(n2427), .S(n2451), .Z(n2071) );
  MUX2_X1 U8764 ( .A(n88), .B(n2428), .S(n2451), .Z(n2070) );
  MUX2_X1 U8765 ( .A(n362), .B(n2429), .S(n2451), .Z(n2069) );
  MUX2_X1 U8766 ( .A(n2938), .B(n2430), .S(n2451), .Z(n2068) );
  MUX2_X1 U8767 ( .A(n2944), .B(n2431), .S(n2451), .Z(n2067) );
  MUX2_X1 U8768 ( .A(n2950), .B(n2432), .S(n2451), .Z(n2066) );
  MUX2_X1 U8769 ( .A(n2956), .B(n2433), .S(n2451), .Z(n2065) );
  MUX2_X1 U8770 ( .A(n2962), .B(n2434), .S(n2451), .Z(n2064) );
  MUX2_X1 U8771 ( .A(n2968), .B(n2435), .S(n2451), .Z(n2063) );
  MUX2_X1 U8772 ( .A(n2974), .B(n2436), .S(n2451), .Z(n2062) );
  MUX2_X1 U8773 ( .A(n833), .B(n2437), .S(n2451), .Z(n2061) );
  MUX2_X1 U8774 ( .A(n834), .B(n2438), .S(n2451), .Z(n2060) );
  MUX2_X1 U8775 ( .A(n835), .B(n2439), .S(n2451), .Z(n2059) );
  MUX2_X1 U8776 ( .A(n836), .B(n2440), .S(n2451), .Z(n2058) );
  MUX2_X1 U8777 ( .A(n837), .B(n2441), .S(n2451), .Z(n2057) );
  MUX2_X1 U8778 ( .A(n838), .B(n2442), .S(n2451), .Z(n2056) );
  MUX2_X1 U8779 ( .A(n839), .B(n2443), .S(n2451), .Z(n2055) );
  MUX2_X1 U8780 ( .A(n840), .B(n2444), .S(n2451), .Z(n2054) );
  MUX2_X1 U8781 ( .A(n397), .B(n2412), .S(n2453), .Z(n2053) );
  MUX2_X1 U8782 ( .A(n398), .B(n2414), .S(n2453), .Z(n2052) );
  MUX2_X1 U8783 ( .A(n399), .B(n2415), .S(n2453), .Z(n2051) );
  MUX2_X1 U8784 ( .A(n400), .B(n2416), .S(n2453), .Z(n2050) );
  MUX2_X1 U8785 ( .A(n401), .B(n2417), .S(n2453), .Z(n2049) );
  MUX2_X1 U8786 ( .A(n402), .B(n2418), .S(n2453), .Z(n2048) );
  MUX2_X1 U8787 ( .A(n403), .B(n2419), .S(n2453), .Z(n2047) );
  MUX2_X1 U8788 ( .A(n404), .B(n2420), .S(n2453), .Z(n2046) );
  MUX2_X1 U8789 ( .A(n405), .B(n2421), .S(n2453), .Z(n2045) );
  MUX2_X1 U8790 ( .A(n406), .B(n2422), .S(n2453), .Z(n2044) );
  MUX2_X1 U8791 ( .A(n407), .B(n2423), .S(n2453), .Z(n2043) );
  MUX2_X1 U8792 ( .A(n408), .B(n2424), .S(n2453), .Z(n2042) );
  MUX2_X1 U8793 ( .A(n409), .B(n2425), .S(n2453), .Z(n2041) );
  MUX2_X1 U8794 ( .A(n410), .B(n2426), .S(n2453), .Z(n2040) );
  MUX2_X1 U8795 ( .A(n411), .B(n2427), .S(n2453), .Z(n2039) );
  MUX2_X1 U8796 ( .A(n412), .B(n2428), .S(n2453), .Z(n2038) );
  MUX2_X1 U8797 ( .A(n360), .B(n2429), .S(n2453), .Z(n2037) );
  MUX2_X1 U8798 ( .A(n2937), .B(n2430), .S(n2453), .Z(n2036) );
  MUX2_X1 U8799 ( .A(n2943), .B(n2431), .S(n2453), .Z(n2035) );
  MUX2_X1 U8800 ( .A(n2949), .B(n2432), .S(n2453), .Z(n2034) );
  MUX2_X1 U8801 ( .A(n2955), .B(n2433), .S(n2453), .Z(n2033) );
  MUX2_X1 U8802 ( .A(n2961), .B(n2434), .S(n2453), .Z(n2032) );
  MUX2_X1 U8803 ( .A(n2967), .B(n2435), .S(n2453), .Z(n2031) );
  MUX2_X1 U8804 ( .A(n2973), .B(n2436), .S(n2453), .Z(n2030) );
  MUX2_X1 U8805 ( .A(n729), .B(n2437), .S(n2453), .Z(n2029) );
  MUX2_X1 U8806 ( .A(n730), .B(n2438), .S(n2453), .Z(n2028) );
  MUX2_X1 U8807 ( .A(n731), .B(n2439), .S(n2453), .Z(n2027) );
  MUX2_X1 U8808 ( .A(n732), .B(n2440), .S(n2453), .Z(n2026) );
  MUX2_X1 U8809 ( .A(n733), .B(n2441), .S(n2453), .Z(n2025) );
  MUX2_X1 U8810 ( .A(n734), .B(n2442), .S(n2453), .Z(n2024) );
  MUX2_X1 U8811 ( .A(n735), .B(n2443), .S(n2453), .Z(n2023) );
  MUX2_X1 U8812 ( .A(n736), .B(n2444), .S(n2453), .Z(n2022) );
  MUX2_X1 U8813 ( .A(n309), .B(n2412), .S(n2454), .Z(n2021) );
  MUX2_X1 U8814 ( .A(n310), .B(n2414), .S(n2454), .Z(n2020) );
  MUX2_X1 U8815 ( .A(n311), .B(n2415), .S(n2454), .Z(n2019) );
  MUX2_X1 U8816 ( .A(n312), .B(n2416), .S(n2454), .Z(n2018) );
  MUX2_X1 U8817 ( .A(n313), .B(n2417), .S(n2454), .Z(n2017) );
  MUX2_X1 U8818 ( .A(n314), .B(n2418), .S(n2454), .Z(n2016) );
  MUX2_X1 U8819 ( .A(n315), .B(n2419), .S(n2454), .Z(n2015) );
  MUX2_X1 U8820 ( .A(n316), .B(n2420), .S(n2454), .Z(n2014) );
  MUX2_X1 U8821 ( .A(n317), .B(n2421), .S(n2454), .Z(n2013) );
  MUX2_X1 U8822 ( .A(n318), .B(n2422), .S(n2454), .Z(n2012) );
  MUX2_X1 U8823 ( .A(n319), .B(n2423), .S(n2454), .Z(n2011) );
  MUX2_X1 U8824 ( .A(n320), .B(n2424), .S(n2454), .Z(n2010) );
  MUX2_X1 U8825 ( .A(n321), .B(n2425), .S(n2454), .Z(n2009) );
  MUX2_X1 U8826 ( .A(n322), .B(n2426), .S(n2454), .Z(n2008) );
  MUX2_X1 U8827 ( .A(n323), .B(n2427), .S(n2454), .Z(n2007) );
  MUX2_X1 U8828 ( .A(n324), .B(n2428), .S(n2454), .Z(n2006) );
  MUX2_X1 U8829 ( .A(n358), .B(n2429), .S(n2454), .Z(n2005) );
  MUX2_X1 U8830 ( .A(n22), .B(n2430), .S(n2454), .Z(n2004) );
  MUX2_X1 U8831 ( .A(n30), .B(n2431), .S(n2454), .Z(n2003) );
  MUX2_X1 U8832 ( .A(n38), .B(n2432), .S(n2454), .Z(n2002) );
  MUX2_X1 U8833 ( .A(n46), .B(n2433), .S(n2454), .Z(n2001) );
  MUX2_X1 U8834 ( .A(n54), .B(n2434), .S(n2454), .Z(n2000) );
  MUX2_X1 U8835 ( .A(n62), .B(n2435), .S(n2454), .Z(n1999) );
  MUX2_X1 U8836 ( .A(n70), .B(n2436), .S(n2454), .Z(n1998) );
  MUX2_X1 U8837 ( .A(n2978), .B(n2437), .S(n2454), .Z(n1997) );
  MUX2_X1 U8838 ( .A(n2986), .B(n2438), .S(n2454), .Z(n1996) );
  MUX2_X1 U8839 ( .A(n2994), .B(n2439), .S(n2454), .Z(n1995) );
  MUX2_X1 U8840 ( .A(n3002), .B(n2440), .S(n2454), .Z(n1994) );
  MUX2_X1 U8841 ( .A(n3010), .B(n2441), .S(n2454), .Z(n1993) );
  MUX2_X1 U8842 ( .A(n3018), .B(n2442), .S(n2454), .Z(n1992) );
  MUX2_X1 U8843 ( .A(n3026), .B(n2443), .S(n2454), .Z(n1991) );
  MUX2_X1 U8844 ( .A(n3034), .B(n2444), .S(n2454), .Z(n1990) );
  MUX2_X1 U8845 ( .A(n2917), .B(n2412), .S(n2455), .Z(n1989) );
  MUX2_X1 U8846 ( .A(n2918), .B(n2414), .S(n2455), .Z(n1988) );
  MUX2_X1 U8847 ( .A(n2919), .B(n2415), .S(n2455), .Z(n1987) );
  MUX2_X1 U8848 ( .A(n2920), .B(n2416), .S(n2455), .Z(n1986) );
  MUX2_X1 U8849 ( .A(n2921), .B(n2417), .S(n2455), .Z(n1985) );
  MUX2_X1 U8850 ( .A(n2922), .B(n2418), .S(n2455), .Z(n1984) );
  MUX2_X1 U8851 ( .A(n2923), .B(n2419), .S(n2455), .Z(n1983) );
  MUX2_X1 U8852 ( .A(n2924), .B(n2420), .S(n2455), .Z(n1982) );
  MUX2_X1 U8853 ( .A(n2925), .B(n2421), .S(n2455), .Z(n1981) );
  MUX2_X1 U8854 ( .A(n2926), .B(n2422), .S(n2455), .Z(n1980) );
  MUX2_X1 U8855 ( .A(n2927), .B(n2423), .S(n2455), .Z(n1979) );
  MUX2_X1 U8856 ( .A(n2928), .B(n2424), .S(n2455), .Z(n1978) );
  MUX2_X1 U8857 ( .A(n2929), .B(n2425), .S(n2455), .Z(n1977) );
  MUX2_X1 U8858 ( .A(n2930), .B(n2426), .S(n2455), .Z(n1976) );
  MUX2_X1 U8859 ( .A(n2931), .B(n2427), .S(n2455), .Z(n1975) );
  MUX2_X1 U8860 ( .A(n2932), .B(n2428), .S(n2455), .Z(n1974) );
  MUX2_X1 U8861 ( .A(n364), .B(n2429), .S(n2455), .Z(n1973) );
  MUX2_X1 U8862 ( .A(n258), .B(n2430), .S(n2455), .Z(n1972) );
  MUX2_X1 U8863 ( .A(n266), .B(n2431), .S(n2455), .Z(n1971) );
  MUX2_X1 U8864 ( .A(n274), .B(n2432), .S(n2455), .Z(n1970) );
  MUX2_X1 U8865 ( .A(n282), .B(n2433), .S(n2455), .Z(n1969) );
  MUX2_X1 U8866 ( .A(n290), .B(n2434), .S(n2455), .Z(n1968) );
  MUX2_X1 U8867 ( .A(n298), .B(n2435), .S(n2455), .Z(n1967) );
  MUX2_X1 U8868 ( .A(n306), .B(n2436), .S(n2455), .Z(n1966) );
  MUX2_X1 U8869 ( .A(n2977), .B(n2437), .S(n2455), .Z(n1965) );
  MUX2_X1 U8870 ( .A(n2985), .B(n2438), .S(n2455), .Z(n1964) );
  MUX2_X1 U8871 ( .A(n2993), .B(n2439), .S(n2455), .Z(n1963) );
  MUX2_X1 U8872 ( .A(n3001), .B(n2440), .S(n2455), .Z(n1962) );
  MUX2_X1 U8873 ( .A(n3009), .B(n2441), .S(n2455), .Z(n1961) );
  MUX2_X1 U8874 ( .A(n3017), .B(n2442), .S(n2455), .Z(n1960) );
  MUX2_X1 U8875 ( .A(n3025), .B(n2443), .S(n2455), .Z(n1959) );
  MUX2_X1 U8876 ( .A(n3033), .B(n2444), .S(n2455), .Z(n1958) );
  AND2_X1 U8877 ( .A1(n2449), .A2(n2456), .ZN(n2452) );
  MUX2_X1 U8878 ( .A(n325), .B(n2412), .S(n2457), .Z(n1957) );
  MUX2_X1 U8879 ( .A(n326), .B(n2414), .S(n2457), .Z(n1956) );
  MUX2_X1 U8880 ( .A(n327), .B(n2415), .S(n2457), .Z(n1955) );
  MUX2_X1 U8881 ( .A(n328), .B(n2416), .S(n2457), .Z(n1954) );
  MUX2_X1 U8882 ( .A(n329), .B(n2417), .S(n2457), .Z(n1953) );
  MUX2_X1 U8883 ( .A(n330), .B(n2418), .S(n2457), .Z(n1952) );
  MUX2_X1 U8884 ( .A(n331), .B(n2419), .S(n2457), .Z(n1951) );
  MUX2_X1 U8885 ( .A(n332), .B(n2420), .S(n2457), .Z(n1950) );
  MUX2_X1 U8886 ( .A(n333), .B(n2421), .S(n2457), .Z(n1949) );
  MUX2_X1 U8887 ( .A(n334), .B(n2422), .S(n2457), .Z(n1948) );
  MUX2_X1 U8888 ( .A(n335), .B(n2423), .S(n2457), .Z(n1947) );
  MUX2_X1 U8889 ( .A(n336), .B(n2424), .S(n2457), .Z(n1946) );
  MUX2_X1 U8890 ( .A(n337), .B(n2425), .S(n2457), .Z(n1945) );
  MUX2_X1 U8891 ( .A(n338), .B(n2426), .S(n2457), .Z(n1944) );
  MUX2_X1 U8892 ( .A(n339), .B(n2427), .S(n2457), .Z(n1943) );
  MUX2_X1 U8893 ( .A(n340), .B(n2428), .S(n2457), .Z(n1942) );
  MUX2_X1 U8894 ( .A(n841), .B(n2429), .S(n2457), .Z(n1941) );
  MUX2_X1 U8895 ( .A(n24), .B(n2430), .S(n2457), .Z(n1940) );
  MUX2_X1 U8896 ( .A(n32), .B(n2431), .S(n2457), .Z(n1939) );
  MUX2_X1 U8897 ( .A(n40), .B(n2432), .S(n2457), .Z(n1938) );
  MUX2_X1 U8898 ( .A(n48), .B(n2433), .S(n2457), .Z(n1937) );
  MUX2_X1 U8899 ( .A(n56), .B(n2434), .S(n2457), .Z(n1936) );
  MUX2_X1 U8900 ( .A(n64), .B(n2435), .S(n2457), .Z(n1935) );
  MUX2_X1 U8901 ( .A(n72), .B(n2436), .S(n2457), .Z(n1934) );
  MUX2_X1 U8902 ( .A(n842), .B(n2437), .S(n2457), .Z(n1933) );
  MUX2_X1 U8903 ( .A(n843), .B(n2438), .S(n2457), .Z(n1932) );
  MUX2_X1 U8904 ( .A(n844), .B(n2439), .S(n2457), .Z(n1931) );
  MUX2_X1 U8905 ( .A(n845), .B(n2440), .S(n2457), .Z(n1930) );
  MUX2_X1 U8906 ( .A(n846), .B(n2441), .S(n2457), .Z(n1929) );
  MUX2_X1 U8907 ( .A(n847), .B(n2442), .S(n2457), .Z(n1928) );
  MUX2_X1 U8908 ( .A(n848), .B(n2443), .S(n2457), .Z(n1927) );
  MUX2_X1 U8909 ( .A(n849), .B(n2444), .S(n2457), .Z(n1926) );
  MUX2_X1 U8910 ( .A(n737), .B(n2412), .S(n2459), .Z(n1925) );
  MUX2_X1 U8911 ( .A(n738), .B(n2414), .S(n2459), .Z(n1924) );
  MUX2_X1 U8912 ( .A(n739), .B(n2415), .S(n2459), .Z(n1923) );
  MUX2_X1 U8913 ( .A(n740), .B(n2416), .S(n2459), .Z(n1922) );
  MUX2_X1 U8914 ( .A(n741), .B(n2417), .S(n2459), .Z(n1921) );
  MUX2_X1 U8915 ( .A(n742), .B(n2418), .S(n2459), .Z(n1920) );
  MUX2_X1 U8916 ( .A(n743), .B(n2419), .S(n2459), .Z(n1919) );
  MUX2_X1 U8917 ( .A(n744), .B(n2420), .S(n2459), .Z(n1918) );
  MUX2_X1 U8918 ( .A(n745), .B(n2421), .S(n2459), .Z(n1917) );
  MUX2_X1 U8919 ( .A(n746), .B(n2422), .S(n2459), .Z(n1916) );
  MUX2_X1 U8920 ( .A(n747), .B(n2423), .S(n2459), .Z(n1915) );
  MUX2_X1 U8921 ( .A(n748), .B(n2424), .S(n2459), .Z(n1914) );
  MUX2_X1 U8922 ( .A(n749), .B(n2425), .S(n2459), .Z(n1913) );
  MUX2_X1 U8923 ( .A(n750), .B(n2426), .S(n2459), .Z(n1912) );
  MUX2_X1 U8924 ( .A(n751), .B(n2427), .S(n2459), .Z(n1911) );
  MUX2_X1 U8925 ( .A(n752), .B(n2428), .S(n2459), .Z(n1910) );
  MUX2_X1 U8926 ( .A(n850), .B(n2429), .S(n2459), .Z(n1909) );
  MUX2_X1 U8927 ( .A(n260), .B(n2430), .S(n2459), .Z(n1908) );
  MUX2_X1 U8928 ( .A(n268), .B(n2431), .S(n2459), .Z(n1907) );
  MUX2_X1 U8929 ( .A(n276), .B(n2432), .S(n2459), .Z(n1906) );
  MUX2_X1 U8930 ( .A(n284), .B(n2433), .S(n2459), .Z(n1905) );
  MUX2_X1 U8931 ( .A(n292), .B(n2434), .S(n2459), .Z(n1904) );
  MUX2_X1 U8932 ( .A(n300), .B(n2435), .S(n2459), .Z(n1903) );
  MUX2_X1 U8933 ( .A(n308), .B(n2436), .S(n2459), .Z(n1902) );
  MUX2_X1 U8934 ( .A(n753), .B(n2437), .S(n2459), .Z(n1901) );
  MUX2_X1 U8935 ( .A(n754), .B(n2438), .S(n2459), .Z(n1900) );
  MUX2_X1 U8936 ( .A(n755), .B(n2439), .S(n2459), .Z(n1899) );
  MUX2_X1 U8937 ( .A(n756), .B(n2440), .S(n2459), .Z(n1898) );
  MUX2_X1 U8938 ( .A(n757), .B(n2441), .S(n2459), .Z(n1897) );
  MUX2_X1 U8939 ( .A(n758), .B(n2442), .S(n2459), .Z(n1896) );
  MUX2_X1 U8940 ( .A(n759), .B(n2443), .S(n2459), .Z(n1895) );
  MUX2_X1 U8941 ( .A(n760), .B(n2444), .S(n2459), .Z(n1894) );
  MUX2_X1 U8942 ( .A(n89), .B(n2412), .S(n2460), .Z(n1893) );
  MUX2_X1 U8943 ( .A(n90), .B(n2414), .S(n2460), .Z(n1892) );
  MUX2_X1 U8944 ( .A(n91), .B(n2415), .S(n2460), .Z(n1891) );
  MUX2_X1 U8945 ( .A(n92), .B(n2416), .S(n2460), .Z(n1890) );
  MUX2_X1 U8946 ( .A(n93), .B(n2417), .S(n2460), .Z(n1889) );
  MUX2_X1 U8947 ( .A(n94), .B(n2418), .S(n2460), .Z(n1888) );
  MUX2_X1 U8948 ( .A(n95), .B(n2419), .S(n2460), .Z(n1887) );
  MUX2_X1 U8949 ( .A(n96), .B(n2420), .S(n2460), .Z(n1886) );
  MUX2_X1 U8950 ( .A(n97), .B(n2421), .S(n2460), .Z(n1885) );
  MUX2_X1 U8951 ( .A(n98), .B(n2422), .S(n2460), .Z(n1884) );
  MUX2_X1 U8952 ( .A(n99), .B(n2423), .S(n2460), .Z(n1883) );
  MUX2_X1 U8953 ( .A(n100), .B(n2424), .S(n2460), .Z(n1882) );
  MUX2_X1 U8954 ( .A(n101), .B(n2425), .S(n2460), .Z(n1881) );
  MUX2_X1 U8955 ( .A(n102), .B(n2426), .S(n2460), .Z(n1880) );
  MUX2_X1 U8956 ( .A(n103), .B(n2427), .S(n2460), .Z(n1879) );
  MUX2_X1 U8957 ( .A(n104), .B(n2428), .S(n2460), .Z(n1878) );
  MUX2_X1 U8958 ( .A(n851), .B(n2429), .S(n2460), .Z(n1877) );
  MUX2_X1 U8959 ( .A(n473), .B(n2430), .S(n2460), .Z(n1876) );
  MUX2_X1 U8960 ( .A(n474), .B(n2431), .S(n2460), .Z(n1875) );
  MUX2_X1 U8961 ( .A(n475), .B(n2432), .S(n2460), .Z(n1874) );
  MUX2_X1 U8962 ( .A(n476), .B(n2433), .S(n2460), .Z(n1873) );
  MUX2_X1 U8963 ( .A(n477), .B(n2434), .S(n2460), .Z(n1872) );
  MUX2_X1 U8964 ( .A(n478), .B(n2435), .S(n2460), .Z(n1871) );
  MUX2_X1 U8965 ( .A(n479), .B(n2436), .S(n2460), .Z(n1870) );
  MUX2_X1 U8966 ( .A(n365), .B(n2437), .S(n2460), .Z(n1869) );
  MUX2_X1 U8967 ( .A(n369), .B(n2438), .S(n2460), .Z(n1868) );
  MUX2_X1 U8968 ( .A(n373), .B(n2439), .S(n2460), .Z(n1867) );
  MUX2_X1 U8969 ( .A(n377), .B(n2440), .S(n2460), .Z(n1866) );
  MUX2_X1 U8970 ( .A(n381), .B(n2441), .S(n2460), .Z(n1865) );
  MUX2_X1 U8971 ( .A(n385), .B(n2442), .S(n2460), .Z(n1864) );
  MUX2_X1 U8972 ( .A(n389), .B(n2443), .S(n2460), .Z(n1863) );
  MUX2_X1 U8973 ( .A(n393), .B(n2444), .S(n2460), .Z(n1862) );
  MUX2_X1 U8974 ( .A(n852), .B(n2412), .S(n2461), .Z(n1861) );
  MUX2_X1 U8975 ( .A(n853), .B(n2414), .S(n2461), .Z(n1860) );
  MUX2_X1 U8976 ( .A(n854), .B(n2415), .S(n2461), .Z(n1859) );
  MUX2_X1 U8977 ( .A(n855), .B(n2416), .S(n2461), .Z(n1858) );
  MUX2_X1 U8978 ( .A(n856), .B(n2417), .S(n2461), .Z(n1857) );
  MUX2_X1 U8979 ( .A(n857), .B(n2418), .S(n2461), .Z(n1856) );
  MUX2_X1 U8980 ( .A(n858), .B(n2419), .S(n2461), .Z(n1855) );
  MUX2_X1 U8981 ( .A(n859), .B(n2420), .S(n2461), .Z(n1854) );
  MUX2_X1 U8982 ( .A(n860), .B(n2421), .S(n2461), .Z(n1853) );
  MUX2_X1 U8983 ( .A(n861), .B(n2422), .S(n2461), .Z(n1852) );
  MUX2_X1 U8984 ( .A(n862), .B(n2423), .S(n2461), .Z(n1851) );
  MUX2_X1 U8985 ( .A(n863), .B(n2424), .S(n2461), .Z(n1850) );
  MUX2_X1 U8986 ( .A(n864), .B(n2425), .S(n2461), .Z(n1849) );
  MUX2_X1 U8987 ( .A(n865), .B(n2426), .S(n2461), .Z(n1848) );
  MUX2_X1 U8988 ( .A(n866), .B(n2427), .S(n2461), .Z(n1847) );
  MUX2_X1 U8989 ( .A(n867), .B(n2428), .S(n2461), .Z(n1846) );
  MUX2_X1 U8990 ( .A(n868), .B(n2429), .S(n2461), .Z(n1845) );
  MUX2_X1 U8991 ( .A(n597), .B(n2430), .S(n2461), .Z(n1844) );
  MUX2_X1 U8992 ( .A(n598), .B(n2431), .S(n2461), .Z(n1843) );
  MUX2_X1 U8993 ( .A(n599), .B(n2432), .S(n2461), .Z(n1842) );
  MUX2_X1 U8994 ( .A(n600), .B(n2433), .S(n2461), .Z(n1841) );
  MUX2_X1 U8995 ( .A(n601), .B(n2434), .S(n2461), .Z(n1840) );
  MUX2_X1 U8996 ( .A(n602), .B(n2435), .S(n2461), .Z(n1839) );
  MUX2_X1 U8997 ( .A(n603), .B(n2436), .S(n2461), .Z(n1838) );
  MUX2_X1 U8998 ( .A(n129), .B(n2437), .S(n2461), .Z(n1837) );
  MUX2_X1 U8999 ( .A(n133), .B(n2438), .S(n2461), .Z(n1836) );
  MUX2_X1 U9000 ( .A(n137), .B(n2439), .S(n2461), .Z(n1835) );
  MUX2_X1 U9001 ( .A(n141), .B(n2440), .S(n2461), .Z(n1834) );
  MUX2_X1 U9002 ( .A(n145), .B(n2441), .S(n2461), .Z(n1833) );
  MUX2_X1 U9003 ( .A(n149), .B(n2442), .S(n2461), .Z(n1832) );
  MUX2_X1 U9004 ( .A(n153), .B(n2443), .S(n2461), .Z(n1831) );
  MUX2_X1 U9005 ( .A(n157), .B(n2444), .S(n2461), .Z(n1830) );
  AND2_X1 U9006 ( .A1(n2449), .A2(n2462), .ZN(n2458) );
  MUX2_X1 U9007 ( .A(n105), .B(n2412), .S(n2463), .Z(n1829) );
  MUX2_X1 U9008 ( .A(n106), .B(n2414), .S(n2463), .Z(n1828) );
  MUX2_X1 U9009 ( .A(n107), .B(n2415), .S(n2463), .Z(n1827) );
  MUX2_X1 U9010 ( .A(n108), .B(n2416), .S(n2463), .Z(n1826) );
  MUX2_X1 U9011 ( .A(n109), .B(n2417), .S(n2463), .Z(n1825) );
  MUX2_X1 U9012 ( .A(n110), .B(n2418), .S(n2463), .Z(n1824) );
  MUX2_X1 U9013 ( .A(n111), .B(n2419), .S(n2463), .Z(n1823) );
  MUX2_X1 U9014 ( .A(n112), .B(n2420), .S(n2463), .Z(n1822) );
  MUX2_X1 U9015 ( .A(n113), .B(n2421), .S(n2463), .Z(n1821) );
  MUX2_X1 U9016 ( .A(n114), .B(n2422), .S(n2463), .Z(n1820) );
  MUX2_X1 U9017 ( .A(n115), .B(n2423), .S(n2463), .Z(n1819) );
  MUX2_X1 U9018 ( .A(n116), .B(n2424), .S(n2463), .Z(n1818) );
  MUX2_X1 U9019 ( .A(n117), .B(n2425), .S(n2463), .Z(n1817) );
  MUX2_X1 U9020 ( .A(n118), .B(n2426), .S(n2463), .Z(n1816) );
  MUX2_X1 U9021 ( .A(n119), .B(n2427), .S(n2463), .Z(n1815) );
  MUX2_X1 U9022 ( .A(n120), .B(n2428), .S(n2463), .Z(n1814) );
  MUX2_X1 U9023 ( .A(n761), .B(n2429), .S(n2463), .Z(n1813) );
  MUX2_X1 U9024 ( .A(n23), .B(n2430), .S(n2463), .Z(n1812) );
  MUX2_X1 U9025 ( .A(n31), .B(n2431), .S(n2463), .Z(n1811) );
  MUX2_X1 U9026 ( .A(n39), .B(n2432), .S(n2463), .Z(n1810) );
  MUX2_X1 U9027 ( .A(n47), .B(n2433), .S(n2463), .Z(n1809) );
  MUX2_X1 U9028 ( .A(n55), .B(n2434), .S(n2463), .Z(n1808) );
  MUX2_X1 U9029 ( .A(n63), .B(n2435), .S(n2463), .Z(n1807) );
  MUX2_X1 U9030 ( .A(n71), .B(n2436), .S(n2463), .Z(n1806) );
  MUX2_X1 U9031 ( .A(n869), .B(n2437), .S(n2463), .Z(n1805) );
  MUX2_X1 U9032 ( .A(n870), .B(n2438), .S(n2463), .Z(n1804) );
  MUX2_X1 U9033 ( .A(n871), .B(n2439), .S(n2463), .Z(n1803) );
  MUX2_X1 U9034 ( .A(n872), .B(n2440), .S(n2463), .Z(n1802) );
  MUX2_X1 U9035 ( .A(n873), .B(n2441), .S(n2463), .Z(n1801) );
  MUX2_X1 U9036 ( .A(n874), .B(n2442), .S(n2463), .Z(n1800) );
  MUX2_X1 U9037 ( .A(n875), .B(n2443), .S(n2463), .Z(n1799) );
  MUX2_X1 U9038 ( .A(n876), .B(n2444), .S(n2463), .Z(n1798) );
  MUX2_X1 U9039 ( .A(n877), .B(n2412), .S(n2465), .Z(n1797) );
  MUX2_X1 U9040 ( .A(n878), .B(n2414), .S(n2465), .Z(n1796) );
  MUX2_X1 U9041 ( .A(n879), .B(n2415), .S(n2465), .Z(n1795) );
  MUX2_X1 U9042 ( .A(n880), .B(n2416), .S(n2465), .Z(n1794) );
  MUX2_X1 U9043 ( .A(n881), .B(n2417), .S(n2465), .Z(n1793) );
  MUX2_X1 U9044 ( .A(n882), .B(n2418), .S(n2465), .Z(n1792) );
  MUX2_X1 U9045 ( .A(n883), .B(n2419), .S(n2465), .Z(n1791) );
  MUX2_X1 U9046 ( .A(n884), .B(n2420), .S(n2465), .Z(n1790) );
  MUX2_X1 U9047 ( .A(n885), .B(n2421), .S(n2465), .Z(n1789) );
  MUX2_X1 U9048 ( .A(n886), .B(n2422), .S(n2465), .Z(n1788) );
  MUX2_X1 U9049 ( .A(n887), .B(n2423), .S(n2465), .Z(n1787) );
  MUX2_X1 U9050 ( .A(n888), .B(n2424), .S(n2465), .Z(n1786) );
  MUX2_X1 U9051 ( .A(n889), .B(n2425), .S(n2465), .Z(n1785) );
  MUX2_X1 U9052 ( .A(n890), .B(n2426), .S(n2465), .Z(n1784) );
  MUX2_X1 U9053 ( .A(n891), .B(n2427), .S(n2465), .Z(n1783) );
  MUX2_X1 U9054 ( .A(n892), .B(n2428), .S(n2465), .Z(n1782) );
  MUX2_X1 U9055 ( .A(n762), .B(n2429), .S(n2465), .Z(n1781) );
  MUX2_X1 U9056 ( .A(n259), .B(n2430), .S(n2465), .Z(n1780) );
  MUX2_X1 U9057 ( .A(n267), .B(n2431), .S(n2465), .Z(n1779) );
  MUX2_X1 U9058 ( .A(n275), .B(n2432), .S(n2465), .Z(n1778) );
  MUX2_X1 U9059 ( .A(n283), .B(n2433), .S(n2465), .Z(n1777) );
  MUX2_X1 U9060 ( .A(n291), .B(n2434), .S(n2465), .Z(n1776) );
  MUX2_X1 U9061 ( .A(n299), .B(n2435), .S(n2465), .Z(n1775) );
  MUX2_X1 U9062 ( .A(n307), .B(n2436), .S(n2465), .Z(n1774) );
  MUX2_X1 U9063 ( .A(n763), .B(n2437), .S(n2465), .Z(n1773) );
  MUX2_X1 U9064 ( .A(n764), .B(n2438), .S(n2465), .Z(n1772) );
  MUX2_X1 U9065 ( .A(n765), .B(n2439), .S(n2465), .Z(n1771) );
  MUX2_X1 U9066 ( .A(n766), .B(n2440), .S(n2465), .Z(n1770) );
  MUX2_X1 U9067 ( .A(n767), .B(n2441), .S(n2465), .Z(n1769) );
  MUX2_X1 U9068 ( .A(n768), .B(n2442), .S(n2465), .Z(n1768) );
  MUX2_X1 U9069 ( .A(n769), .B(n2443), .S(n2465), .Z(n1767) );
  MUX2_X1 U9070 ( .A(n770), .B(n2444), .S(n2465), .Z(n1766) );
  MUX2_X1 U9071 ( .A(n893), .B(n2412), .S(n2466), .Z(n1765) );
  MUX2_X1 U9072 ( .A(n894), .B(n2414), .S(n2466), .Z(n1764) );
  MUX2_X1 U9073 ( .A(n895), .B(n2415), .S(n2466), .Z(n1763) );
  MUX2_X1 U9074 ( .A(n896), .B(n2416), .S(n2466), .Z(n1762) );
  MUX2_X1 U9075 ( .A(n897), .B(n2417), .S(n2466), .Z(n1761) );
  MUX2_X1 U9076 ( .A(n898), .B(n2418), .S(n2466), .Z(n1760) );
  MUX2_X1 U9077 ( .A(n899), .B(n2419), .S(n2466), .Z(n1759) );
  MUX2_X1 U9078 ( .A(n900), .B(n2420), .S(n2466), .Z(n1758) );
  MUX2_X1 U9079 ( .A(n901), .B(n2421), .S(n2466), .Z(n1757) );
  MUX2_X1 U9080 ( .A(n902), .B(n2422), .S(n2466), .Z(n1756) );
  MUX2_X1 U9081 ( .A(n903), .B(n2423), .S(n2466), .Z(n1755) );
  MUX2_X1 U9082 ( .A(n904), .B(n2424), .S(n2466), .Z(n1754) );
  MUX2_X1 U9083 ( .A(n905), .B(n2425), .S(n2466), .Z(n1753) );
  MUX2_X1 U9084 ( .A(n906), .B(n2426), .S(n2466), .Z(n1752) );
  MUX2_X1 U9085 ( .A(n907), .B(n2427), .S(n2466), .Z(n1751) );
  MUX2_X1 U9086 ( .A(n908), .B(n2428), .S(n2466), .Z(n1750) );
  MUX2_X1 U9087 ( .A(n771), .B(n2429), .S(n2466), .Z(n1749) );
  MUX2_X1 U9088 ( .A(n480), .B(n2430), .S(n2466), .Z(n1748) );
  MUX2_X1 U9089 ( .A(n481), .B(n2431), .S(n2466), .Z(n1747) );
  MUX2_X1 U9090 ( .A(n482), .B(n2432), .S(n2466), .Z(n1746) );
  MUX2_X1 U9091 ( .A(n483), .B(n2433), .S(n2466), .Z(n1745) );
  MUX2_X1 U9092 ( .A(n484), .B(n2434), .S(n2466), .Z(n1744) );
  MUX2_X1 U9093 ( .A(n485), .B(n2435), .S(n2466), .Z(n1743) );
  MUX2_X1 U9094 ( .A(n486), .B(n2436), .S(n2466), .Z(n1742) );
  MUX2_X1 U9095 ( .A(n366), .B(n2437), .S(n2466), .Z(n1741) );
  MUX2_X1 U9096 ( .A(n370), .B(n2438), .S(n2466), .Z(n1740) );
  MUX2_X1 U9097 ( .A(n374), .B(n2439), .S(n2466), .Z(n1739) );
  MUX2_X1 U9098 ( .A(n378), .B(n2440), .S(n2466), .Z(n1738) );
  MUX2_X1 U9099 ( .A(n382), .B(n2441), .S(n2466), .Z(n1737) );
  MUX2_X1 U9100 ( .A(n386), .B(n2442), .S(n2466), .Z(n1736) );
  MUX2_X1 U9101 ( .A(n390), .B(n2443), .S(n2466), .Z(n1735) );
  MUX2_X1 U9102 ( .A(n394), .B(n2444), .S(n2466), .Z(n1734) );
  MUX2_X1 U9103 ( .A(n772), .B(n2412), .S(n2467), .Z(n1733) );
  MUX2_X1 U9104 ( .A(n773), .B(n2414), .S(n2467), .Z(n1732) );
  MUX2_X1 U9105 ( .A(n774), .B(n2415), .S(n2467), .Z(n1731) );
  MUX2_X1 U9106 ( .A(n775), .B(n2416), .S(n2467), .Z(n1730) );
  MUX2_X1 U9107 ( .A(n776), .B(n2417), .S(n2467), .Z(n1729) );
  MUX2_X1 U9108 ( .A(n777), .B(n2418), .S(n2467), .Z(n1728) );
  MUX2_X1 U9109 ( .A(n778), .B(n2419), .S(n2467), .Z(n1727) );
  MUX2_X1 U9110 ( .A(n779), .B(n2420), .S(n2467), .Z(n1726) );
  MUX2_X1 U9111 ( .A(n780), .B(n2421), .S(n2467), .Z(n1725) );
  MUX2_X1 U9112 ( .A(n781), .B(n2422), .S(n2467), .Z(n1724) );
  MUX2_X1 U9113 ( .A(n782), .B(n2423), .S(n2467), .Z(n1723) );
  MUX2_X1 U9114 ( .A(n783), .B(n2424), .S(n2467), .Z(n1722) );
  MUX2_X1 U9115 ( .A(n784), .B(n2425), .S(n2467), .Z(n1721) );
  MUX2_X1 U9116 ( .A(n785), .B(n2426), .S(n2467), .Z(n1720) );
  MUX2_X1 U9117 ( .A(n786), .B(n2427), .S(n2467), .Z(n1719) );
  MUX2_X1 U9118 ( .A(n787), .B(n2428), .S(n2467), .Z(n1718) );
  MUX2_X1 U9119 ( .A(n788), .B(n2429), .S(n2467), .Z(n1717) );
  MUX2_X1 U9120 ( .A(n604), .B(n2430), .S(n2467), .Z(n1716) );
  MUX2_X1 U9121 ( .A(n605), .B(n2431), .S(n2467), .Z(n1715) );
  MUX2_X1 U9122 ( .A(n606), .B(n2432), .S(n2467), .Z(n1714) );
  MUX2_X1 U9123 ( .A(n607), .B(n2433), .S(n2467), .Z(n1713) );
  MUX2_X1 U9124 ( .A(n608), .B(n2434), .S(n2467), .Z(n1712) );
  MUX2_X1 U9125 ( .A(n609), .B(n2435), .S(n2467), .Z(n1711) );
  MUX2_X1 U9126 ( .A(n610), .B(n2436), .S(n2467), .Z(n1710) );
  MUX2_X1 U9127 ( .A(n130), .B(n2437), .S(n2467), .Z(n1709) );
  MUX2_X1 U9128 ( .A(n134), .B(n2438), .S(n2467), .Z(n1708) );
  MUX2_X1 U9129 ( .A(n138), .B(n2439), .S(n2467), .Z(n1707) );
  MUX2_X1 U9130 ( .A(n142), .B(n2440), .S(n2467), .Z(n1706) );
  MUX2_X1 U9131 ( .A(n146), .B(n2441), .S(n2467), .Z(n1705) );
  MUX2_X1 U9132 ( .A(n150), .B(n2442), .S(n2467), .Z(n1704) );
  MUX2_X1 U9133 ( .A(n154), .B(n2443), .S(n2467), .Z(n1703) );
  MUX2_X1 U9134 ( .A(n158), .B(n2444), .S(n2467), .Z(n1702) );
  AND2_X1 U9135 ( .A1(n2449), .A2(n2468), .ZN(n2464) );
  AND3_X1 U9136 ( .A1(EN), .A2(n2469), .A3(WM), .ZN(n2449) );
  MUX2_X1 U9137 ( .A(n611), .B(n2412), .S(n2470), .Z(n1701) );
  MUX2_X1 U9138 ( .A(n612), .B(n2414), .S(n2470), .Z(n1700) );
  MUX2_X1 U9139 ( .A(n613), .B(n2415), .S(n2470), .Z(n1699) );
  MUX2_X1 U9140 ( .A(n614), .B(n2416), .S(n2470), .Z(n1698) );
  MUX2_X1 U9141 ( .A(n615), .B(n2417), .S(n2470), .Z(n1697) );
  MUX2_X1 U9142 ( .A(n616), .B(n2418), .S(n2470), .Z(n1696) );
  MUX2_X1 U9143 ( .A(n617), .B(n2419), .S(n2470), .Z(n1695) );
  MUX2_X1 U9144 ( .A(n618), .B(n2420), .S(n2470), .Z(n1694) );
  MUX2_X1 U9145 ( .A(n619), .B(n2421), .S(n2470), .Z(n1693) );
  MUX2_X1 U9146 ( .A(n620), .B(n2422), .S(n2470), .Z(n1692) );
  MUX2_X1 U9147 ( .A(n621), .B(n2423), .S(n2470), .Z(n1691) );
  MUX2_X1 U9148 ( .A(n622), .B(n2424), .S(n2470), .Z(n1690) );
  MUX2_X1 U9149 ( .A(n623), .B(n2425), .S(n2470), .Z(n1689) );
  MUX2_X1 U9150 ( .A(n624), .B(n2426), .S(n2470), .Z(n1688) );
  MUX2_X1 U9151 ( .A(n625), .B(n2427), .S(n2470), .Z(n1687) );
  MUX2_X1 U9152 ( .A(n626), .B(n2428), .S(n2470), .Z(n1686) );
  MUX2_X1 U9153 ( .A(n125), .B(n2429), .S(n2470), .Z(n1685) );
  MUX2_X1 U9154 ( .A(n2936), .B(n2430), .S(n2470), .Z(n1684) );
  MUX2_X1 U9155 ( .A(n2942), .B(n2431), .S(n2470), .Z(n1683) );
  MUX2_X1 U9156 ( .A(n2948), .B(n2432), .S(n2470), .Z(n1682) );
  MUX2_X1 U9157 ( .A(n2954), .B(n2433), .S(n2470), .Z(n1681) );
  MUX2_X1 U9158 ( .A(n2960), .B(n2434), .S(n2470), .Z(n1680) );
  MUX2_X1 U9159 ( .A(n2966), .B(n2435), .S(n2470), .Z(n1679) );
  MUX2_X1 U9160 ( .A(n2972), .B(n2436), .S(n2470), .Z(n1678) );
  MUX2_X1 U9161 ( .A(n909), .B(n2437), .S(n2470), .Z(n1677) );
  MUX2_X1 U9162 ( .A(n910), .B(n2438), .S(n2470), .Z(n1676) );
  MUX2_X1 U9163 ( .A(n911), .B(n2439), .S(n2470), .Z(n1675) );
  MUX2_X1 U9164 ( .A(n912), .B(n2440), .S(n2470), .Z(n1674) );
  MUX2_X1 U9165 ( .A(n913), .B(n2441), .S(n2470), .Z(n1673) );
  MUX2_X1 U9166 ( .A(n914), .B(n2442), .S(n2470), .Z(n1672) );
  MUX2_X1 U9167 ( .A(n915), .B(n2443), .S(n2470), .Z(n1671) );
  MUX2_X1 U9168 ( .A(n916), .B(n2444), .S(n2470), .Z(n1670) );
  MUX2_X1 U9169 ( .A(n341), .B(n2412), .S(n2472), .Z(n1669) );
  MUX2_X1 U9170 ( .A(n342), .B(n2414), .S(n2472), .Z(n1668) );
  MUX2_X1 U9171 ( .A(n343), .B(n2415), .S(n2472), .Z(n1667) );
  MUX2_X1 U9172 ( .A(n344), .B(n2416), .S(n2472), .Z(n1666) );
  MUX2_X1 U9173 ( .A(n345), .B(n2417), .S(n2472), .Z(n1665) );
  MUX2_X1 U9174 ( .A(n346), .B(n2418), .S(n2472), .Z(n1664) );
  MUX2_X1 U9175 ( .A(n347), .B(n2419), .S(n2472), .Z(n1663) );
  MUX2_X1 U9176 ( .A(n348), .B(n2420), .S(n2472), .Z(n1662) );
  MUX2_X1 U9177 ( .A(n349), .B(n2421), .S(n2472), .Z(n1661) );
  MUX2_X1 U9178 ( .A(n350), .B(n2422), .S(n2472), .Z(n1660) );
  MUX2_X1 U9179 ( .A(n351), .B(n2423), .S(n2472), .Z(n1659) );
  MUX2_X1 U9180 ( .A(n352), .B(n2424), .S(n2472), .Z(n1658) );
  MUX2_X1 U9181 ( .A(n353), .B(n2425), .S(n2472), .Z(n1657) );
  MUX2_X1 U9182 ( .A(n354), .B(n2426), .S(n2472), .Z(n1656) );
  MUX2_X1 U9183 ( .A(n355), .B(n2427), .S(n2472), .Z(n1655) );
  MUX2_X1 U9184 ( .A(n356), .B(n2428), .S(n2472), .Z(n1654) );
  MUX2_X1 U9185 ( .A(n123), .B(n2429), .S(n2472), .Z(n1653) );
  MUX2_X1 U9186 ( .A(n2935), .B(n2430), .S(n2472), .Z(n1652) );
  MUX2_X1 U9187 ( .A(n2941), .B(n2431), .S(n2472), .Z(n1651) );
  MUX2_X1 U9188 ( .A(n2947), .B(n2432), .S(n2472), .Z(n1650) );
  MUX2_X1 U9189 ( .A(n2953), .B(n2433), .S(n2472), .Z(n1649) );
  MUX2_X1 U9190 ( .A(n2959), .B(n2434), .S(n2472), .Z(n1648) );
  MUX2_X1 U9191 ( .A(n2965), .B(n2435), .S(n2472), .Z(n1647) );
  MUX2_X1 U9192 ( .A(n2971), .B(n2436), .S(n2472), .Z(n1646) );
  MUX2_X1 U9193 ( .A(n789), .B(n2437), .S(n2472), .Z(n1645) );
  MUX2_X1 U9194 ( .A(n790), .B(n2438), .S(n2472), .Z(n1644) );
  MUX2_X1 U9195 ( .A(n791), .B(n2439), .S(n2472), .Z(n1643) );
  MUX2_X1 U9196 ( .A(n792), .B(n2440), .S(n2472), .Z(n1642) );
  MUX2_X1 U9197 ( .A(n793), .B(n2441), .S(n2472), .Z(n1641) );
  MUX2_X1 U9198 ( .A(n794), .B(n2442), .S(n2472), .Z(n1640) );
  MUX2_X1 U9199 ( .A(n795), .B(n2443), .S(n2472), .Z(n1639) );
  MUX2_X1 U9200 ( .A(n796), .B(n2444), .S(n2472), .Z(n1638) );
  MUX2_X1 U9201 ( .A(n487), .B(n2412), .S(n2473), .Z(n1637) );
  MUX2_X1 U9202 ( .A(n488), .B(n2414), .S(n2473), .Z(n1636) );
  MUX2_X1 U9203 ( .A(n489), .B(n2415), .S(n2473), .Z(n1635) );
  MUX2_X1 U9204 ( .A(n490), .B(n2416), .S(n2473), .Z(n1634) );
  MUX2_X1 U9205 ( .A(n491), .B(n2417), .S(n2473), .Z(n1633) );
  MUX2_X1 U9206 ( .A(n492), .B(n2418), .S(n2473), .Z(n1632) );
  MUX2_X1 U9207 ( .A(n493), .B(n2419), .S(n2473), .Z(n1631) );
  MUX2_X1 U9208 ( .A(n494), .B(n2420), .S(n2473), .Z(n1630) );
  MUX2_X1 U9209 ( .A(n495), .B(n2421), .S(n2473), .Z(n1629) );
  MUX2_X1 U9210 ( .A(n496), .B(n2422), .S(n2473), .Z(n1628) );
  MUX2_X1 U9211 ( .A(n497), .B(n2423), .S(n2473), .Z(n1627) );
  MUX2_X1 U9212 ( .A(n498), .B(n2424), .S(n2473), .Z(n1626) );
  MUX2_X1 U9213 ( .A(n499), .B(n2425), .S(n2473), .Z(n1625) );
  MUX2_X1 U9214 ( .A(n500), .B(n2426), .S(n2473), .Z(n1624) );
  MUX2_X1 U9215 ( .A(n501), .B(n2427), .S(n2473), .Z(n1623) );
  MUX2_X1 U9216 ( .A(n502), .B(n2428), .S(n2473), .Z(n1622) );
  MUX2_X1 U9217 ( .A(n121), .B(n2429), .S(n2473), .Z(n1621) );
  MUX2_X1 U9218 ( .A(n17), .B(n2430), .S(n2473), .Z(n1620) );
  MUX2_X1 U9219 ( .A(n25), .B(n2431), .S(n2473), .Z(n1619) );
  MUX2_X1 U9220 ( .A(n33), .B(n2432), .S(n2473), .Z(n1618) );
  MUX2_X1 U9221 ( .A(n41), .B(n2433), .S(n2473), .Z(n1617) );
  MUX2_X1 U9222 ( .A(n49), .B(n2434), .S(n2473), .Z(n1616) );
  MUX2_X1 U9223 ( .A(n57), .B(n2435), .S(n2473), .Z(n1615) );
  MUX2_X1 U9224 ( .A(n65), .B(n2436), .S(n2473), .Z(n1614) );
  MUX2_X1 U9225 ( .A(n2980), .B(n2437), .S(n2473), .Z(n1613) );
  MUX2_X1 U9226 ( .A(n2988), .B(n2438), .S(n2473), .Z(n1612) );
  MUX2_X1 U9227 ( .A(n2996), .B(n2439), .S(n2473), .Z(n1611) );
  MUX2_X1 U9228 ( .A(n3004), .B(n2440), .S(n2473), .Z(n1610) );
  MUX2_X1 U9229 ( .A(n3012), .B(n2441), .S(n2473), .Z(n1609) );
  MUX2_X1 U9230 ( .A(n3020), .B(n2442), .S(n2473), .Z(n1608) );
  MUX2_X1 U9231 ( .A(n3028), .B(n2443), .S(n2473), .Z(n1607) );
  MUX2_X1 U9232 ( .A(n3036), .B(n2444), .S(n2473), .Z(n1606) );
  MUX2_X1 U9233 ( .A(n627), .B(n2412), .S(n2474), .Z(n1605) );
  MUX2_X1 U9234 ( .A(n628), .B(n2414), .S(n2474), .Z(n1604) );
  MUX2_X1 U9235 ( .A(n629), .B(n2415), .S(n2474), .Z(n1603) );
  MUX2_X1 U9236 ( .A(n630), .B(n2416), .S(n2474), .Z(n1602) );
  MUX2_X1 U9237 ( .A(n631), .B(n2417), .S(n2474), .Z(n1601) );
  MUX2_X1 U9238 ( .A(n632), .B(n2418), .S(n2474), .Z(n1600) );
  MUX2_X1 U9239 ( .A(n633), .B(n2419), .S(n2474), .Z(n1599) );
  MUX2_X1 U9240 ( .A(n634), .B(n2420), .S(n2474), .Z(n1598) );
  MUX2_X1 U9241 ( .A(n635), .B(n2421), .S(n2474), .Z(n1597) );
  MUX2_X1 U9242 ( .A(n636), .B(n2422), .S(n2474), .Z(n1596) );
  MUX2_X1 U9243 ( .A(n637), .B(n2423), .S(n2474), .Z(n1595) );
  MUX2_X1 U9244 ( .A(n638), .B(n2424), .S(n2474), .Z(n1594) );
  MUX2_X1 U9245 ( .A(n639), .B(n2425), .S(n2474), .Z(n1593) );
  MUX2_X1 U9246 ( .A(n640), .B(n2426), .S(n2474), .Z(n1592) );
  MUX2_X1 U9247 ( .A(n641), .B(n2427), .S(n2474), .Z(n1591) );
  MUX2_X1 U9248 ( .A(n642), .B(n2428), .S(n2474), .Z(n1590) );
  MUX2_X1 U9249 ( .A(n127), .B(n2429), .S(n2474), .Z(n1589) );
  MUX2_X1 U9250 ( .A(n253), .B(n2430), .S(n2474), .Z(n1588) );
  MUX2_X1 U9251 ( .A(n261), .B(n2431), .S(n2474), .Z(n1587) );
  MUX2_X1 U9252 ( .A(n269), .B(n2432), .S(n2474), .Z(n1586) );
  MUX2_X1 U9253 ( .A(n277), .B(n2433), .S(n2474), .Z(n1585) );
  MUX2_X1 U9254 ( .A(n285), .B(n2434), .S(n2474), .Z(n1584) );
  MUX2_X1 U9255 ( .A(n293), .B(n2435), .S(n2474), .Z(n1583) );
  MUX2_X1 U9256 ( .A(n301), .B(n2436), .S(n2474), .Z(n1582) );
  MUX2_X1 U9257 ( .A(n2979), .B(n2437), .S(n2474), .Z(n1581) );
  MUX2_X1 U9258 ( .A(n2987), .B(n2438), .S(n2474), .Z(n1580) );
  MUX2_X1 U9259 ( .A(n2995), .B(n2439), .S(n2474), .Z(n1579) );
  MUX2_X1 U9260 ( .A(n3003), .B(n2440), .S(n2474), .Z(n1578) );
  MUX2_X1 U9261 ( .A(n3011), .B(n2441), .S(n2474), .Z(n1577) );
  MUX2_X1 U9262 ( .A(n3019), .B(n2442), .S(n2474), .Z(n1576) );
  MUX2_X1 U9263 ( .A(n3027), .B(n2443), .S(n2474), .Z(n1575) );
  MUX2_X1 U9264 ( .A(n3035), .B(n2444), .S(n2474), .Z(n1574) );
  AND2_X1 U9265 ( .A1(n2475), .A2(n2450), .ZN(n2471) );
  MUX2_X1 U9266 ( .A(n643), .B(n2412), .S(n2476), .Z(n1573) );
  MUX2_X1 U9267 ( .A(n644), .B(n2414), .S(n2476), .Z(n1572) );
  MUX2_X1 U9268 ( .A(n645), .B(n2415), .S(n2476), .Z(n1571) );
  MUX2_X1 U9269 ( .A(n646), .B(n2416), .S(n2476), .Z(n1570) );
  MUX2_X1 U9270 ( .A(n647), .B(n2417), .S(n2476), .Z(n1569) );
  MUX2_X1 U9271 ( .A(n648), .B(n2418), .S(n2476), .Z(n1568) );
  MUX2_X1 U9272 ( .A(n649), .B(n2419), .S(n2476), .Z(n1567) );
  MUX2_X1 U9273 ( .A(n650), .B(n2420), .S(n2476), .Z(n1566) );
  MUX2_X1 U9274 ( .A(n651), .B(n2421), .S(n2476), .Z(n1565) );
  MUX2_X1 U9275 ( .A(n652), .B(n2422), .S(n2476), .Z(n1564) );
  MUX2_X1 U9276 ( .A(n653), .B(n2423), .S(n2476), .Z(n1563) );
  MUX2_X1 U9277 ( .A(n654), .B(n2424), .S(n2476), .Z(n1562) );
  MUX2_X1 U9278 ( .A(n655), .B(n2425), .S(n2476), .Z(n1561) );
  MUX2_X1 U9279 ( .A(n656), .B(n2426), .S(n2476), .Z(n1560) );
  MUX2_X1 U9280 ( .A(n657), .B(n2427), .S(n2476), .Z(n1559) );
  MUX2_X1 U9281 ( .A(n658), .B(n2428), .S(n2476), .Z(n1558) );
  MUX2_X1 U9282 ( .A(n361), .B(n2429), .S(n2476), .Z(n1557) );
  MUX2_X1 U9283 ( .A(n2934), .B(n2430), .S(n2476), .Z(n1556) );
  MUX2_X1 U9284 ( .A(n2940), .B(n2431), .S(n2476), .Z(n1555) );
  MUX2_X1 U9285 ( .A(n2946), .B(n2432), .S(n2476), .Z(n1554) );
  MUX2_X1 U9286 ( .A(n2952), .B(n2433), .S(n2476), .Z(n1553) );
  MUX2_X1 U9287 ( .A(n2958), .B(n2434), .S(n2476), .Z(n1552) );
  MUX2_X1 U9288 ( .A(n2964), .B(n2435), .S(n2476), .Z(n1551) );
  MUX2_X1 U9289 ( .A(n2970), .B(n2436), .S(n2476), .Z(n1550) );
  MUX2_X1 U9290 ( .A(n917), .B(n2437), .S(n2476), .Z(n1549) );
  MUX2_X1 U9291 ( .A(n918), .B(n2438), .S(n2476), .Z(n1548) );
  MUX2_X1 U9292 ( .A(n919), .B(n2439), .S(n2476), .Z(n1547) );
  MUX2_X1 U9293 ( .A(n920), .B(n2440), .S(n2476), .Z(n1546) );
  MUX2_X1 U9294 ( .A(n921), .B(n2441), .S(n2476), .Z(n1545) );
  MUX2_X1 U9295 ( .A(n922), .B(n2442), .S(n2476), .Z(n1544) );
  MUX2_X1 U9296 ( .A(n923), .B(n2443), .S(n2476), .Z(n1543) );
  MUX2_X1 U9297 ( .A(n924), .B(n2444), .S(n2476), .Z(n1542) );
  MUX2_X1 U9298 ( .A(n503), .B(n2412), .S(n2478), .Z(n1541) );
  MUX2_X1 U9299 ( .A(n504), .B(n2414), .S(n2478), .Z(n1540) );
  MUX2_X1 U9300 ( .A(n505), .B(n2415), .S(n2478), .Z(n1539) );
  MUX2_X1 U9301 ( .A(n506), .B(n2416), .S(n2478), .Z(n1538) );
  MUX2_X1 U9302 ( .A(n507), .B(n2417), .S(n2478), .Z(n1537) );
  MUX2_X1 U9303 ( .A(n508), .B(n2418), .S(n2478), .Z(n1536) );
  MUX2_X1 U9304 ( .A(n509), .B(n2419), .S(n2478), .Z(n1535) );
  MUX2_X1 U9305 ( .A(n510), .B(n2420), .S(n2478), .Z(n1534) );
  MUX2_X1 U9306 ( .A(n511), .B(n2421), .S(n2478), .Z(n1533) );
  MUX2_X1 U9307 ( .A(n512), .B(n2422), .S(n2478), .Z(n1532) );
  MUX2_X1 U9308 ( .A(n513), .B(n2423), .S(n2478), .Z(n1531) );
  MUX2_X1 U9309 ( .A(n514), .B(n2424), .S(n2478), .Z(n1530) );
  MUX2_X1 U9310 ( .A(n515), .B(n2425), .S(n2478), .Z(n1529) );
  MUX2_X1 U9311 ( .A(n516), .B(n2426), .S(n2478), .Z(n1528) );
  MUX2_X1 U9312 ( .A(n517), .B(n2427), .S(n2478), .Z(n1527) );
  MUX2_X1 U9313 ( .A(n518), .B(n2428), .S(n2478), .Z(n1526) );
  MUX2_X1 U9314 ( .A(n359), .B(n2429), .S(n2478), .Z(n1525) );
  MUX2_X1 U9315 ( .A(n2933), .B(n2430), .S(n2478), .Z(n1524) );
  MUX2_X1 U9316 ( .A(n2939), .B(n2431), .S(n2478), .Z(n1523) );
  MUX2_X1 U9317 ( .A(n2945), .B(n2432), .S(n2478), .Z(n1522) );
  MUX2_X1 U9318 ( .A(n2951), .B(n2433), .S(n2478), .Z(n1521) );
  MUX2_X1 U9319 ( .A(n2957), .B(n2434), .S(n2478), .Z(n1520) );
  MUX2_X1 U9320 ( .A(n2963), .B(n2435), .S(n2478), .Z(n1519) );
  MUX2_X1 U9321 ( .A(n2969), .B(n2436), .S(n2478), .Z(n1518) );
  MUX2_X1 U9322 ( .A(n797), .B(n2437), .S(n2478), .Z(n1517) );
  MUX2_X1 U9323 ( .A(n798), .B(n2438), .S(n2478), .Z(n1516) );
  MUX2_X1 U9324 ( .A(n799), .B(n2439), .S(n2478), .Z(n1515) );
  MUX2_X1 U9325 ( .A(n800), .B(n2440), .S(n2478), .Z(n1514) );
  MUX2_X1 U9326 ( .A(n801), .B(n2441), .S(n2478), .Z(n1513) );
  MUX2_X1 U9327 ( .A(n802), .B(n2442), .S(n2478), .Z(n1512) );
  MUX2_X1 U9328 ( .A(n803), .B(n2443), .S(n2478), .Z(n1511) );
  MUX2_X1 U9329 ( .A(n804), .B(n2444), .S(n2478), .Z(n1510) );
  MUX2_X1 U9330 ( .A(n519), .B(n2412), .S(n2479), .Z(n1509) );
  MUX2_X1 U9331 ( .A(n520), .B(n2414), .S(n2479), .Z(n1508) );
  MUX2_X1 U9332 ( .A(n521), .B(n2415), .S(n2479), .Z(n1507) );
  MUX2_X1 U9333 ( .A(n522), .B(n2416), .S(n2479), .Z(n1506) );
  MUX2_X1 U9334 ( .A(n523), .B(n2417), .S(n2479), .Z(n1505) );
  MUX2_X1 U9335 ( .A(n524), .B(n2418), .S(n2479), .Z(n1504) );
  MUX2_X1 U9336 ( .A(n525), .B(n2419), .S(n2479), .Z(n1503) );
  MUX2_X1 U9337 ( .A(n526), .B(n2420), .S(n2479), .Z(n1502) );
  MUX2_X1 U9338 ( .A(n527), .B(n2421), .S(n2479), .Z(n1501) );
  MUX2_X1 U9339 ( .A(n528), .B(n2422), .S(n2479), .Z(n1500) );
  MUX2_X1 U9340 ( .A(n529), .B(n2423), .S(n2479), .Z(n1499) );
  MUX2_X1 U9341 ( .A(n530), .B(n2424), .S(n2479), .Z(n1498) );
  MUX2_X1 U9342 ( .A(n531), .B(n2425), .S(n2479), .Z(n1497) );
  MUX2_X1 U9343 ( .A(n532), .B(n2426), .S(n2479), .Z(n1496) );
  MUX2_X1 U9344 ( .A(n533), .B(n2427), .S(n2479), .Z(n1495) );
  MUX2_X1 U9345 ( .A(n534), .B(n2428), .S(n2479), .Z(n1494) );
  MUX2_X1 U9346 ( .A(n357), .B(n2429), .S(n2479), .Z(n1493) );
  MUX2_X1 U9347 ( .A(n18), .B(n2430), .S(n2479), .Z(n1492) );
  MUX2_X1 U9348 ( .A(n26), .B(n2431), .S(n2479), .Z(n1491) );
  MUX2_X1 U9349 ( .A(n34), .B(n2432), .S(n2479), .Z(n1490) );
  MUX2_X1 U9350 ( .A(n42), .B(n2433), .S(n2479), .Z(n1489) );
  MUX2_X1 U9351 ( .A(n50), .B(n2434), .S(n2479), .Z(n1488) );
  MUX2_X1 U9352 ( .A(n58), .B(n2435), .S(n2479), .Z(n1487) );
  MUX2_X1 U9353 ( .A(n66), .B(n2436), .S(n2479), .Z(n1486) );
  MUX2_X1 U9354 ( .A(n2982), .B(n2437), .S(n2479), .Z(n1485) );
  MUX2_X1 U9355 ( .A(n2990), .B(n2438), .S(n2479), .Z(n1484) );
  MUX2_X1 U9356 ( .A(n2998), .B(n2439), .S(n2479), .Z(n1483) );
  MUX2_X1 U9357 ( .A(n3006), .B(n2440), .S(n2479), .Z(n1482) );
  MUX2_X1 U9358 ( .A(n3014), .B(n2441), .S(n2479), .Z(n1481) );
  MUX2_X1 U9359 ( .A(n3022), .B(n2442), .S(n2479), .Z(n1480) );
  MUX2_X1 U9360 ( .A(n3030), .B(n2443), .S(n2479), .Z(n1479) );
  MUX2_X1 U9361 ( .A(n3038), .B(n2444), .S(n2479), .Z(n1478) );
  MUX2_X1 U9362 ( .A(n659), .B(n2412), .S(n2480), .Z(n1477) );
  MUX2_X1 U9363 ( .A(n660), .B(n2414), .S(n2480), .Z(n1476) );
  MUX2_X1 U9364 ( .A(n661), .B(n2415), .S(n2480), .Z(n1475) );
  MUX2_X1 U9365 ( .A(n662), .B(n2416), .S(n2480), .Z(n1474) );
  MUX2_X1 U9366 ( .A(n663), .B(n2417), .S(n2480), .Z(n1473) );
  MUX2_X1 U9367 ( .A(n664), .B(n2418), .S(n2480), .Z(n1472) );
  MUX2_X1 U9368 ( .A(n665), .B(n2419), .S(n2480), .Z(n1471) );
  MUX2_X1 U9369 ( .A(n666), .B(n2420), .S(n2480), .Z(n1470) );
  MUX2_X1 U9370 ( .A(n667), .B(n2421), .S(n2480), .Z(n1469) );
  MUX2_X1 U9371 ( .A(n668), .B(n2422), .S(n2480), .Z(n1468) );
  MUX2_X1 U9372 ( .A(n669), .B(n2423), .S(n2480), .Z(n1467) );
  MUX2_X1 U9373 ( .A(n670), .B(n2424), .S(n2480), .Z(n1466) );
  MUX2_X1 U9374 ( .A(n671), .B(n2425), .S(n2480), .Z(n1465) );
  MUX2_X1 U9375 ( .A(n672), .B(n2426), .S(n2480), .Z(n1464) );
  MUX2_X1 U9376 ( .A(n673), .B(n2427), .S(n2480), .Z(n1463) );
  MUX2_X1 U9377 ( .A(n674), .B(n2428), .S(n2480), .Z(n1462) );
  MUX2_X1 U9378 ( .A(n363), .B(n2429), .S(n2480), .Z(n1461) );
  MUX2_X1 U9379 ( .A(n254), .B(n2430), .S(n2480), .Z(n1460) );
  MUX2_X1 U9380 ( .A(n262), .B(n2431), .S(n2480), .Z(n1459) );
  MUX2_X1 U9381 ( .A(n270), .B(n2432), .S(n2480), .Z(n1458) );
  MUX2_X1 U9382 ( .A(n278), .B(n2433), .S(n2480), .Z(n1457) );
  MUX2_X1 U9383 ( .A(n286), .B(n2434), .S(n2480), .Z(n1456) );
  MUX2_X1 U9384 ( .A(n294), .B(n2435), .S(n2480), .Z(n1455) );
  MUX2_X1 U9385 ( .A(n302), .B(n2436), .S(n2480), .Z(n1454) );
  MUX2_X1 U9386 ( .A(n2981), .B(n2437), .S(n2480), .Z(n1453) );
  MUX2_X1 U9387 ( .A(n2989), .B(n2438), .S(n2480), .Z(n1452) );
  MUX2_X1 U9388 ( .A(n2997), .B(n2439), .S(n2480), .Z(n1451) );
  MUX2_X1 U9389 ( .A(n3005), .B(n2440), .S(n2480), .Z(n1450) );
  MUX2_X1 U9390 ( .A(n3013), .B(n2441), .S(n2480), .Z(n1449) );
  MUX2_X1 U9391 ( .A(n3021), .B(n2442), .S(n2480), .Z(n1448) );
  MUX2_X1 U9392 ( .A(n3029), .B(n2443), .S(n2480), .Z(n1447) );
  MUX2_X1 U9393 ( .A(n3037), .B(n2444), .S(n2480), .Z(n1446) );
  AND2_X1 U9394 ( .A1(n2475), .A2(n2456), .ZN(n2477) );
  MUX2_X1 U9395 ( .A(n675), .B(n2412), .S(n2481), .Z(n1445) );
  MUX2_X1 U9396 ( .A(n676), .B(n2414), .S(n2481), .Z(n1444) );
  MUX2_X1 U9397 ( .A(n677), .B(n2415), .S(n2481), .Z(n1443) );
  MUX2_X1 U9398 ( .A(n678), .B(n2416), .S(n2481), .Z(n1442) );
  MUX2_X1 U9399 ( .A(n679), .B(n2417), .S(n2481), .Z(n1441) );
  MUX2_X1 U9400 ( .A(n680), .B(n2418), .S(n2481), .Z(n1440) );
  MUX2_X1 U9401 ( .A(n681), .B(n2419), .S(n2481), .Z(n1439) );
  MUX2_X1 U9402 ( .A(n682), .B(n2420), .S(n2481), .Z(n1438) );
  MUX2_X1 U9403 ( .A(n683), .B(n2421), .S(n2481), .Z(n1437) );
  MUX2_X1 U9404 ( .A(n684), .B(n2422), .S(n2481), .Z(n1436) );
  MUX2_X1 U9405 ( .A(n685), .B(n2423), .S(n2481), .Z(n1435) );
  MUX2_X1 U9406 ( .A(n686), .B(n2424), .S(n2481), .Z(n1434) );
  MUX2_X1 U9407 ( .A(n687), .B(n2425), .S(n2481), .Z(n1433) );
  MUX2_X1 U9408 ( .A(n688), .B(n2426), .S(n2481), .Z(n1432) );
  MUX2_X1 U9409 ( .A(n689), .B(n2427), .S(n2481), .Z(n1431) );
  MUX2_X1 U9410 ( .A(n690), .B(n2428), .S(n2481), .Z(n1430) );
  MUX2_X1 U9411 ( .A(n925), .B(n2429), .S(n2481), .Z(n1429) );
  MUX2_X1 U9412 ( .A(n20), .B(n2430), .S(n2481), .Z(n1428) );
  MUX2_X1 U9413 ( .A(n28), .B(n2431), .S(n2481), .Z(n1427) );
  MUX2_X1 U9414 ( .A(n36), .B(n2432), .S(n2481), .Z(n1426) );
  MUX2_X1 U9415 ( .A(n44), .B(n2433), .S(n2481), .Z(n1425) );
  MUX2_X1 U9416 ( .A(n52), .B(n2434), .S(n2481), .Z(n1424) );
  MUX2_X1 U9417 ( .A(n60), .B(n2435), .S(n2481), .Z(n1423) );
  MUX2_X1 U9418 ( .A(n68), .B(n2436), .S(n2481), .Z(n1422) );
  MUX2_X1 U9419 ( .A(n926), .B(n2437), .S(n2481), .Z(n1421) );
  MUX2_X1 U9420 ( .A(n927), .B(n2438), .S(n2481), .Z(n1420) );
  MUX2_X1 U9421 ( .A(n928), .B(n2439), .S(n2481), .Z(n1419) );
  MUX2_X1 U9422 ( .A(n929), .B(n2440), .S(n2481), .Z(n1418) );
  MUX2_X1 U9423 ( .A(n930), .B(n2441), .S(n2481), .Z(n1417) );
  MUX2_X1 U9424 ( .A(n931), .B(n2442), .S(n2481), .Z(n1416) );
  MUX2_X1 U9425 ( .A(n932), .B(n2443), .S(n2481), .Z(n1415) );
  MUX2_X1 U9426 ( .A(n933), .B(n2444), .S(n2481), .Z(n1414) );
  MUX2_X1 U9427 ( .A(n535), .B(n2412), .S(n2483), .Z(n1413) );
  MUX2_X1 U9428 ( .A(n536), .B(n2414), .S(n2483), .Z(n1412) );
  MUX2_X1 U9429 ( .A(n537), .B(n2415), .S(n2483), .Z(n1411) );
  MUX2_X1 U9430 ( .A(n538), .B(n2416), .S(n2483), .Z(n1410) );
  MUX2_X1 U9431 ( .A(n539), .B(n2417), .S(n2483), .Z(n1409) );
  MUX2_X1 U9432 ( .A(n540), .B(n2418), .S(n2483), .Z(n1408) );
  MUX2_X1 U9433 ( .A(n541), .B(n2419), .S(n2483), .Z(n1407) );
  MUX2_X1 U9434 ( .A(n542), .B(n2420), .S(n2483), .Z(n1406) );
  MUX2_X1 U9435 ( .A(n543), .B(n2421), .S(n2483), .Z(n1405) );
  MUX2_X1 U9436 ( .A(n544), .B(n2422), .S(n2483), .Z(n1404) );
  MUX2_X1 U9437 ( .A(n545), .B(n2423), .S(n2483), .Z(n1403) );
  MUX2_X1 U9438 ( .A(n546), .B(n2424), .S(n2483), .Z(n1402) );
  MUX2_X1 U9439 ( .A(n547), .B(n2425), .S(n2483), .Z(n1401) );
  MUX2_X1 U9440 ( .A(n548), .B(n2426), .S(n2483), .Z(n1400) );
  MUX2_X1 U9441 ( .A(n549), .B(n2427), .S(n2483), .Z(n1399) );
  MUX2_X1 U9442 ( .A(n550), .B(n2428), .S(n2483), .Z(n1398) );
  MUX2_X1 U9443 ( .A(n934), .B(n2429), .S(n2483), .Z(n1397) );
  MUX2_X1 U9444 ( .A(n256), .B(n2430), .S(n2483), .Z(n1396) );
  MUX2_X1 U9445 ( .A(n264), .B(n2431), .S(n2483), .Z(n1395) );
  MUX2_X1 U9446 ( .A(n272), .B(n2432), .S(n2483), .Z(n1394) );
  MUX2_X1 U9447 ( .A(n280), .B(n2433), .S(n2483), .Z(n1393) );
  MUX2_X1 U9448 ( .A(n288), .B(n2434), .S(n2483), .Z(n1392) );
  MUX2_X1 U9449 ( .A(n296), .B(n2435), .S(n2483), .Z(n1391) );
  MUX2_X1 U9450 ( .A(n304), .B(n2436), .S(n2483), .Z(n1390) );
  MUX2_X1 U9451 ( .A(n805), .B(n2437), .S(n2483), .Z(n1389) );
  MUX2_X1 U9452 ( .A(n806), .B(n2438), .S(n2483), .Z(n1388) );
  MUX2_X1 U9453 ( .A(n807), .B(n2439), .S(n2483), .Z(n1387) );
  MUX2_X1 U9454 ( .A(n808), .B(n2440), .S(n2483), .Z(n1386) );
  MUX2_X1 U9455 ( .A(n809), .B(n2441), .S(n2483), .Z(n1385) );
  MUX2_X1 U9456 ( .A(n810), .B(n2442), .S(n2483), .Z(n1384) );
  MUX2_X1 U9457 ( .A(n811), .B(n2443), .S(n2483), .Z(n1383) );
  MUX2_X1 U9458 ( .A(n812), .B(n2444), .S(n2483), .Z(n1382) );
  MUX2_X1 U9459 ( .A(n551), .B(n2412), .S(n2484), .Z(n1381) );
  MUX2_X1 U9460 ( .A(n552), .B(n2414), .S(n2484), .Z(n1380) );
  MUX2_X1 U9461 ( .A(n553), .B(n2415), .S(n2484), .Z(n1379) );
  MUX2_X1 U9462 ( .A(n554), .B(n2416), .S(n2484), .Z(n1378) );
  MUX2_X1 U9463 ( .A(n555), .B(n2417), .S(n2484), .Z(n1377) );
  MUX2_X1 U9464 ( .A(n556), .B(n2418), .S(n2484), .Z(n1376) );
  MUX2_X1 U9465 ( .A(n557), .B(n2419), .S(n2484), .Z(n1375) );
  MUX2_X1 U9466 ( .A(n558), .B(n2420), .S(n2484), .Z(n1374) );
  MUX2_X1 U9467 ( .A(n559), .B(n2421), .S(n2484), .Z(n1373) );
  MUX2_X1 U9468 ( .A(n560), .B(n2422), .S(n2484), .Z(n1372) );
  MUX2_X1 U9469 ( .A(n561), .B(n2423), .S(n2484), .Z(n1371) );
  MUX2_X1 U9470 ( .A(n562), .B(n2424), .S(n2484), .Z(n1370) );
  MUX2_X1 U9471 ( .A(n563), .B(n2425), .S(n2484), .Z(n1369) );
  INV_X1 U9472 ( .A(Rst), .ZN(n13687) );
  MUX2_X1 U9473 ( .A(n564), .B(n2426), .S(n2484), .Z(n1368) );
  MUX2_X1 U9474 ( .A(n565), .B(n2427), .S(n2484), .Z(n1367) );
  MUX2_X1 U9475 ( .A(n566), .B(n2428), .S(n2484), .Z(n1366) );
  MUX2_X1 U9476 ( .A(n935), .B(n2429), .S(n2484), .Z(n1365) );
  MUX2_X1 U9477 ( .A(n567), .B(n2430), .S(n2484), .Z(n1364) );
  MUX2_X1 U9478 ( .A(n568), .B(n2431), .S(n2484), .Z(n1363) );
  MUX2_X1 U9479 ( .A(n569), .B(n2432), .S(n2484), .Z(n1362) );
  MUX2_X1 U9480 ( .A(n570), .B(n2433), .S(n2484), .Z(n1361) );
  MUX2_X1 U9481 ( .A(n571), .B(n2434), .S(n2484), .Z(n1360) );
  MUX2_X1 U9482 ( .A(n572), .B(n2435), .S(n2484), .Z(n1359) );
  MUX2_X1 U9483 ( .A(n573), .B(n2436), .S(n2484), .Z(n1358) );
  MUX2_X1 U9484 ( .A(n367), .B(n2437), .S(n2484), .Z(n1357) );
  MUX2_X1 U9485 ( .A(n371), .B(n2438), .S(n2484), .Z(n1356) );
  MUX2_X1 U9486 ( .A(n375), .B(n2439), .S(n2484), .Z(n1355) );
  MUX2_X1 U9487 ( .A(n379), .B(n2440), .S(n2484), .Z(n1354) );
  MUX2_X1 U9488 ( .A(n383), .B(n2441), .S(n2484), .Z(n1353) );
  MUX2_X1 U9489 ( .A(n387), .B(n2442), .S(n2484), .Z(n1352) );
  MUX2_X1 U9490 ( .A(n391), .B(n2443), .S(n2484), .Z(n1351) );
  MUX2_X1 U9491 ( .A(n395), .B(n2444), .S(n2484), .Z(n1350) );
  MUX2_X1 U9492 ( .A(n221), .B(n2412), .S(n2485), .Z(n1349) );
  MUX2_X1 U9493 ( .A(n222), .B(n2414), .S(n2485), .Z(n1348) );
  MUX2_X1 U9494 ( .A(n223), .B(n2415), .S(n2485), .Z(n1347) );
  MUX2_X1 U9495 ( .A(n224), .B(n2416), .S(n2485), .Z(n1346) );
  MUX2_X1 U9496 ( .A(n225), .B(n2417), .S(n2485), .Z(n1345) );
  MUX2_X1 U9497 ( .A(n226), .B(n2418), .S(n2485), .Z(n1344) );
  MUX2_X1 U9498 ( .A(n227), .B(n2419), .S(n2485), .Z(n1343) );
  MUX2_X1 U9499 ( .A(n228), .B(n2420), .S(n2485), .Z(n1342) );
  MUX2_X1 U9500 ( .A(n229), .B(n2421), .S(n2485), .Z(n1341) );
  MUX2_X1 U9501 ( .A(n230), .B(n2422), .S(n2485), .Z(n1340) );
  MUX2_X1 U9502 ( .A(n231), .B(n2423), .S(n2485), .Z(n1339) );
  MUX2_X1 U9503 ( .A(n232), .B(n2424), .S(n2485), .Z(n1338) );
  MUX2_X1 U9504 ( .A(n233), .B(n2425), .S(n2485), .Z(n1337) );
  MUX2_X1 U9505 ( .A(n234), .B(n2426), .S(n2485), .Z(n1336) );
  MUX2_X1 U9506 ( .A(n235), .B(n2427), .S(n2485), .Z(n1335) );
  MUX2_X1 U9507 ( .A(n236), .B(n2428), .S(n2485), .Z(n1334) );
  MUX2_X1 U9508 ( .A(n936), .B(n2429), .S(n2485), .Z(n1333) );
  MUX2_X1 U9509 ( .A(n691), .B(n2430), .S(n2485), .Z(n1332) );
  MUX2_X1 U9510 ( .A(n692), .B(n2431), .S(n2485), .Z(n1331) );
  MUX2_X1 U9511 ( .A(n693), .B(n2432), .S(n2485), .Z(n1330) );
  MUX2_X1 U9512 ( .A(n694), .B(n2433), .S(n2485), .Z(n1329) );
  MUX2_X1 U9513 ( .A(n695), .B(n2434), .S(n2485), .Z(n1328) );
  MUX2_X1 U9514 ( .A(n696), .B(n2435), .S(n2485), .Z(n1327) );
  MUX2_X1 U9515 ( .A(n697), .B(n2436), .S(n2485), .Z(n1326) );
  MUX2_X1 U9516 ( .A(n131), .B(n2437), .S(n2485), .Z(n1325) );
  MUX2_X1 U9517 ( .A(n135), .B(n2438), .S(n2485), .Z(n1324) );
  MUX2_X1 U9518 ( .A(n139), .B(n2439), .S(n2485), .Z(n1323) );
  MUX2_X1 U9519 ( .A(n143), .B(n2440), .S(n2485), .Z(n1322) );
  MUX2_X1 U9520 ( .A(n147), .B(n2441), .S(n2485), .Z(n1321) );
  MUX2_X1 U9521 ( .A(n151), .B(n2442), .S(n2485), .Z(n1320) );
  MUX2_X1 U9522 ( .A(n155), .B(n2443), .S(n2485), .Z(n1319) );
  MUX2_X1 U9523 ( .A(n159), .B(n2444), .S(n2485), .Z(n1318) );
  AND2_X1 U9524 ( .A1(n2475), .A2(n2462), .ZN(n2482) );
  MUX2_X1 U9525 ( .A(n237), .B(n2412), .S(n2486), .Z(n1317) );
  MUX2_X1 U9526 ( .A(n238), .B(n2414), .S(n2486), .Z(n1316) );
  MUX2_X1 U9527 ( .A(n239), .B(n2415), .S(n2486), .Z(n1315) );
  MUX2_X1 U9528 ( .A(n240), .B(n2416), .S(n2486), .Z(n1314) );
  MUX2_X1 U9529 ( .A(n241), .B(n2417), .S(n2486), .Z(n1313) );
  MUX2_X1 U9530 ( .A(n242), .B(n2418), .S(n2486), .Z(n1312) );
  MUX2_X1 U9531 ( .A(n243), .B(n2419), .S(n2486), .Z(n1311) );
  MUX2_X1 U9532 ( .A(n244), .B(n2420), .S(n2486), .Z(n1310) );
  MUX2_X1 U9533 ( .A(n245), .B(n2421), .S(n2486), .Z(n1309) );
  MUX2_X1 U9534 ( .A(n246), .B(n2422), .S(n2486), .Z(n1308) );
  MUX2_X1 U9535 ( .A(n247), .B(n2423), .S(n2486), .Z(n1307) );
  MUX2_X1 U9536 ( .A(n248), .B(n2424), .S(n2486), .Z(n1306) );
  MUX2_X1 U9537 ( .A(n249), .B(n2425), .S(n2486), .Z(n1305) );
  MUX2_X1 U9538 ( .A(n250), .B(n2426), .S(n2486), .Z(n1304) );
  MUX2_X1 U9539 ( .A(n251), .B(n2427), .S(n2486), .Z(n1303) );
  MUX2_X1 U9540 ( .A(n252), .B(n2428), .S(n2486), .Z(n1302) );
  MUX2_X1 U9541 ( .A(n813), .B(n2429), .S(n2486), .Z(n1301) );
  MUX2_X1 U9542 ( .A(n19), .B(n2430), .S(n2486), .Z(n1300) );
  MUX2_X1 U9543 ( .A(n27), .B(n2431), .S(n2486), .Z(n1299) );
  MUX2_X1 U9544 ( .A(n35), .B(n2432), .S(n2486), .Z(n1298) );
  MUX2_X1 U9545 ( .A(n43), .B(n2433), .S(n2486), .Z(n1297) );
  MUX2_X1 U9546 ( .A(n51), .B(n2434), .S(n2486), .Z(n1296) );
  MUX2_X1 U9547 ( .A(n59), .B(n2435), .S(n2486), .Z(n1295) );
  MUX2_X1 U9548 ( .A(n67), .B(n2436), .S(n2486), .Z(n1294) );
  MUX2_X1 U9549 ( .A(n937), .B(n2437), .S(n2486), .Z(n1293) );
  MUX2_X1 U9550 ( .A(n938), .B(n2438), .S(n2486), .Z(n1292) );
  MUX2_X1 U9551 ( .A(n939), .B(n2439), .S(n2486), .Z(n1291) );
  MUX2_X1 U9552 ( .A(n940), .B(n2440), .S(n2486), .Z(n1290) );
  MUX2_X1 U9553 ( .A(n941), .B(n2441), .S(n2486), .Z(n1289) );
  MUX2_X1 U9554 ( .A(n942), .B(n2442), .S(n2486), .Z(n1288) );
  MUX2_X1 U9555 ( .A(n943), .B(n2443), .S(n2486), .Z(n1287) );
  MUX2_X1 U9556 ( .A(n944), .B(n2444), .S(n2486), .Z(n1286) );
  MUX2_X1 U9557 ( .A(n574), .B(n2412), .S(n2488), .Z(n1285) );
  MUX2_X1 U9558 ( .A(n575), .B(n2414), .S(n2488), .Z(n1284) );
  MUX2_X1 U9559 ( .A(n576), .B(n2415), .S(n2488), .Z(n1283) );
  MUX2_X1 U9560 ( .A(n577), .B(n2416), .S(n2488), .Z(n1282) );
  MUX2_X1 U9561 ( .A(n578), .B(n2417), .S(n2488), .Z(n1281) );
  MUX2_X1 U9562 ( .A(n579), .B(n2418), .S(n2488), .Z(n1280) );
  MUX2_X1 U9563 ( .A(n580), .B(n2419), .S(n2488), .Z(n1279) );
  MUX2_X1 U9564 ( .A(n581), .B(n2420), .S(n2488), .Z(n1278) );
  MUX2_X1 U9565 ( .A(n582), .B(n2421), .S(n2488), .Z(n1277) );
  MUX2_X1 U9566 ( .A(n583), .B(n2422), .S(n2488), .Z(n1276) );
  MUX2_X1 U9567 ( .A(n584), .B(n2423), .S(n2488), .Z(n1275) );
  MUX2_X1 U9568 ( .A(n585), .B(n2424), .S(n2488), .Z(n1274) );
  MUX2_X1 U9569 ( .A(n586), .B(n2425), .S(n2488), .Z(n1273) );
  MUX2_X1 U9570 ( .A(n587), .B(n2426), .S(n2488), .Z(n1272) );
  MUX2_X1 U9571 ( .A(n588), .B(n2427), .S(n2488), .Z(n1271) );
  MUX2_X1 U9572 ( .A(n589), .B(n2428), .S(n2488), .Z(n1270) );
  MUX2_X1 U9573 ( .A(n814), .B(n2429), .S(n2488), .Z(n1269) );
  MUX2_X1 U9574 ( .A(n255), .B(n2430), .S(n2488), .Z(n1268) );
  MUX2_X1 U9575 ( .A(n263), .B(n2431), .S(n2488), .Z(n1267) );
  MUX2_X1 U9576 ( .A(n271), .B(n2432), .S(n2488), .Z(n1266) );
  MUX2_X1 U9577 ( .A(n279), .B(n2433), .S(n2488), .Z(n1265) );
  MUX2_X1 U9578 ( .A(n287), .B(n2434), .S(n2488), .Z(n1264) );
  MUX2_X1 U9579 ( .A(n295), .B(n2435), .S(n2488), .Z(n1263) );
  MUX2_X1 U9580 ( .A(n303), .B(n2436), .S(n2488), .Z(n1262) );
  MUX2_X1 U9581 ( .A(n815), .B(n2437), .S(n2488), .Z(n1261) );
  MUX2_X1 U9582 ( .A(n816), .B(n2438), .S(n2488), .Z(n1260) );
  MUX2_X1 U9583 ( .A(n817), .B(n2439), .S(n2488), .Z(n1259) );
  MUX2_X1 U9584 ( .A(n818), .B(n2440), .S(n2488), .Z(n1258) );
  MUX2_X1 U9585 ( .A(n819), .B(n2441), .S(n2488), .Z(n1257) );
  MUX2_X1 U9586 ( .A(n820), .B(n2442), .S(n2488), .Z(n1256) );
  MUX2_X1 U9587 ( .A(n821), .B(n2443), .S(n2488), .Z(n1255) );
  MUX2_X1 U9588 ( .A(n822), .B(n2444), .S(n2488), .Z(n1254) );
  MUX2_X1 U9589 ( .A(n1), .B(n2412), .S(n2489), .Z(n1253) );
  MUX2_X1 U9590 ( .A(n2), .B(n2414), .S(n2489), .Z(n1252) );
  MUX2_X1 U9591 ( .A(n3), .B(n2415), .S(n2489), .Z(n1251) );
  MUX2_X1 U9592 ( .A(n4), .B(n2416), .S(n2489), .Z(n1250) );
  MUX2_X1 U9593 ( .A(n5), .B(n2417), .S(n2489), .Z(n1249) );
  MUX2_X1 U9594 ( .A(n6), .B(n2418), .S(n2489), .Z(n1248) );
  MUX2_X1 U9595 ( .A(n7), .B(n2419), .S(n2489), .Z(n1247) );
  MUX2_X1 U9596 ( .A(n8), .B(n2420), .S(n2489), .Z(n1246) );
  MUX2_X1 U9597 ( .A(n9), .B(n2421), .S(n2489), .Z(n1245) );
  MUX2_X1 U9598 ( .A(n10), .B(n2422), .S(n2489), .Z(n1244) );
  MUX2_X1 U9599 ( .A(n11), .B(n2423), .S(n2489), .Z(n1243) );
  MUX2_X1 U9600 ( .A(n12), .B(n2424), .S(n2489), .Z(n1242) );
  MUX2_X1 U9601 ( .A(n13), .B(n2425), .S(n2489), .Z(n1241) );
  MUX2_X1 U9602 ( .A(n14), .B(n2426), .S(n2489), .Z(n1240) );
  MUX2_X1 U9603 ( .A(n15), .B(n2427), .S(n2489), .Z(n1239) );
  MUX2_X1 U9604 ( .A(n16), .B(n2428), .S(n2489), .Z(n1238) );
  MUX2_X1 U9605 ( .A(n823), .B(n2429), .S(n2489), .Z(n1237) );
  MUX2_X1 U9606 ( .A(n590), .B(n2430), .S(n2489), .Z(n1236) );
  MUX2_X1 U9607 ( .A(n591), .B(n2431), .S(n2489), .Z(n1235) );
  MUX2_X1 U9608 ( .A(n592), .B(n2432), .S(n2489), .Z(n1234) );
  MUX2_X1 U9609 ( .A(n593), .B(n2433), .S(n2489), .Z(n1233) );
  MUX2_X1 U9610 ( .A(n594), .B(n2434), .S(n2489), .Z(n1232) );
  MUX2_X1 U9611 ( .A(n595), .B(n2435), .S(n2489), .Z(n1231) );
  MUX2_X1 U9612 ( .A(n596), .B(n2436), .S(n2489), .Z(n1230) );
  MUX2_X1 U9613 ( .A(n368), .B(n2437), .S(n2489), .Z(n1229) );
  MUX2_X1 U9614 ( .A(n372), .B(n2438), .S(n2489), .Z(n1228) );
  MUX2_X1 U9615 ( .A(n376), .B(n2439), .S(n2489), .Z(n1227) );
  MUX2_X1 U9616 ( .A(n380), .B(n2440), .S(n2489), .Z(n1226) );
  MUX2_X1 U9617 ( .A(n384), .B(n2441), .S(n2489), .Z(n1225) );
  MUX2_X1 U9618 ( .A(n388), .B(n2442), .S(n2489), .Z(n1224) );
  MUX2_X1 U9619 ( .A(n392), .B(n2443), .S(n2489), .Z(n1223) );
  MUX2_X1 U9620 ( .A(n396), .B(n2444), .S(n2489), .Z(n1222) );
  MUX2_X1 U9621 ( .A(n698), .B(n2412), .S(n2490), .Z(n1221) );
  INV_X1 U9622 ( .A(n2491), .ZN(n2412) );
  OAI21_X1 U9623 ( .B1(Din[31]), .B2(n2492), .A(n2493), .ZN(n2491) );
  MUX2_X1 U9624 ( .A(n699), .B(n2414), .S(n2490), .Z(n1220) );
  INV_X1 U9625 ( .A(n2494), .ZN(n2414) );
  OAI21_X1 U9626 ( .B1(Din[30]), .B2(n2492), .A(n2493), .ZN(n2494) );
  MUX2_X1 U9627 ( .A(n700), .B(n2415), .S(n2490), .Z(n1219) );
  INV_X1 U9628 ( .A(n2495), .ZN(n2415) );
  OAI21_X1 U9629 ( .B1(Din[29]), .B2(n2492), .A(n2493), .ZN(n2495) );
  MUX2_X1 U9630 ( .A(n701), .B(n2416), .S(n2490), .Z(n1218) );
  INV_X1 U9631 ( .A(n2496), .ZN(n2416) );
  OAI21_X1 U9632 ( .B1(Din[28]), .B2(n2492), .A(n2493), .ZN(n2496) );
  MUX2_X1 U9633 ( .A(n702), .B(n2417), .S(n2490), .Z(n1217) );
  INV_X1 U9634 ( .A(n2497), .ZN(n2417) );
  OAI21_X1 U9635 ( .B1(Din[27]), .B2(n2492), .A(n2493), .ZN(n2497) );
  MUX2_X1 U9636 ( .A(n703), .B(n2418), .S(n2490), .Z(n1216) );
  INV_X1 U9637 ( .A(n2498), .ZN(n2418) );
  OAI21_X1 U9638 ( .B1(Din[26]), .B2(n2492), .A(n2493), .ZN(n2498) );
  MUX2_X1 U9639 ( .A(n704), .B(n2419), .S(n2490), .Z(n1215) );
  INV_X1 U9640 ( .A(n2499), .ZN(n2419) );
  OAI21_X1 U9641 ( .B1(Din[25]), .B2(n2492), .A(n2493), .ZN(n2499) );
  MUX2_X1 U9642 ( .A(n705), .B(n2420), .S(n2490), .Z(n1214) );
  INV_X1 U9643 ( .A(n2500), .ZN(n2420) );
  OAI21_X1 U9644 ( .B1(Din[24]), .B2(n2492), .A(n2493), .ZN(n2500) );
  MUX2_X1 U9645 ( .A(n706), .B(n2421), .S(n2490), .Z(n1213) );
  INV_X1 U9646 ( .A(n2501), .ZN(n2421) );
  OAI21_X1 U9647 ( .B1(Din[23]), .B2(n2492), .A(n2493), .ZN(n2501) );
  MUX2_X1 U9648 ( .A(n707), .B(n2422), .S(n2490), .Z(n1212) );
  INV_X1 U9649 ( .A(n2502), .ZN(n2422) );
  OAI21_X1 U9650 ( .B1(Din[22]), .B2(n2492), .A(n2493), .ZN(n2502) );
  MUX2_X1 U9651 ( .A(n708), .B(n2423), .S(n2490), .Z(n1211) );
  INV_X1 U9652 ( .A(n2503), .ZN(n2423) );
  OAI21_X1 U9653 ( .B1(Din[21]), .B2(n2492), .A(n2493), .ZN(n2503) );
  MUX2_X1 U9654 ( .A(n709), .B(n2424), .S(n2490), .Z(n1210) );
  INV_X1 U9655 ( .A(n2504), .ZN(n2424) );
  OAI21_X1 U9656 ( .B1(Din[20]), .B2(n2492), .A(n2493), .ZN(n2504) );
  MUX2_X1 U9657 ( .A(n710), .B(n2425), .S(n2490), .Z(n1209) );
  INV_X1 U9658 ( .A(n2505), .ZN(n2425) );
  OAI21_X1 U9659 ( .B1(Din[19]), .B2(n2492), .A(n2493), .ZN(n2505) );
  MUX2_X1 U9660 ( .A(n711), .B(n2426), .S(n2490), .Z(n1208) );
  INV_X1 U9661 ( .A(n2506), .ZN(n2426) );
  OAI21_X1 U9662 ( .B1(Din[18]), .B2(n2492), .A(n2493), .ZN(n2506) );
  MUX2_X1 U9663 ( .A(n712), .B(n2427), .S(n2490), .Z(n1207) );
  INV_X1 U9664 ( .A(n2507), .ZN(n2427) );
  OAI21_X1 U9665 ( .B1(Din[17]), .B2(n2492), .A(n2493), .ZN(n2507) );
  MUX2_X1 U9666 ( .A(n713), .B(n2428), .S(n2490), .Z(n1206) );
  INV_X1 U9667 ( .A(n2508), .ZN(n2428) );
  OAI21_X1 U9668 ( .B1(Din[16]), .B2(n2492), .A(n2493), .ZN(n2508) );
  MUX2_X1 U9669 ( .A(n824), .B(n2429), .S(n2490), .Z(n1205) );
  INV_X1 U9670 ( .A(n2509), .ZN(n2429) );
  OAI21_X1 U9671 ( .B1(Din[15]), .B2(n2492), .A(n2493), .ZN(n2509) );
  OR2_X1 U9672 ( .A1(n2492), .A2(n2402), .ZN(n2493) );
  INV_X1 U9673 ( .A(n2510), .ZN(n2492) );
  AOI21_X1 U9674 ( .B1(n2408), .B2(Din[15]), .A(n2511), .ZN(n2510) );
  MUX2_X1 U9675 ( .A(n714), .B(n2430), .S(n2490), .Z(n1204) );
  INV_X1 U9676 ( .A(n2512), .ZN(n2430) );
  OAI21_X1 U9677 ( .B1(Din[14]), .B2(n2511), .A(n2513), .ZN(n2512) );
  MUX2_X1 U9678 ( .A(n715), .B(n2431), .S(n2490), .Z(n1203) );
  INV_X1 U9679 ( .A(n2514), .ZN(n2431) );
  OAI21_X1 U9680 ( .B1(Din[13]), .B2(n2511), .A(n2513), .ZN(n2514) );
  MUX2_X1 U9681 ( .A(n716), .B(n2432), .S(n2490), .Z(n1202) );
  INV_X1 U9682 ( .A(n2515), .ZN(n2432) );
  OAI21_X1 U9683 ( .B1(Din[12]), .B2(n2511), .A(n2513), .ZN(n2515) );
  MUX2_X1 U9684 ( .A(n717), .B(n2433), .S(n2490), .Z(n1201) );
  INV_X1 U9685 ( .A(n2516), .ZN(n2433) );
  OAI21_X1 U9686 ( .B1(Din[11]), .B2(n2511), .A(n2513), .ZN(n2516) );
  MUX2_X1 U9687 ( .A(n718), .B(n2434), .S(n2490), .Z(n1200) );
  INV_X1 U9688 ( .A(n2517), .ZN(n2434) );
  OAI21_X1 U9689 ( .B1(Din[10]), .B2(n2511), .A(n2513), .ZN(n2517) );
  MUX2_X1 U9690 ( .A(n719), .B(n2435), .S(n2490), .Z(n1199) );
  INV_X1 U9691 ( .A(n2518), .ZN(n2435) );
  OAI21_X1 U9692 ( .B1(Din[9]), .B2(n2511), .A(n2513), .ZN(n2518) );
  MUX2_X1 U9693 ( .A(n720), .B(n2436), .S(n2490), .Z(n1198) );
  INV_X1 U9694 ( .A(n2519), .ZN(n2436) );
  OAI21_X1 U9695 ( .B1(Din[8]), .B2(n2511), .A(n2513), .ZN(n2519) );
  INV_X1 U9696 ( .A(n2520), .ZN(n2511) );
  MUX2_X1 U9697 ( .A(n132), .B(n2437), .S(n2490), .Z(n1197) );
  AND2_X1 U9698 ( .A1(Din[7]), .A2(n2513), .ZN(n2437) );
  NAND2_X1 U9699 ( .A1(n2521), .A2(n2520), .ZN(n2513) );
  NAND2_X1 U9700 ( .A1(Din[7]), .A2(n2522), .ZN(n2520) );
  MUX2_X1 U9701 ( .A(n136), .B(n2438), .S(n2490), .Z(n1196) );
  AND2_X1 U9702 ( .A1(Din[6]), .A2(n2523), .ZN(n2438) );
  MUX2_X1 U9703 ( .A(n140), .B(n2439), .S(n2490), .Z(n1195) );
  AND2_X1 U9704 ( .A1(Din[5]), .A2(n2523), .ZN(n2439) );
  MUX2_X1 U9705 ( .A(n144), .B(n2440), .S(n2490), .Z(n1194) );
  AND2_X1 U9706 ( .A1(Din[4]), .A2(n2523), .ZN(n2440) );
  MUX2_X1 U9707 ( .A(n148), .B(n2441), .S(n2490), .Z(n1193) );
  AND2_X1 U9708 ( .A1(Din[3]), .A2(n2523), .ZN(n2441) );
  MUX2_X1 U9709 ( .A(n152), .B(n2442), .S(n2490), .Z(n1192) );
  AND2_X1 U9710 ( .A1(Din[2]), .A2(n2523), .ZN(n2442) );
  MUX2_X1 U9711 ( .A(n156), .B(n2443), .S(n2490), .Z(n1191) );
  AND2_X1 U9712 ( .A1(Din[1]), .A2(n2523), .ZN(n2443) );
  MUX2_X1 U9713 ( .A(n160), .B(n2444), .S(n2490), .Z(n1190) );
  AND2_X1 U9714 ( .A1(n2475), .A2(n2468), .ZN(n2487) );
  AND3_X1 U9715 ( .A1(EN), .A2(Addr[4]), .A3(WM), .ZN(n2475) );
  AND2_X1 U9716 ( .A1(Din[0]), .A2(n2523), .ZN(n2444) );
  OAI21_X1 U9717 ( .B1(Sel[2]), .B2(Sel[1]), .A(n2521), .ZN(n2523) );
  AND2_X1 U9718 ( .A1(RM), .A2(EN), .ZN(N598) );
  OAI21_X1 U9719 ( .B1(n2405), .B2(n2524), .A(n2407), .ZN(N581) );
  INV_X1 U9720 ( .A(n2525), .ZN(n2524) );
  AND4_X1 U9721 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2529), .ZN(n2405)
         );
  OAI21_X1 U9722 ( .B1(n2530), .B2(n2531), .A(n2410), .ZN(n2529) );
  OAI221_X1 U9723 ( .B1(n3509), .B2(n2532), .C1(n3459), .C2(n2533), .A(n2534), 
        .ZN(n2531) );
  AOI22_X1 U9724 ( .A1(n2383), .A2(n121), .B1(n2398), .B2(n357), .ZN(n2534) );
  OAI221_X1 U9725 ( .B1(n3217), .B2(n2535), .C1(n3135), .C2(n2536), .A(n2537), 
        .ZN(n2530) );
  AOI22_X1 U9726 ( .A1(n2393), .A2(n122), .B1(n2391), .B2(n358), .ZN(n2537) );
  OAI21_X1 U9727 ( .B1(n2538), .B2(n2539), .A(n2403), .ZN(n2528) );
  OAI221_X1 U9728 ( .B1(n3500), .B2(n2532), .C1(n3434), .C2(n2533), .A(n2540), 
        .ZN(n2539) );
  AOI22_X1 U9729 ( .A1(n2383), .A2(n123), .B1(n2398), .B2(n359), .ZN(n2540) );
  OAI221_X1 U9730 ( .B1(n3192), .B2(n2535), .C1(n3126), .C2(n2536), .A(n2541), 
        .ZN(n2538) );
  AOI22_X1 U9731 ( .A1(n2393), .A2(n124), .B1(n2391), .B2(n360), .ZN(n2541) );
  OAI21_X1 U9732 ( .B1(n2542), .B2(n2543), .A(n2409), .ZN(n2527) );
  OAI221_X1 U9733 ( .B1(n3475), .B2(n2532), .C1(n3409), .C2(n2533), .A(n2544), 
        .ZN(n2543) );
  AOI22_X1 U9734 ( .A1(n2383), .A2(n125), .B1(n2398), .B2(n361), .ZN(n2544) );
  OAI221_X1 U9735 ( .B1(n3167), .B2(n2535), .C1(n3101), .C2(n2536), .A(n2545), 
        .ZN(n2542) );
  AOI22_X1 U9736 ( .A1(n2393), .A2(n126), .B1(n2391), .B2(n362), .ZN(n2545) );
  OAI21_X1 U9737 ( .B1(n2546), .B2(n2547), .A(n2411), .ZN(n2526) );
  OAI221_X1 U9738 ( .B1(n3533), .B2(n2532), .C1(n3467), .C2(n2533), .A(n2548), 
        .ZN(n2547) );
  AOI22_X1 U9739 ( .A1(n2383), .A2(n127), .B1(n2398), .B2(n363), .ZN(n2548) );
  OAI221_X1 U9740 ( .B1(n3241), .B2(n2535), .C1(n3159), .C2(n2536), .A(n2549), 
        .ZN(n2546) );
  AOI22_X1 U9741 ( .A1(n2393), .A2(n128), .B1(n2391), .B2(n364), .ZN(n2549) );
  NAND2_X1 U9742 ( .A1(n2407), .A2(n2550), .ZN(N580) );
  OAI21_X1 U9743 ( .B1(n2551), .B2(n2552), .A(n2525), .ZN(n2550) );
  NAND4_X1 U9744 ( .A1(n2553), .A2(n2554), .A3(n2555), .A4(n2556), .ZN(n2552)
         );
  AOI221_X1 U9745 ( .B1(n2557), .B2(n253), .C1(n2558), .C2(n17), .A(n2559), 
        .ZN(n2556) );
  OAI22_X1 U9746 ( .A1(n2560), .A2(n429), .B1(n2561), .B2(n177), .ZN(n2559) );
  AOI221_X1 U9747 ( .B1(n2562), .B2(n254), .C1(n2563), .C2(n18), .A(n2564), 
        .ZN(n2555) );
  OAI22_X1 U9748 ( .A1(n2565), .A2(n430), .B1(n2566), .B2(n178), .ZN(n2564) );
  AOI221_X1 U9749 ( .B1(n2567), .B2(n255), .C1(n2568), .C2(n19), .A(n2569), 
        .ZN(n2554) );
  OAI22_X1 U9750 ( .A1(n3510), .A2(n2570), .B1(n3534), .B2(n2571), .ZN(n2569)
         );
  AOI221_X1 U9751 ( .B1(n2572), .B2(n256), .C1(n2573), .C2(n20), .A(n2574), 
        .ZN(n2553) );
  OAI22_X1 U9752 ( .A1(n3460), .A2(n2575), .B1(n3468), .B2(n2576), .ZN(n2574)
         );
  NAND4_X1 U9753 ( .A1(n2577), .A2(n2578), .A3(n2579), .A4(n2580), .ZN(n2551)
         );
  AOI221_X1 U9754 ( .B1(n2581), .B2(n257), .C1(n2582), .C2(n21), .A(n2583), 
        .ZN(n2580) );
  OAI22_X1 U9755 ( .A1(n2584), .A2(n431), .B1(n2585), .B2(n179), .ZN(n2583) );
  AOI221_X1 U9756 ( .B1(n2586), .B2(n258), .C1(n2587), .C2(n22), .A(n2588), 
        .ZN(n2579) );
  OAI22_X1 U9757 ( .A1(n2589), .A2(n432), .B1(n2590), .B2(n180), .ZN(n2588) );
  AOI221_X1 U9758 ( .B1(n2591), .B2(n259), .C1(n2592), .C2(n23), .A(n2593), 
        .ZN(n2578) );
  OAI22_X1 U9759 ( .A1(n3218), .A2(n2594), .B1(n3242), .B2(n2595), .ZN(n2593)
         );
  AOI221_X1 U9760 ( .B1(n2596), .B2(n260), .C1(n2597), .C2(n24), .A(n2598), 
        .ZN(n2577) );
  OAI22_X1 U9761 ( .A1(n3136), .A2(n2599), .B1(n3160), .B2(n2600), .ZN(n2598)
         );
  NAND2_X1 U9762 ( .A1(n2407), .A2(n2601), .ZN(N579) );
  OAI21_X1 U9763 ( .B1(n2602), .B2(n2603), .A(n2525), .ZN(n2601) );
  NAND4_X1 U9764 ( .A1(n2604), .A2(n2605), .A3(n2606), .A4(n2607), .ZN(n2603)
         );
  AOI221_X1 U9765 ( .B1(n2557), .B2(n261), .C1(n2558), .C2(n25), .A(n2608), 
        .ZN(n2607) );
  OAI22_X1 U9766 ( .A1(n2560), .A2(n433), .B1(n2561), .B2(n181), .ZN(n2608) );
  AOI221_X1 U9767 ( .B1(n2562), .B2(n262), .C1(n2563), .C2(n26), .A(n2609), 
        .ZN(n2606) );
  OAI22_X1 U9768 ( .A1(n2565), .A2(n434), .B1(n2566), .B2(n182), .ZN(n2609) );
  AOI221_X1 U9769 ( .B1(n2567), .B2(n263), .C1(n2568), .C2(n27), .A(n2610), 
        .ZN(n2605) );
  OAI22_X1 U9770 ( .A1(n3511), .A2(n2570), .B1(n3535), .B2(n2571), .ZN(n2610)
         );
  AOI221_X1 U9771 ( .B1(n2572), .B2(n264), .C1(n2573), .C2(n28), .A(n2611), 
        .ZN(n2604) );
  OAI22_X1 U9772 ( .A1(n3461), .A2(n2575), .B1(n3469), .B2(n2576), .ZN(n2611)
         );
  NAND4_X1 U9773 ( .A1(n2612), .A2(n2613), .A3(n2614), .A4(n2615), .ZN(n2602)
         );
  AOI221_X1 U9774 ( .B1(n2581), .B2(n265), .C1(n2582), .C2(n29), .A(n2616), 
        .ZN(n2615) );
  OAI22_X1 U9775 ( .A1(n2584), .A2(n435), .B1(n2585), .B2(n183), .ZN(n2616) );
  AOI221_X1 U9776 ( .B1(n2586), .B2(n266), .C1(n2587), .C2(n30), .A(n2617), 
        .ZN(n2614) );
  OAI22_X1 U9777 ( .A1(n2589), .A2(n436), .B1(n2590), .B2(n184), .ZN(n2617) );
  AOI221_X1 U9778 ( .B1(n2591), .B2(n267), .C1(n2592), .C2(n31), .A(n2618), 
        .ZN(n2613) );
  OAI22_X1 U9779 ( .A1(n3219), .A2(n2594), .B1(n3243), .B2(n2595), .ZN(n2618)
         );
  AOI221_X1 U9780 ( .B1(n2596), .B2(n268), .C1(n2597), .C2(n32), .A(n2619), 
        .ZN(n2612) );
  OAI22_X1 U9781 ( .A1(n3137), .A2(n2599), .B1(n3161), .B2(n2600), .ZN(n2619)
         );
  NAND2_X1 U9782 ( .A1(n2407), .A2(n2620), .ZN(N578) );
  OAI21_X1 U9783 ( .B1(n2621), .B2(n2622), .A(n2525), .ZN(n2620) );
  NAND4_X1 U9784 ( .A1(n2623), .A2(n2624), .A3(n2625), .A4(n2626), .ZN(n2622)
         );
  AOI221_X1 U9785 ( .B1(n2557), .B2(n269), .C1(n2558), .C2(n33), .A(n2627), 
        .ZN(n2626) );
  OAI22_X1 U9786 ( .A1(n2560), .A2(n437), .B1(n2561), .B2(n185), .ZN(n2627) );
  AOI221_X1 U9787 ( .B1(n2562), .B2(n270), .C1(n2563), .C2(n34), .A(n2628), 
        .ZN(n2625) );
  OAI22_X1 U9788 ( .A1(n2565), .A2(n438), .B1(n2566), .B2(n186), .ZN(n2628) );
  AOI221_X1 U9789 ( .B1(n2567), .B2(n271), .C1(n2568), .C2(n35), .A(n2629), 
        .ZN(n2624) );
  OAI22_X1 U9790 ( .A1(n3512), .A2(n2570), .B1(n3536), .B2(n2571), .ZN(n2629)
         );
  AOI221_X1 U9791 ( .B1(n2572), .B2(n272), .C1(n2573), .C2(n36), .A(n2630), 
        .ZN(n2623) );
  OAI22_X1 U9792 ( .A1(n3462), .A2(n2575), .B1(n3470), .B2(n2576), .ZN(n2630)
         );
  NAND4_X1 U9793 ( .A1(n2631), .A2(n2632), .A3(n2633), .A4(n2634), .ZN(n2621)
         );
  AOI221_X1 U9794 ( .B1(n2581), .B2(n273), .C1(n2582), .C2(n37), .A(n2635), 
        .ZN(n2634) );
  OAI22_X1 U9795 ( .A1(n2584), .A2(n439), .B1(n2585), .B2(n187), .ZN(n2635) );
  AOI221_X1 U9796 ( .B1(n2586), .B2(n274), .C1(n2587), .C2(n38), .A(n2636), 
        .ZN(n2633) );
  OAI22_X1 U9797 ( .A1(n2589), .A2(n440), .B1(n2590), .B2(n188), .ZN(n2636) );
  AOI221_X1 U9798 ( .B1(n2591), .B2(n275), .C1(n2592), .C2(n39), .A(n2637), 
        .ZN(n2632) );
  OAI22_X1 U9799 ( .A1(n3220), .A2(n2594), .B1(n3244), .B2(n2595), .ZN(n2637)
         );
  AOI221_X1 U9800 ( .B1(n2596), .B2(n276), .C1(n2597), .C2(n40), .A(n2638), 
        .ZN(n2631) );
  OAI22_X1 U9801 ( .A1(n3138), .A2(n2599), .B1(n3162), .B2(n2600), .ZN(n2638)
         );
  NAND2_X1 U9802 ( .A1(n2407), .A2(n2639), .ZN(N577) );
  OAI21_X1 U9803 ( .B1(n2640), .B2(n2641), .A(n2525), .ZN(n2639) );
  NAND4_X1 U9804 ( .A1(n2642), .A2(n2643), .A3(n2644), .A4(n2645), .ZN(n2641)
         );
  AOI221_X1 U9805 ( .B1(n2557), .B2(n277), .C1(n2558), .C2(n41), .A(n2646), 
        .ZN(n2645) );
  OAI22_X1 U9806 ( .A1(n2560), .A2(n441), .B1(n2561), .B2(n189), .ZN(n2646) );
  AOI221_X1 U9807 ( .B1(n2562), .B2(n278), .C1(n2563), .C2(n42), .A(n2647), 
        .ZN(n2644) );
  OAI22_X1 U9808 ( .A1(n2565), .A2(n442), .B1(n2566), .B2(n190), .ZN(n2647) );
  AOI221_X1 U9809 ( .B1(n2567), .B2(n279), .C1(n2568), .C2(n43), .A(n2648), 
        .ZN(n2643) );
  OAI22_X1 U9810 ( .A1(n3513), .A2(n2570), .B1(n3537), .B2(n2571), .ZN(n2648)
         );
  AOI221_X1 U9811 ( .B1(n2572), .B2(n280), .C1(n2573), .C2(n44), .A(n2649), 
        .ZN(n2642) );
  OAI22_X1 U9812 ( .A1(n3463), .A2(n2575), .B1(n3471), .B2(n2576), .ZN(n2649)
         );
  NAND4_X1 U9813 ( .A1(n2650), .A2(n2651), .A3(n2652), .A4(n2653), .ZN(n2640)
         );
  AOI221_X1 U9814 ( .B1(n2581), .B2(n281), .C1(n2582), .C2(n45), .A(n2654), 
        .ZN(n2653) );
  OAI22_X1 U9815 ( .A1(n2584), .A2(n443), .B1(n2585), .B2(n191), .ZN(n2654) );
  AOI221_X1 U9816 ( .B1(n2586), .B2(n282), .C1(n2587), .C2(n46), .A(n2655), 
        .ZN(n2652) );
  OAI22_X1 U9817 ( .A1(n2589), .A2(n444), .B1(n2590), .B2(n192), .ZN(n2655) );
  AOI221_X1 U9818 ( .B1(n2591), .B2(n283), .C1(n2592), .C2(n47), .A(n2656), 
        .ZN(n2651) );
  OAI22_X1 U9819 ( .A1(n3221), .A2(n2594), .B1(n3245), .B2(n2595), .ZN(n2656)
         );
  AOI221_X1 U9820 ( .B1(n2596), .B2(n284), .C1(n2597), .C2(n48), .A(n2657), 
        .ZN(n2650) );
  OAI22_X1 U9821 ( .A1(n3139), .A2(n2599), .B1(n3163), .B2(n2600), .ZN(n2657)
         );
  NAND2_X1 U9822 ( .A1(n2407), .A2(n2658), .ZN(N576) );
  OAI21_X1 U9823 ( .B1(n2659), .B2(n2660), .A(n2525), .ZN(n2658) );
  NAND4_X1 U9824 ( .A1(n2661), .A2(n2662), .A3(n2663), .A4(n2664), .ZN(n2660)
         );
  AOI221_X1 U9825 ( .B1(n2557), .B2(n285), .C1(n2558), .C2(n49), .A(n2665), 
        .ZN(n2664) );
  OAI22_X1 U9826 ( .A1(n2560), .A2(n445), .B1(n2561), .B2(n193), .ZN(n2665) );
  AOI221_X1 U9827 ( .B1(n2562), .B2(n286), .C1(n2563), .C2(n50), .A(n2666), 
        .ZN(n2663) );
  OAI22_X1 U9828 ( .A1(n2565), .A2(n446), .B1(n2566), .B2(n194), .ZN(n2666) );
  AOI221_X1 U9829 ( .B1(n2567), .B2(n287), .C1(n2568), .C2(n51), .A(n2667), 
        .ZN(n2662) );
  OAI22_X1 U9830 ( .A1(n3514), .A2(n2570), .B1(n3538), .B2(n2571), .ZN(n2667)
         );
  AOI221_X1 U9831 ( .B1(n2572), .B2(n288), .C1(n2573), .C2(n52), .A(n2668), 
        .ZN(n2661) );
  OAI22_X1 U9832 ( .A1(n3464), .A2(n2575), .B1(n3472), .B2(n2576), .ZN(n2668)
         );
  NAND4_X1 U9833 ( .A1(n2669), .A2(n2670), .A3(n2671), .A4(n2672), .ZN(n2659)
         );
  AOI221_X1 U9834 ( .B1(n2581), .B2(n289), .C1(n2582), .C2(n53), .A(n2673), 
        .ZN(n2672) );
  OAI22_X1 U9835 ( .A1(n2584), .A2(n447), .B1(n2585), .B2(n195), .ZN(n2673) );
  AOI221_X1 U9836 ( .B1(n2586), .B2(n290), .C1(n2587), .C2(n54), .A(n2674), 
        .ZN(n2671) );
  OAI22_X1 U9837 ( .A1(n2589), .A2(n448), .B1(n2590), .B2(n196), .ZN(n2674) );
  AOI221_X1 U9838 ( .B1(n2591), .B2(n291), .C1(n2592), .C2(n55), .A(n2675), 
        .ZN(n2670) );
  OAI22_X1 U9839 ( .A1(n3222), .A2(n2594), .B1(n3246), .B2(n2595), .ZN(n2675)
         );
  AOI221_X1 U9840 ( .B1(n2596), .B2(n292), .C1(n2597), .C2(n56), .A(n2676), 
        .ZN(n2669) );
  OAI22_X1 U9841 ( .A1(n3140), .A2(n2599), .B1(n3164), .B2(n2600), .ZN(n2676)
         );
  NAND2_X1 U9842 ( .A1(n2407), .A2(n2677), .ZN(N575) );
  OAI21_X1 U9843 ( .B1(n2678), .B2(n2679), .A(n2525), .ZN(n2677) );
  NAND4_X1 U9844 ( .A1(n2680), .A2(n2681), .A3(n2682), .A4(n2683), .ZN(n2679)
         );
  AOI221_X1 U9845 ( .B1(n2557), .B2(n293), .C1(n2558), .C2(n57), .A(n2684), 
        .ZN(n2683) );
  OAI22_X1 U9846 ( .A1(n2560), .A2(n449), .B1(n2561), .B2(n197), .ZN(n2684) );
  AOI221_X1 U9847 ( .B1(n2562), .B2(n294), .C1(n2563), .C2(n58), .A(n2685), 
        .ZN(n2682) );
  OAI22_X1 U9848 ( .A1(n2565), .A2(n450), .B1(n2566), .B2(n198), .ZN(n2685) );
  AOI221_X1 U9849 ( .B1(n2567), .B2(n295), .C1(n2568), .C2(n59), .A(n2686), 
        .ZN(n2681) );
  OAI22_X1 U9850 ( .A1(n3515), .A2(n2570), .B1(n3539), .B2(n2571), .ZN(n2686)
         );
  AOI221_X1 U9851 ( .B1(n2572), .B2(n296), .C1(n2573), .C2(n60), .A(n2687), 
        .ZN(n2680) );
  OAI22_X1 U9852 ( .A1(n3465), .A2(n2575), .B1(n3473), .B2(n2576), .ZN(n2687)
         );
  NAND4_X1 U9853 ( .A1(n2688), .A2(n2689), .A3(n2690), .A4(n2691), .ZN(n2678)
         );
  AOI221_X1 U9854 ( .B1(n2581), .B2(n297), .C1(n2582), .C2(n61), .A(n2692), 
        .ZN(n2691) );
  OAI22_X1 U9855 ( .A1(n2584), .A2(n451), .B1(n2585), .B2(n199), .ZN(n2692) );
  AOI221_X1 U9856 ( .B1(n2586), .B2(n298), .C1(n2587), .C2(n62), .A(n2693), 
        .ZN(n2690) );
  OAI22_X1 U9857 ( .A1(n2589), .A2(n452), .B1(n2590), .B2(n200), .ZN(n2693) );
  AOI221_X1 U9858 ( .B1(n2591), .B2(n299), .C1(n2592), .C2(n63), .A(n2694), 
        .ZN(n2689) );
  OAI22_X1 U9859 ( .A1(n3223), .A2(n2594), .B1(n3247), .B2(n2595), .ZN(n2694)
         );
  AOI221_X1 U9860 ( .B1(n2596), .B2(n300), .C1(n2597), .C2(n64), .A(n2695), 
        .ZN(n2688) );
  OAI22_X1 U9861 ( .A1(n3141), .A2(n2599), .B1(n3165), .B2(n2600), .ZN(n2695)
         );
  NAND2_X1 U9862 ( .A1(n2407), .A2(n2696), .ZN(N574) );
  OAI21_X1 U9863 ( .B1(n2697), .B2(n2698), .A(n2525), .ZN(n2696) );
  NAND2_X1 U9864 ( .A1(n2521), .A2(n2699), .ZN(n2525) );
  NOR2_X1 U9865 ( .A1(n2402), .A2(n2408), .ZN(n2521) );
  NOR3_X1 U9866 ( .A1(Sel[0]), .A2(Sel[2]), .A3(n2700), .ZN(n2408) );
  NOR2_X1 U9867 ( .A1(n2699), .A2(Sel[2]), .ZN(n2402) );
  NAND4_X1 U9868 ( .A1(n2701), .A2(n2702), .A3(n2703), .A4(n2704), .ZN(n2698)
         );
  AOI221_X1 U9869 ( .B1(n2557), .B2(n301), .C1(n2558), .C2(n65), .A(n2705), 
        .ZN(n2704) );
  OAI22_X1 U9870 ( .A1(n2560), .A2(n453), .B1(n2561), .B2(n201), .ZN(n2705) );
  AOI221_X1 U9871 ( .B1(n2562), .B2(n302), .C1(n2563), .C2(n66), .A(n2706), 
        .ZN(n2703) );
  OAI22_X1 U9872 ( .A1(n2565), .A2(n454), .B1(n2566), .B2(n202), .ZN(n2706) );
  AOI221_X1 U9873 ( .B1(n2567), .B2(n303), .C1(n2568), .C2(n67), .A(n2707), 
        .ZN(n2702) );
  OAI22_X1 U9874 ( .A1(n3516), .A2(n2570), .B1(n3540), .B2(n2571), .ZN(n2707)
         );
  INV_X1 U9875 ( .A(n2708), .ZN(n2568) );
  INV_X1 U9876 ( .A(n2709), .ZN(n2567) );
  AOI221_X1 U9877 ( .B1(n2572), .B2(n304), .C1(n2573), .C2(n68), .A(n2710), 
        .ZN(n2701) );
  OAI22_X1 U9878 ( .A1(n3466), .A2(n2575), .B1(n3474), .B2(n2576), .ZN(n2710)
         );
  INV_X1 U9879 ( .A(n2711), .ZN(n2573) );
  INV_X1 U9880 ( .A(n2712), .ZN(n2572) );
  NAND4_X1 U9881 ( .A1(n2713), .A2(n2714), .A3(n2715), .A4(n2716), .ZN(n2697)
         );
  AOI221_X1 U9882 ( .B1(n2581), .B2(n305), .C1(n2582), .C2(n69), .A(n2717), 
        .ZN(n2716) );
  OAI22_X1 U9883 ( .A1(n2584), .A2(n455), .B1(n2585), .B2(n203), .ZN(n2717) );
  AOI221_X1 U9884 ( .B1(n2586), .B2(n306), .C1(n2587), .C2(n70), .A(n2718), 
        .ZN(n2715) );
  OAI22_X1 U9885 ( .A1(n2589), .A2(n456), .B1(n2590), .B2(n204), .ZN(n2718) );
  AOI221_X1 U9886 ( .B1(n2591), .B2(n307), .C1(n2592), .C2(n71), .A(n2719), 
        .ZN(n2714) );
  OAI22_X1 U9887 ( .A1(n3224), .A2(n2594), .B1(n3248), .B2(n2595), .ZN(n2719)
         );
  INV_X1 U9888 ( .A(n2720), .ZN(n2592) );
  INV_X1 U9889 ( .A(n2721), .ZN(n2591) );
  AOI221_X1 U9890 ( .B1(n2596), .B2(n308), .C1(n2597), .C2(n72), .A(n2722), 
        .ZN(n2713) );
  OAI22_X1 U9891 ( .A1(n3142), .A2(n2599), .B1(n3166), .B2(n2600), .ZN(n2722)
         );
  INV_X1 U9892 ( .A(n2723), .ZN(n2597) );
  INV_X1 U9893 ( .A(n2724), .ZN(n2596) );
  NAND2_X1 U9894 ( .A1(n2522), .A2(n2725), .ZN(n2407) );
  NOR3_X1 U9895 ( .A1(Sel[1]), .A2(Sel[2]), .A3(n2726), .ZN(n2522) );
  NOR2_X1 U9896 ( .A1(n2727), .A2(n2728), .ZN(N573) );
  INV_X1 U9897 ( .A(n2725), .ZN(n2727) );
  NAND2_X1 U9898 ( .A1(n2729), .A2(n2730), .ZN(n2725) );
  NOR4_X1 U9899 ( .A1(n2731), .A2(n2732), .A3(n2733), .A4(n2734), .ZN(n2730)
         );
  OAI221_X1 U9900 ( .B1(n3127), .B2(n2724), .C1(n3102), .C2(n2723), .A(n2735), 
        .ZN(n2734) );
  AOI22_X1 U9901 ( .A1(n2736), .A2(n129), .B1(n2737), .B2(n365), .ZN(n2735) );
  OAI221_X1 U9902 ( .B1(n3193), .B2(n2721), .C1(n3168), .C2(n2720), .A(n2738), 
        .ZN(n2733) );
  AOI22_X1 U9903 ( .A1(n2739), .A2(n130), .B1(n2740), .B2(n366), .ZN(n2738) );
  OAI221_X1 U9904 ( .B1(n3093), .B2(n2590), .C1(n3085), .C2(n2589), .A(n2741), 
        .ZN(n2732) );
  AOI22_X1 U9905 ( .A1(n2977), .A2(n2586), .B1(n2978), .B2(n2587), .ZN(n2741)
         );
  OAI221_X1 U9906 ( .B1(n3077), .B2(n2585), .C1(n3062), .C2(n2584), .A(n2742), 
        .ZN(n2731) );
  AOI22_X1 U9907 ( .A1(n2975), .A2(n2581), .B1(n2976), .B2(n2582), .ZN(n2742)
         );
  NOR4_X1 U9908 ( .A1(n2743), .A2(n2744), .A3(n2745), .A4(n2746), .ZN(n2729)
         );
  OAI221_X1 U9909 ( .B1(n3435), .B2(n2712), .C1(n3410), .C2(n2711), .A(n2747), 
        .ZN(n2746) );
  AOI22_X1 U9910 ( .A1(n2748), .A2(n131), .B1(n2749), .B2(n367), .ZN(n2747) );
  OAI221_X1 U9911 ( .B1(n3501), .B2(n2709), .C1(n3476), .C2(n2708), .A(n2750), 
        .ZN(n2745) );
  AOI22_X1 U9912 ( .A1(n2751), .A2(n132), .B1(n2752), .B2(n368), .ZN(n2750) );
  OAI221_X1 U9913 ( .B1(n3353), .B2(n2566), .C1(n3329), .C2(n2565), .A(n2753), 
        .ZN(n2744) );
  AOI22_X1 U9914 ( .A1(n2981), .A2(n2562), .B1(n2982), .B2(n2563), .ZN(n2753)
         );
  OAI221_X1 U9915 ( .B1(n3273), .B2(n2561), .C1(n3265), .C2(n2560), .A(n2754), 
        .ZN(n2743) );
  AOI22_X1 U9916 ( .A1(n2979), .A2(n2557), .B1(n2980), .B2(n2558), .ZN(n2754)
         );
  AOI21_X1 U9917 ( .B1(n2755), .B2(n2756), .A(n2728), .ZN(N572) );
  NOR4_X1 U9918 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .ZN(n2756)
         );
  OAI221_X1 U9919 ( .B1(n3128), .B2(n2724), .C1(n3103), .C2(n2723), .A(n2761), 
        .ZN(n2760) );
  AOI22_X1 U9920 ( .A1(n2736), .A2(n133), .B1(n2737), .B2(n369), .ZN(n2761) );
  OAI221_X1 U9921 ( .B1(n3194), .B2(n2721), .C1(n3169), .C2(n2720), .A(n2762), 
        .ZN(n2759) );
  AOI22_X1 U9922 ( .A1(n2739), .A2(n134), .B1(n2740), .B2(n370), .ZN(n2762) );
  OAI221_X1 U9923 ( .B1(n3094), .B2(n2590), .C1(n3086), .C2(n2589), .A(n2763), 
        .ZN(n2758) );
  AOI22_X1 U9924 ( .A1(n2985), .A2(n2586), .B1(n2986), .B2(n2587), .ZN(n2763)
         );
  OAI221_X1 U9925 ( .B1(n3078), .B2(n2585), .C1(n3063), .C2(n2584), .A(n2764), 
        .ZN(n2757) );
  AOI22_X1 U9926 ( .A1(n2983), .A2(n2581), .B1(n2984), .B2(n2582), .ZN(n2764)
         );
  NOR4_X1 U9927 ( .A1(n2765), .A2(n2766), .A3(n2767), .A4(n2768), .ZN(n2755)
         );
  OAI221_X1 U9928 ( .B1(n3436), .B2(n2712), .C1(n3411), .C2(n2711), .A(n2769), 
        .ZN(n2768) );
  AOI22_X1 U9929 ( .A1(n2748), .A2(n135), .B1(n2749), .B2(n371), .ZN(n2769) );
  OAI221_X1 U9930 ( .B1(n3502), .B2(n2709), .C1(n3477), .C2(n2708), .A(n2770), 
        .ZN(n2767) );
  AOI22_X1 U9931 ( .A1(n2751), .A2(n136), .B1(n2752), .B2(n372), .ZN(n2770) );
  OAI221_X1 U9932 ( .B1(n3354), .B2(n2566), .C1(n3330), .C2(n2565), .A(n2771), 
        .ZN(n2766) );
  AOI22_X1 U9933 ( .A1(n2989), .A2(n2562), .B1(n2990), .B2(n2563), .ZN(n2771)
         );
  OAI221_X1 U9934 ( .B1(n3274), .B2(n2561), .C1(n3266), .C2(n2560), .A(n2772), 
        .ZN(n2765) );
  AOI22_X1 U9935 ( .A1(n2987), .A2(n2557), .B1(n2988), .B2(n2558), .ZN(n2772)
         );
  AOI21_X1 U9936 ( .B1(n2773), .B2(n2774), .A(n2728), .ZN(N571) );
  NOR4_X1 U9937 ( .A1(n2775), .A2(n2776), .A3(n2777), .A4(n2778), .ZN(n2774)
         );
  OAI221_X1 U9938 ( .B1(n3129), .B2(n2724), .C1(n3104), .C2(n2723), .A(n2779), 
        .ZN(n2778) );
  AOI22_X1 U9939 ( .A1(n2736), .A2(n137), .B1(n2737), .B2(n373), .ZN(n2779) );
  OAI221_X1 U9940 ( .B1(n3195), .B2(n2721), .C1(n3170), .C2(n2720), .A(n2780), 
        .ZN(n2777) );
  AOI22_X1 U9941 ( .A1(n2739), .A2(n138), .B1(n2740), .B2(n374), .ZN(n2780) );
  OAI221_X1 U9942 ( .B1(n3095), .B2(n2590), .C1(n3087), .C2(n2589), .A(n2781), 
        .ZN(n2776) );
  AOI22_X1 U9943 ( .A1(n2993), .A2(n2586), .B1(n2994), .B2(n2587), .ZN(n2781)
         );
  OAI221_X1 U9944 ( .B1(n3079), .B2(n2585), .C1(n3064), .C2(n2584), .A(n2782), 
        .ZN(n2775) );
  AOI22_X1 U9945 ( .A1(n2991), .A2(n2581), .B1(n2992), .B2(n2582), .ZN(n2782)
         );
  NOR4_X1 U9946 ( .A1(n2783), .A2(n2784), .A3(n2785), .A4(n2786), .ZN(n2773)
         );
  OAI221_X1 U9947 ( .B1(n3437), .B2(n2712), .C1(n3412), .C2(n2711), .A(n2787), 
        .ZN(n2786) );
  AOI22_X1 U9948 ( .A1(n2748), .A2(n139), .B1(n2749), .B2(n375), .ZN(n2787) );
  OAI221_X1 U9949 ( .B1(n3503), .B2(n2709), .C1(n3478), .C2(n2708), .A(n2788), 
        .ZN(n2785) );
  AOI22_X1 U9950 ( .A1(n2751), .A2(n140), .B1(n2752), .B2(n376), .ZN(n2788) );
  OAI221_X1 U9951 ( .B1(n3355), .B2(n2566), .C1(n3331), .C2(n2565), .A(n2789), 
        .ZN(n2784) );
  AOI22_X1 U9952 ( .A1(n2997), .A2(n2562), .B1(n2998), .B2(n2563), .ZN(n2789)
         );
  OAI221_X1 U9953 ( .B1(n3275), .B2(n2561), .C1(n3267), .C2(n2560), .A(n2790), 
        .ZN(n2783) );
  AOI22_X1 U9954 ( .A1(n2995), .A2(n2557), .B1(n2996), .B2(n2558), .ZN(n2790)
         );
  AOI21_X1 U9955 ( .B1(n2791), .B2(n2792), .A(n2728), .ZN(N570) );
  NOR4_X1 U9956 ( .A1(n2793), .A2(n2794), .A3(n2795), .A4(n2796), .ZN(n2792)
         );
  OAI221_X1 U9957 ( .B1(n3130), .B2(n2724), .C1(n3105), .C2(n2723), .A(n2797), 
        .ZN(n2796) );
  AOI22_X1 U9958 ( .A1(n2736), .A2(n141), .B1(n2737), .B2(n377), .ZN(n2797) );
  OAI221_X1 U9959 ( .B1(n3196), .B2(n2721), .C1(n3171), .C2(n2720), .A(n2798), 
        .ZN(n2795) );
  AOI22_X1 U9960 ( .A1(n2739), .A2(n142), .B1(n2740), .B2(n378), .ZN(n2798) );
  OAI221_X1 U9961 ( .B1(n3096), .B2(n2590), .C1(n3088), .C2(n2589), .A(n2799), 
        .ZN(n2794) );
  AOI22_X1 U9962 ( .A1(n3001), .A2(n2586), .B1(n3002), .B2(n2587), .ZN(n2799)
         );
  OAI221_X1 U9963 ( .B1(n3080), .B2(n2585), .C1(n3065), .C2(n2584), .A(n2800), 
        .ZN(n2793) );
  AOI22_X1 U9964 ( .A1(n2999), .A2(n2581), .B1(n3000), .B2(n2582), .ZN(n2800)
         );
  NOR4_X1 U9965 ( .A1(n2801), .A2(n2802), .A3(n2803), .A4(n2804), .ZN(n2791)
         );
  OAI221_X1 U9966 ( .B1(n3438), .B2(n2712), .C1(n3413), .C2(n2711), .A(n2805), 
        .ZN(n2804) );
  AOI22_X1 U9967 ( .A1(n2748), .A2(n143), .B1(n2749), .B2(n379), .ZN(n2805) );
  OAI221_X1 U9968 ( .B1(n3504), .B2(n2709), .C1(n3479), .C2(n2708), .A(n2806), 
        .ZN(n2803) );
  AOI22_X1 U9969 ( .A1(n2751), .A2(n144), .B1(n2752), .B2(n380), .ZN(n2806) );
  OAI221_X1 U9970 ( .B1(n3356), .B2(n2566), .C1(n3332), .C2(n2565), .A(n2807), 
        .ZN(n2802) );
  AOI22_X1 U9971 ( .A1(n3005), .A2(n2562), .B1(n3006), .B2(n2563), .ZN(n2807)
         );
  OAI221_X1 U9972 ( .B1(n3276), .B2(n2561), .C1(n3268), .C2(n2560), .A(n2808), 
        .ZN(n2801) );
  AOI22_X1 U9973 ( .A1(n3003), .A2(n2557), .B1(n3004), .B2(n2558), .ZN(n2808)
         );
  AOI21_X1 U9974 ( .B1(n2809), .B2(n2810), .A(n2728), .ZN(N569) );
  NOR4_X1 U9975 ( .A1(n2811), .A2(n2812), .A3(n2813), .A4(n2814), .ZN(n2810)
         );
  OAI221_X1 U9976 ( .B1(n3131), .B2(n2724), .C1(n3106), .C2(n2723), .A(n2815), 
        .ZN(n2814) );
  AOI22_X1 U9977 ( .A1(n2736), .A2(n145), .B1(n2737), .B2(n381), .ZN(n2815) );
  OAI221_X1 U9978 ( .B1(n3197), .B2(n2721), .C1(n3172), .C2(n2720), .A(n2816), 
        .ZN(n2813) );
  AOI22_X1 U9979 ( .A1(n2739), .A2(n146), .B1(n2740), .B2(n382), .ZN(n2816) );
  OAI221_X1 U9980 ( .B1(n3097), .B2(n2590), .C1(n3089), .C2(n2589), .A(n2817), 
        .ZN(n2812) );
  AOI22_X1 U9981 ( .A1(n3009), .A2(n2586), .B1(n3010), .B2(n2587), .ZN(n2817)
         );
  OAI221_X1 U9982 ( .B1(n3081), .B2(n2585), .C1(n3066), .C2(n2584), .A(n2818), 
        .ZN(n2811) );
  AOI22_X1 U9983 ( .A1(n3007), .A2(n2581), .B1(n3008), .B2(n2582), .ZN(n2818)
         );
  NOR4_X1 U9984 ( .A1(n2819), .A2(n2820), .A3(n2821), .A4(n2822), .ZN(n2809)
         );
  OAI221_X1 U9985 ( .B1(n3439), .B2(n2712), .C1(n3414), .C2(n2711), .A(n2823), 
        .ZN(n2822) );
  AOI22_X1 U9986 ( .A1(n2748), .A2(n147), .B1(n2749), .B2(n383), .ZN(n2823) );
  OAI221_X1 U9987 ( .B1(n3505), .B2(n2709), .C1(n3480), .C2(n2708), .A(n2824), 
        .ZN(n2821) );
  AOI22_X1 U9988 ( .A1(n2751), .A2(n148), .B1(n2752), .B2(n384), .ZN(n2824) );
  OAI221_X1 U9989 ( .B1(n3357), .B2(n2566), .C1(n3333), .C2(n2565), .A(n2825), 
        .ZN(n2820) );
  AOI22_X1 U9990 ( .A1(n3013), .A2(n2562), .B1(n3014), .B2(n2563), .ZN(n2825)
         );
  OAI221_X1 U9991 ( .B1(n3277), .B2(n2561), .C1(n3269), .C2(n2560), .A(n2826), 
        .ZN(n2819) );
  AOI22_X1 U9992 ( .A1(n3011), .A2(n2557), .B1(n3012), .B2(n2558), .ZN(n2826)
         );
  AOI21_X1 U9993 ( .B1(n2827), .B2(n2828), .A(n2728), .ZN(N568) );
  NOR4_X1 U9994 ( .A1(n2829), .A2(n2830), .A3(n2831), .A4(n2832), .ZN(n2828)
         );
  OAI221_X1 U9995 ( .B1(n3132), .B2(n2724), .C1(n3107), .C2(n2723), .A(n2833), 
        .ZN(n2832) );
  AOI22_X1 U9996 ( .A1(n2736), .A2(n149), .B1(n2737), .B2(n385), .ZN(n2833) );
  OAI221_X1 U9997 ( .B1(n3198), .B2(n2721), .C1(n3173), .C2(n2720), .A(n2834), 
        .ZN(n2831) );
  AOI22_X1 U9998 ( .A1(n2739), .A2(n150), .B1(n2740), .B2(n386), .ZN(n2834) );
  OAI221_X1 U9999 ( .B1(n3098), .B2(n2590), .C1(n3090), .C2(n2589), .A(n2835), 
        .ZN(n2830) );
  AOI22_X1 U10000 ( .A1(n3017), .A2(n2586), .B1(n3018), .B2(n2587), .ZN(n2835)
         );
  OAI221_X1 U10001 ( .B1(n3082), .B2(n2585), .C1(n3067), .C2(n2584), .A(n2836), 
        .ZN(n2829) );
  AOI22_X1 U10002 ( .A1(n3015), .A2(n2581), .B1(n3016), .B2(n2582), .ZN(n2836)
         );
  NOR4_X1 U10003 ( .A1(n2837), .A2(n2838), .A3(n2839), .A4(n2840), .ZN(n2827)
         );
  OAI221_X1 U10004 ( .B1(n3440), .B2(n2712), .C1(n3415), .C2(n2711), .A(n2841), 
        .ZN(n2840) );
  AOI22_X1 U10005 ( .A1(n2748), .A2(n151), .B1(n2749), .B2(n387), .ZN(n2841)
         );
  OAI221_X1 U10006 ( .B1(n3506), .B2(n2709), .C1(n3481), .C2(n2708), .A(n2842), 
        .ZN(n2839) );
  AOI22_X1 U10007 ( .A1(n2751), .A2(n152), .B1(n2752), .B2(n388), .ZN(n2842)
         );
  OAI221_X1 U10008 ( .B1(n3358), .B2(n2566), .C1(n3334), .C2(n2565), .A(n2843), 
        .ZN(n2838) );
  AOI22_X1 U10009 ( .A1(n3021), .A2(n2562), .B1(n3022), .B2(n2563), .ZN(n2843)
         );
  OAI221_X1 U10010 ( .B1(n3278), .B2(n2561), .C1(n3270), .C2(n2560), .A(n2844), 
        .ZN(n2837) );
  AOI22_X1 U10011 ( .A1(n3019), .A2(n2557), .B1(n3020), .B2(n2558), .ZN(n2844)
         );
  AOI21_X1 U10012 ( .B1(n2845), .B2(n2846), .A(n2728), .ZN(N567) );
  NOR4_X1 U10013 ( .A1(n2847), .A2(n2848), .A3(n2849), .A4(n2850), .ZN(n2846)
         );
  OAI221_X1 U10014 ( .B1(n3133), .B2(n2724), .C1(n3108), .C2(n2723), .A(n2851), 
        .ZN(n2850) );
  AOI22_X1 U10015 ( .A1(n2736), .A2(n153), .B1(n2737), .B2(n389), .ZN(n2851)
         );
  OAI221_X1 U10016 ( .B1(n3199), .B2(n2721), .C1(n3174), .C2(n2720), .A(n2852), 
        .ZN(n2849) );
  AOI22_X1 U10017 ( .A1(n2739), .A2(n154), .B1(n2740), .B2(n390), .ZN(n2852)
         );
  OAI221_X1 U10018 ( .B1(n3099), .B2(n2590), .C1(n3091), .C2(n2589), .A(n2853), 
        .ZN(n2848) );
  AOI22_X1 U10019 ( .A1(n3025), .A2(n2586), .B1(n3026), .B2(n2587), .ZN(n2853)
         );
  OAI221_X1 U10020 ( .B1(n3083), .B2(n2585), .C1(n3068), .C2(n2584), .A(n2854), 
        .ZN(n2847) );
  AOI22_X1 U10021 ( .A1(n3023), .A2(n2581), .B1(n3024), .B2(n2582), .ZN(n2854)
         );
  NOR4_X1 U10022 ( .A1(n2855), .A2(n2856), .A3(n2857), .A4(n2858), .ZN(n2845)
         );
  OAI221_X1 U10023 ( .B1(n3441), .B2(n2712), .C1(n3416), .C2(n2711), .A(n2859), 
        .ZN(n2858) );
  AOI22_X1 U10024 ( .A1(n2748), .A2(n155), .B1(n2749), .B2(n391), .ZN(n2859)
         );
  OAI221_X1 U10025 ( .B1(n3507), .B2(n2709), .C1(n3482), .C2(n2708), .A(n2860), 
        .ZN(n2857) );
  AOI22_X1 U10026 ( .A1(n2751), .A2(n156), .B1(n2752), .B2(n392), .ZN(n2860)
         );
  OAI221_X1 U10027 ( .B1(n3359), .B2(n2566), .C1(n3335), .C2(n2565), .A(n2861), 
        .ZN(n2856) );
  AOI22_X1 U10028 ( .A1(n3029), .A2(n2562), .B1(n3030), .B2(n2563), .ZN(n2861)
         );
  OAI221_X1 U10029 ( .B1(n3279), .B2(n2561), .C1(n3271), .C2(n2560), .A(n2862), 
        .ZN(n2855) );
  AOI22_X1 U10030 ( .A1(n3027), .A2(n2557), .B1(n3028), .B2(n2558), .ZN(n2862)
         );
  AOI21_X1 U10031 ( .B1(n2863), .B2(n2864), .A(n2728), .ZN(N566) );
  AND2_X1 U10032 ( .A1(Sel[2]), .A2(n2699), .ZN(n2728) );
  NAND2_X1 U10033 ( .A1(n2726), .A2(n2700), .ZN(n2699) );
  INV_X1 U10034 ( .A(Sel[1]), .ZN(n2700) );
  INV_X1 U10035 ( .A(Sel[0]), .ZN(n2726) );
  NOR4_X1 U10036 ( .A1(n2865), .A2(n2866), .A3(n2867), .A4(n2868), .ZN(n2864)
         );
  OAI221_X1 U10037 ( .B1(n3134), .B2(n2724), .C1(n3109), .C2(n2723), .A(n2869), 
        .ZN(n2868) );
  AOI22_X1 U10038 ( .A1(n2736), .A2(n157), .B1(n2737), .B2(n393), .ZN(n2869)
         );
  INV_X1 U10039 ( .A(n2599), .ZN(n2737) );
  NAND2_X1 U10040 ( .A1(n2410), .A2(n2385), .ZN(n2599) );
  INV_X1 U10041 ( .A(n2600), .ZN(n2736) );
  NAND2_X1 U10042 ( .A1(n2411), .A2(n2385), .ZN(n2600) );
  NAND2_X1 U10043 ( .A1(n2409), .A2(n2385), .ZN(n2723) );
  NAND2_X1 U10044 ( .A1(n2403), .A2(n2385), .ZN(n2724) );
  INV_X1 U10045 ( .A(n2536), .ZN(n2385) );
  NAND2_X1 U10046 ( .A1(n2462), .A2(n2469), .ZN(n2536) );
  OAI221_X1 U10047 ( .B1(n3200), .B2(n2721), .C1(n3175), .C2(n2720), .A(n2870), 
        .ZN(n2867) );
  AOI22_X1 U10048 ( .A1(n2739), .A2(n158), .B1(n2740), .B2(n394), .ZN(n2870)
         );
  INV_X1 U10049 ( .A(n2594), .ZN(n2740) );
  NAND2_X1 U10050 ( .A1(n2410), .A2(n2389), .ZN(n2594) );
  INV_X1 U10051 ( .A(n2595), .ZN(n2739) );
  NAND2_X1 U10052 ( .A1(n2411), .A2(n2389), .ZN(n2595) );
  NAND2_X1 U10053 ( .A1(n2409), .A2(n2389), .ZN(n2720) );
  NAND2_X1 U10054 ( .A1(n2403), .A2(n2389), .ZN(n2721) );
  INV_X1 U10055 ( .A(n2535), .ZN(n2389) );
  NAND2_X1 U10056 ( .A1(n2468), .A2(n2469), .ZN(n2535) );
  OAI221_X1 U10057 ( .B1(n3100), .B2(n2590), .C1(n3092), .C2(n2589), .A(n2871), 
        .ZN(n2866) );
  AOI22_X1 U10058 ( .A1(n3033), .A2(n2586), .B1(n3034), .B2(n2587), .ZN(n2871)
         );
  AND2_X1 U10059 ( .A1(n2410), .A2(n2391), .ZN(n2587) );
  AND2_X1 U10060 ( .A1(n2411), .A2(n2391), .ZN(n2586) );
  NAND2_X1 U10061 ( .A1(n2409), .A2(n2391), .ZN(n2589) );
  NAND2_X1 U10062 ( .A1(n2403), .A2(n2391), .ZN(n2590) );
  AND2_X1 U10063 ( .A1(n2456), .A2(n2469), .ZN(n2391) );
  OAI221_X1 U10064 ( .B1(n3084), .B2(n2585), .C1(n3069), .C2(n2584), .A(n2872), 
        .ZN(n2865) );
  AOI22_X1 U10065 ( .A1(n3031), .A2(n2581), .B1(n3032), .B2(n2582), .ZN(n2872)
         );
  AND2_X1 U10066 ( .A1(n2410), .A2(n2393), .ZN(n2582) );
  AND2_X1 U10067 ( .A1(n2411), .A2(n2393), .ZN(n2581) );
  NAND2_X1 U10068 ( .A1(n2409), .A2(n2393), .ZN(n2584) );
  NAND2_X1 U10069 ( .A1(n2403), .A2(n2393), .ZN(n2585) );
  AND2_X1 U10070 ( .A1(n2450), .A2(n2469), .ZN(n2393) );
  INV_X1 U10071 ( .A(Addr[4]), .ZN(n2469) );
  NOR4_X1 U10072 ( .A1(n2873), .A2(n2874), .A3(n2875), .A4(n2876), .ZN(n2863)
         );
  OAI221_X1 U10073 ( .B1(n3442), .B2(n2712), .C1(n3417), .C2(n2711), .A(n2877), 
        .ZN(n2876) );
  AOI22_X1 U10074 ( .A1(n2748), .A2(n159), .B1(n2749), .B2(n395), .ZN(n2877)
         );
  INV_X1 U10075 ( .A(n2575), .ZN(n2749) );
  NAND2_X1 U10076 ( .A1(n2410), .A2(n2401), .ZN(n2575) );
  INV_X1 U10077 ( .A(n2576), .ZN(n2748) );
  NAND2_X1 U10078 ( .A1(n2411), .A2(n2401), .ZN(n2576) );
  NAND2_X1 U10079 ( .A1(n2409), .A2(n2401), .ZN(n2711) );
  NAND2_X1 U10080 ( .A1(n2403), .A2(n2401), .ZN(n2712) );
  INV_X1 U10081 ( .A(n2533), .ZN(n2401) );
  NAND2_X1 U10082 ( .A1(Addr[4]), .A2(n2462), .ZN(n2533) );
  NOR2_X1 U10083 ( .A1(n2878), .A2(Addr[2]), .ZN(n2462) );
  OAI221_X1 U10084 ( .B1(n3508), .B2(n2709), .C1(n3483), .C2(n2708), .A(n2879), 
        .ZN(n2875) );
  AOI22_X1 U10085 ( .A1(n2751), .A2(n160), .B1(n2752), .B2(n396), .ZN(n2879)
         );
  INV_X1 U10086 ( .A(n2570), .ZN(n2752) );
  NAND2_X1 U10087 ( .A1(n2410), .A2(n2399), .ZN(n2570) );
  INV_X1 U10088 ( .A(n2571), .ZN(n2751) );
  NAND2_X1 U10089 ( .A1(n2411), .A2(n2399), .ZN(n2571) );
  NAND2_X1 U10090 ( .A1(n2409), .A2(n2399), .ZN(n2708) );
  NAND2_X1 U10091 ( .A1(n2403), .A2(n2399), .ZN(n2709) );
  INV_X1 U10092 ( .A(n2532), .ZN(n2399) );
  NAND2_X1 U10093 ( .A1(Addr[4]), .A2(n2468), .ZN(n2532) );
  NOR2_X1 U10094 ( .A1(n2878), .A2(n2880), .ZN(n2468) );
  INV_X1 U10095 ( .A(Addr[3]), .ZN(n2878) );
  OAI221_X1 U10096 ( .B1(n3360), .B2(n2566), .C1(n3336), .C2(n2565), .A(n2881), 
        .ZN(n2874) );
  AOI22_X1 U10097 ( .A1(n3037), .A2(n2562), .B1(n3038), .B2(n2563), .ZN(n2881)
         );
  AND2_X1 U10098 ( .A1(n2410), .A2(n2398), .ZN(n2563) );
  AND2_X1 U10099 ( .A1(n2411), .A2(n2398), .ZN(n2562) );
  NAND2_X1 U10100 ( .A1(n2409), .A2(n2398), .ZN(n2565) );
  NAND2_X1 U10101 ( .A1(n2403), .A2(n2398), .ZN(n2566) );
  AND2_X1 U10102 ( .A1(Addr[4]), .A2(n2456), .ZN(n2398) );
  NOR2_X1 U10103 ( .A1(n2880), .A2(Addr[3]), .ZN(n2456) );
  INV_X1 U10104 ( .A(Addr[2]), .ZN(n2880) );
  OAI221_X1 U10105 ( .B1(n3280), .B2(n2561), .C1(n3272), .C2(n2560), .A(n2882), 
        .ZN(n2873) );
  AOI22_X1 U10106 ( .A1(n3035), .A2(n2557), .B1(n3036), .B2(n2558), .ZN(n2882)
         );
  AND2_X1 U10107 ( .A1(n2410), .A2(n2383), .ZN(n2558) );
  AND2_X1 U10108 ( .A1(n2411), .A2(n2383), .ZN(n2557) );
  INV_X1 U10109 ( .A(Addr[1]), .ZN(n2883) );
  NAND2_X1 U10110 ( .A1(n2409), .A2(n2383), .ZN(n2560) );
  NAND2_X1 U10111 ( .A1(n2403), .A2(n2383), .ZN(n2561) );
  AND2_X1 U10112 ( .A1(Addr[4]), .A2(n2450), .ZN(n2383) );
  NOR2_X1 U10113 ( .A1(Addr[2]), .A2(Addr[3]), .ZN(n2450) );
  INV_X1 U10114 ( .A(Addr[0]), .ZN(n2884) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_0 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_63 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_62 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_61 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_60 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_59 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_58 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_57 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_56 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_55 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_54 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_53 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_52 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_51 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_50 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_49 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_48 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_47 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_46 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_45 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_44 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_43 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_42 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_41 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_40 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_39 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_38 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_37 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_36 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_35 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_34 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_33 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_32 MUX21GENI_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 MUX21GENI_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 MUX21GENI_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 MUX21GENI_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_28 MUX21GENI_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_27 MUX21GENI_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_26 MUX21GENI_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_25 MUX21GENI_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_24 MUX21GENI_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_23 MUX21GENI_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_22 MUX21GENI_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_21 MUX21GENI_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_20 MUX21GENI_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_19 MUX21GENI_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_18 MUX21GENI_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_17 MUX21GENI_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_16 MUX21GENI_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_15 MUX21GENI_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_14 MUX21GENI_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_13 MUX21GENI_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_12 MUX21GENI_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_11 MUX21GENI_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_10 MUX21GENI_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_9 MUX21GENI_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_8 MUX21GENI_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_7 MUX21GENI_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_6 MUX21GENI_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_5 MUX21GENI_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_4 MUX21GENI_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_3 MUX21GENI_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_2 MUX21GENI_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_1 MUX21GENI_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module MEMU ( CLK, RST, RM, WM, EN3, S3, S4, MEM_CFG, ALU_OUT, regBout, NPC2in, 
        RD3in, RD3out, WB_DATA );
  input [2:0] MEM_CFG;
  input [31:0] ALU_OUT;
  input [31:0] regBout;
  input [31:0] NPC2in;
  input [4:0] RD3in;
  output [4:0] RD3out;
  output [31:0] WB_DATA;
  input CLK, RST, RM, WM, EN3, S3, S4;

  wire   [31:0] DataMemOut;
  wire   [31:0] wb_prime;
  assign RD3out[4] = RD3in[4];
  assign RD3out[3] = RD3in[3];
  assign RD3out[2] = RD3in[2];
  assign RD3out[1] = RD3in[1];
  assign RD3out[0] = RD3in[0];

  DataMemory_RAM_DEPTH32_WORD_SIZE32 DRAM ( .Rst(RST), .Addr(ALU_OUT), .Din(
        regBout), .Dout(DataMemOut), .Sel(MEM_CFG), .RM(RM), .WM(WM), .EN(EN3), 
        .CLK(CLK) );
  MUX21_GENERIC_NBIT32_0 MUX21_ALMEM ( .A(DataMemOut), .B(ALU_OUT), .SEL(S3), 
        .Y(wb_prime) );
  MUX21_GENERIC_NBIT32_1 MUX21_NPCWB ( .A(NPC2in), .B(wb_prime), .SEL(S4), .Y(
        WB_DATA) );
endmodule

