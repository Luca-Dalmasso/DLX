
module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_2 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_3 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_4 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_5 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_7 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(net85111), .A2(TE), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_8 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_9 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_10 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_11 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_12 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_13 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_14 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_15 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_16 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_17 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_18 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_19 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_20 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_21 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_22 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_23 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_24 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_25 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_26 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_27 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_28 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_29 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_30 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_31 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net85111, n2, n3;
  assign net85111 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net85111), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module register_file_WORD_SIZE32_ADDR_SIZE5 ( CLK, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2, RESET );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, ENABLE, RD1, RD2, WR, RESET;
  wire   N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N444, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n4455), .CK(n4423), .QN(n2584) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n4456), .CK(n4423), .QN(n2585) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n4457), .CK(n4423), .QN(n2586) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n4458), .CK(n4423), .QN(n2587) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n4459), .CK(n4423), .QN(n2588) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n4460), .CK(n4423), .QN(n2589) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n4461), .CK(n4423), .QN(n2590) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n4462), .CK(n4423), .QN(n2591) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n4463), .CK(n4423), .QN(n2592) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n4464), .CK(n4423), .QN(n2593) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n4465), .CK(n4423), .QN(n2594) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n4466), .CK(n4423), .QN(n2595) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n4467), .CK(n4423), .QN(n2596) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n4468), .CK(n4423), .QN(n2597) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n4469), .CK(n4423), .QN(n2598) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n4470), .CK(n4423), .QN(n2599) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n4471), .CK(n4423), .QN(n2600) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n4472), .CK(n4423), .QN(n2601) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n4473), .CK(n4423), .QN(n2602) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n4474), .CK(n4423), .QN(n2603) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n4475), .CK(n4423), .QN(n2604) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n4476), .CK(n4423), .QN(n2605) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n4477), .CK(n4423), .QN(n2606) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n4478), .CK(n4423), .QN(n2607) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n4479), .CK(n4423), .QN(n2608) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n4480), .CK(n4423), .QN(n2609) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n4481), .CK(n4423), .QN(n2610) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n4482), .CK(n4423), .QN(n2611) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n4483), .CK(n4423), .QN(n2612) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n4484), .CK(n4423), .QN(n2613) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n4485), .CK(n4423), .QN(n2614) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n4486), .CK(n4423), .QN(n2615) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n4455), .CK(n4435), .QN(n2616) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n4456), .CK(n4435), .QN(n2617) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n4457), .CK(n4435), .QN(n2618) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n4458), .CK(n4435), .QN(n2619) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n4459), .CK(n4435), .QN(n2620) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n4460), .CK(n4435), .QN(n2621) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n4461), .CK(n4435), .QN(n2622) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n4462), .CK(n4435), .QN(n2623) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n4463), .CK(n4435), .QN(n2624) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n4464), .CK(n4435), .QN(n2625) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n4465), .CK(n4435), .QN(n2626) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n4466), .CK(n4435), .QN(n2627) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n4467), .CK(n4435), .QN(n2628) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n4468), .CK(n4435), .QN(n2629) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n4469), .CK(n4435), .QN(n2630) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n4470), .CK(n4435), .QN(n2631) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n4471), .CK(n4435), .QN(n2632) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n4472), .CK(n4435), .QN(n2633) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n4473), .CK(n4435), .QN(n2634) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n4474), .CK(n4435), .QN(n2635) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n4475), .CK(n4435), .QN(n2636) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n4476), .CK(n4435), .QN(n2637) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n4477), .CK(n4435), .QN(n2638) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n4478), .CK(n4435), .QN(n2639) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n4479), .CK(n4435), .QN(n2640) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n4480), .CK(n4435), .QN(n2641) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n4481), .CK(n4435), .QN(n2642) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n4482), .CK(n4435), .QN(n2643) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n4483), .CK(n4435), .QN(n2644) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n4484), .CK(n4435), .QN(n2645) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n4485), .CK(n4435), .QN(n2646) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n4486), .CK(n4435), .QN(n2647) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n4455), .CK(n4446), .QN(n2648) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n4456), .CK(n4446), .QN(n2649) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n4457), .CK(n4446), .QN(n2650) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n4458), .CK(n4446), .QN(n2651) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n4459), .CK(n4446), .QN(n2652) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n4460), .CK(n4446), .QN(n2653) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n4461), .CK(n4446), .QN(n2654) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n4462), .CK(n4446), .QN(n2655) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n4463), .CK(n4446), .QN(n2656) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n4464), .CK(n4446), .QN(n2657) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n4465), .CK(n4446), .QN(n2658) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n4466), .CK(n4446), .QN(n2659) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n4467), .CK(n4446), .QN(n2660) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n4468), .CK(n4446), .QN(n2661) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n4469), .CK(n4446), .QN(n2662) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n4470), .CK(n4446), .QN(n2663) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n4471), .CK(n4446), .QN(n2664) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n4472), .CK(n4446), .QN(n2665) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n4473), .CK(n4446), .QN(n2666) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n4474), .CK(n4446), .QN(n2667) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n4475), .CK(n4446), .QN(n2668) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n4476), .CK(n4446), .QN(n2669) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n4477), .CK(n4446), .QN(n2670) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n4478), .CK(n4446), .QN(n2671) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n4479), .CK(n4446), .QN(n2672) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n4480), .CK(n4446), .QN(n2673) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n4481), .CK(n4446), .QN(n2674) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n4482), .CK(n4446), .QN(n2675) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n4483), .CK(n4446), .QN(n2676) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n4484), .CK(n4446), .QN(n2677) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n4485), .CK(n4446), .QN(n2678) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n4486), .CK(n4446), .QN(n2679) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n4455), .CK(n4449), .QN(n2680) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n4456), .CK(n4449), .QN(n2681) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n4457), .CK(n4449), .QN(n2682) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n4458), .CK(n4449), .QN(n2683) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n4459), .CK(n4449), .QN(n2684) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n4460), .CK(n4449), .QN(n2685) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n4461), .CK(n4449), .QN(n2686) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n4462), .CK(n4449), .QN(n2687) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n4463), .CK(n4449), .QN(n2688) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n4464), .CK(n4449), .QN(n2689) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n4465), .CK(n4449), .QN(n2690) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n4466), .CK(n4449), .QN(n2691) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n4467), .CK(n4449), .QN(n2692) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n4468), .CK(n4449), .QN(n2693) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n4469), .CK(n4449), .QN(n2694) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n4470), .CK(n4449), .QN(n2695) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n4471), .CK(n4449), .QN(n2696) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n4472), .CK(n4449), .QN(n2697) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n4473), .CK(n4449), .QN(n2698) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n4474), .CK(n4449), .QN(n2699) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n4475), .CK(n4449), .QN(n2700) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n4476), .CK(n4449), .QN(n2701) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n4477), .CK(n4449), .QN(n2702) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n4478), .CK(n4449), .QN(n2703) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n4479), .CK(n4449), .QN(n2704) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n4480), .CK(n4449), .QN(n2705) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n4481), .CK(n4449), .QN(n2706) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n4482), .CK(n4449), .QN(n2707) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n4483), .CK(n4449), .QN(n2708) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n4484), .CK(n4449), .QN(n2709) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n4485), .CK(n4449), .QN(n2710) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n4486), .CK(n4449), .QN(n2711) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n4455), .CK(n4450), .QN(n2712) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n4456), .CK(n4450), .QN(n2713) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n4457), .CK(n4450), .QN(n2714) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n4458), .CK(n4450), .QN(n2715) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n4459), .CK(n4450), .QN(n2716) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n4460), .CK(n4450), .QN(n2717) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n4461), .CK(n4450), .QN(n2718) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n4462), .CK(n4450), .QN(n2719) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n4463), .CK(n4450), .QN(n2720) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n4464), .CK(n4450), .QN(n2721) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n4465), .CK(n4450), .QN(n2722) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n4466), .CK(n4450), .QN(n2723) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n4467), .CK(n4450), .QN(n2724) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n4468), .CK(n4450), .QN(n2725) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n4469), .CK(n4450), .QN(n2726) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n4470), .CK(n4450), .QN(n2727) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n4471), .CK(n4450), .QN(n2728) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n4472), .CK(n4450), .QN(n2729) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n4473), .CK(n4450), .QN(n2730) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n4474), .CK(n4450), .QN(n2731) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n4475), .CK(n4450), .QN(n2732) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n4476), .CK(n4450), .QN(n2733) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n4477), .CK(n4450), .QN(n2734) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n4478), .CK(n4450), .QN(n2735) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n4479), .CK(n4450), .QN(n2736) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n4480), .CK(n4450), .QN(n2737) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n4481), .CK(n4450), .QN(n2738) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n4482), .CK(n4450), .QN(n2739) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n4483), .CK(n4450), .QN(n2740) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n4484), .CK(n4450), .QN(n2741) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n4485), .CK(n4450), .QN(n2742) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n4486), .CK(n4450), .QN(n2743) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n4455), .CK(n4451), .QN(n2744) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n4456), .CK(n4451), .QN(n2745) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n4457), .CK(n4451), .QN(n2746) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n4458), .CK(n4451), .QN(n2747) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n4459), .CK(n4451), .QN(n2748) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n4460), .CK(n4451), .QN(n2749) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n4461), .CK(n4451), .QN(n2750) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n4462), .CK(n4451), .QN(n2751) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n4463), .CK(n4451), .QN(n2752) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n4464), .CK(n4451), .QN(n2753) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n4465), .CK(n4451), .QN(n2754) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n4466), .CK(n4451), .QN(n2755) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n4467), .CK(n4451), .QN(n2756) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n4468), .CK(n4451), .QN(n2757) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n4469), .CK(n4451), .QN(n2758) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n4470), .CK(n4451), .QN(n2759) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n4471), .CK(n4451), .QN(n2760) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n4472), .CK(n4451), .QN(n2761) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n4473), .CK(n4451), .QN(n2762) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n4474), .CK(n4451), .QN(n2763) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n4475), .CK(n4451), .QN(n2764) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n4476), .CK(n4451), .QN(n2765) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n4477), .CK(n4451), .QN(n2766) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n4478), .CK(n4451), .QN(n2767) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n4479), .CK(n4451), .QN(n2768) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n4480), .CK(n4451), .QN(n2769) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n4481), .CK(n4451), .QN(n2770) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n4482), .CK(n4451), .QN(n2771) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n4483), .CK(n4451), .QN(n2772) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n4484), .CK(n4451), .QN(n2773) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n4485), .CK(n4451), .QN(n2774) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n4486), .CK(n4451), .QN(n2775) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n4455), .CK(n4452), .QN(n2776) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n4456), .CK(n4452), .QN(n2777) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n4457), .CK(n4452), .QN(n2778) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n4458), .CK(n4452), .QN(n2779) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n4459), .CK(n4452), .QN(n2780) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n4460), .CK(n4452), .QN(n2781) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n4461), .CK(n4452), .QN(n2782) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n4462), .CK(n4452), .QN(n2783) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n4463), .CK(n4452), .QN(n2784) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n4464), .CK(n4452), .QN(n2785) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n4465), .CK(n4452), .QN(n2786) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n4466), .CK(n4452), .QN(n2787) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n4467), .CK(n4452), .QN(n2788) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n4468), .CK(n4452), .QN(n2789) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n4469), .CK(n4452), .QN(n2790) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n4470), .CK(n4452), .QN(n2791) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n4471), .CK(n4452), .QN(n2792) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n4472), .CK(n4452), .QN(n2793) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n4473), .CK(n4452), .QN(n2794) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n4474), .CK(n4452), .QN(n2795) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n4475), .CK(n4452), .QN(n2796) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n4476), .CK(n4452), .QN(n2797) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n4477), .CK(n4452), .QN(n2798) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n4478), .CK(n4452), .QN(n2799) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n4479), .CK(n4452), .QN(n2800) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n4480), .CK(n4452), .QN(n2801) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n4481), .CK(n4452), .QN(n2802) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n4482), .CK(n4452), .QN(n2803) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n4483), .CK(n4452), .QN(n2804) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n4484), .CK(n4452), .QN(n2805) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n4485), .CK(n4452), .QN(n2806) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n4486), .CK(n4452), .QN(n2807) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n4455), .CK(n4453), .QN(n2808) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n4456), .CK(n4453), .QN(n2809) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n4457), .CK(n4453), .QN(n2810) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n4458), .CK(n4453), .QN(n2811) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n4459), .CK(n4453), .QN(n2812) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n4460), .CK(n4453), .QN(n2813) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n4461), .CK(n4453), .QN(n2814) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n4462), .CK(n4453), .QN(n2815) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n4463), .CK(n4453), .QN(n2816) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n4464), .CK(n4453), .QN(n2817) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n4465), .CK(n4453), .QN(n2818) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n4466), .CK(n4453), .QN(n2819) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n4467), .CK(n4453), .QN(n2820) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n4468), .CK(n4453), .QN(n2821) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n4469), .CK(n4453), .QN(n2822) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n4470), .CK(n4453), .QN(n2823) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n4471), .CK(n4453), .QN(n2824) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n4472), .CK(n4453), .QN(n2825) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n4473), .CK(n4453), .QN(n2826) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n4474), .CK(n4453), .QN(n2827) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n4475), .CK(n4453), .QN(n2828) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n4476), .CK(n4453), .QN(n2829) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n4477), .CK(n4453), .QN(n2830) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n4478), .CK(n4453), .QN(n2831) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n4479), .CK(n4453), .QN(n2832) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n4480), .CK(n4453), .QN(n2833) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n4481), .CK(n4453), .QN(n2834) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n4482), .CK(n4453), .QN(n2835) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n4483), .CK(n4453), .QN(n2836) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n4484), .CK(n4453), .QN(n2837) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n4485), .CK(n4453), .QN(n2838) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n4486), .CK(n4453), .QN(n2839) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n4455), .CK(n4454), .QN(n2840) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n4456), .CK(n4454), .QN(n2841) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n4457), .CK(n4454), .QN(n2842) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n4458), .CK(n4454), .QN(n2843) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n4459), .CK(n4454), .QN(n2844) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n4460), .CK(n4454), .QN(n2845) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n4461), .CK(n4454), .QN(n2846) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n4462), .CK(n4454), .QN(n2847) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n4463), .CK(n4454), .QN(n2848) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n4464), .CK(n4454), .QN(n2849) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n4465), .CK(n4454), .QN(n2850) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n4466), .CK(n4454), .QN(n2851) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n4467), .CK(n4454), .QN(n2852) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n4468), .CK(n4454), .QN(n2853) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n4469), .CK(n4454), .QN(n2854) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n4470), .CK(n4454), .QN(n2855) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n4471), .CK(n4454), .QN(n2856) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n4472), .CK(n4454), .QN(n2857) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n4473), .CK(n4454), .QN(n2858) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n4474), .CK(n4454), .QN(n2859) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n4475), .CK(n4454), .QN(n2860) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n4476), .CK(n4454), .QN(n2861) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n4477), .CK(n4454), .QN(n2862) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n4478), .CK(n4454), .QN(n2863) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n4479), .CK(n4454), .QN(n2864) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n4480), .CK(n4454), .QN(n2865) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n4481), .CK(n4454), .QN(n2866) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n4482), .CK(n4454), .QN(n2867) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n4483), .CK(n4454), .QN(n2868) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n4484), .CK(n4454), .QN(n2869) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n4485), .CK(n4454), .QN(n2870) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n4486), .CK(n4454), .QN(n2871) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n4455), .CK(n4487), .QN(n2872) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n4456), .CK(n4487), .QN(n2873) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n4457), .CK(n4487), .QN(n2874) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n4458), .CK(n4487), .QN(n2875) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n4459), .CK(n4487), .QN(n2876) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n4460), .CK(n4487), .QN(n2877) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n4461), .CK(n4487), .QN(n2878) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n4462), .CK(n4487), .QN(n2879) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n4463), .CK(n4487), .QN(n2880) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n4464), .CK(n4487), .QN(n2881) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n4465), .CK(n4487), .QN(n2882) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n4466), .CK(n4487), .QN(n2883) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n4467), .CK(n4487), .QN(n2884) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n4468), .CK(n4487), .QN(n2885) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n4469), .CK(n4487), .QN(n2886) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n4470), .CK(n4487), .QN(n2887) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n4471), .CK(n4487), .QN(n2888) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n4472), .CK(n4487), .QN(n2889) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n4473), .CK(n4487), .QN(n2890) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n4474), .CK(n4487), .QN(n2891) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n4475), .CK(n4487), .QN(n2892) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n4476), .CK(n4487), .QN(n2893) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n4477), .CK(n4487), .QN(n2894) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n4478), .CK(n4487), .QN(n2895) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n4479), .CK(n4487), .QN(n2896) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n4480), .CK(n4487), .QN(n2897) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n4481), .CK(n4487), .QN(n2898) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n4482), .CK(n4487), .QN(n2899) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n4483), .CK(n4487), .QN(n2900) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n4484), .CK(n4487), .QN(n2901) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n4485), .CK(n4487), .QN(n2902) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n4486), .CK(n4487), .QN(n2903) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n4455), .CK(n4425), .QN(n2904) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n4456), .CK(n4425), .QN(n2905) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n4457), .CK(n4425), .QN(n2906) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n4458), .CK(n4425), .QN(n2907) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n4459), .CK(n4425), .QN(n2908) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n4460), .CK(n4425), .QN(n2909) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n4461), .CK(n4425), .QN(n2910) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n4462), .CK(n4425), .QN(n2911) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n4463), .CK(n4425), .QN(n2912) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n4464), .CK(n4425), .QN(n2913) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n4465), .CK(n4425), .QN(n2914) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n4466), .CK(n4425), .QN(n2915) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n4467), .CK(n4425), .QN(n2916) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n4468), .CK(n4425), .QN(n2917) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n4469), .CK(n4425), .QN(n2918) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n4470), .CK(n4425), .QN(n2919) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n4471), .CK(n4425), .QN(n2920) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n4472), .CK(n4425), .QN(n2921) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n4473), .CK(n4425), .QN(n2922) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n4474), .CK(n4425), .QN(n2923) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n4475), .CK(n4425), .QN(n2924) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n4476), .CK(n4425), .QN(n2925) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n4477), .CK(n4425), .QN(n2926) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n4478), .CK(n4425), .QN(n2927) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n4479), .CK(n4425), .QN(n2928) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n4480), .CK(n4425), .QN(n2929) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n4481), .CK(n4425), .QN(n2930) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n4482), .CK(n4425), .QN(n2931) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n4483), .CK(n4425), .QN(n2932) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n4484), .CK(n4425), .QN(n2933) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n4485), .CK(n4425), .QN(n2934) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n4486), .CK(n4425), .QN(n2935) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n4455), .CK(n4426), .QN(n2936) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n4456), .CK(n4426), .QN(n2937) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n4457), .CK(n4426), .QN(n2938) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n4458), .CK(n4426), .QN(n2939) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n4459), .CK(n4426), .QN(n2940) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n4460), .CK(n4426), .QN(n2941) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n4461), .CK(n4426), .QN(n2942) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n4462), .CK(n4426), .QN(n2943) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n4463), .CK(n4426), .QN(n2944) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n4464), .CK(n4426), .QN(n2945) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n4465), .CK(n4426), .QN(n2946) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n4466), .CK(n4426), .QN(n2947) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n4467), .CK(n4426), .QN(n2948) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n4468), .CK(n4426), .QN(n2949) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n4469), .CK(n4426), .QN(n2950) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n4470), .CK(n4426), .QN(n2951) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n4471), .CK(n4426), .QN(n2952) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n4472), .CK(n4426), .QN(n2953) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n4473), .CK(n4426), .QN(n2954) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n4474), .CK(n4426), .QN(n2955) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n4475), .CK(n4426), .QN(n2956) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n4476), .CK(n4426), .QN(n2957) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n4477), .CK(n4426), .QN(n2958) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n4478), .CK(n4426), .QN(n2959) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n4479), .CK(n4426), .QN(n2960) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n4480), .CK(n4426), .QN(n2961) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n4481), .CK(n4426), .QN(n2962) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n4482), .CK(n4426), .QN(n2963) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n4483), .CK(n4426), .QN(n2964) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n4484), .CK(n4426), .QN(n2965) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n4485), .CK(n4426), .QN(n2966) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n4486), .CK(n4426), .QN(n2967) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n4455), .CK(n4427), .QN(n2968) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n4456), .CK(n4427), .QN(n2969) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n4457), .CK(n4427), .QN(n2970) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n4458), .CK(n4427), .QN(n2971) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n4459), .CK(n4427), .QN(n2972) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n4460), .CK(n4427), .QN(n2973) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n4461), .CK(n4427), .QN(n2974) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n4462), .CK(n4427), .QN(n2975) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n4463), .CK(n4427), .QN(n2976) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n4464), .CK(n4427), .QN(n2977) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n4465), .CK(n4427), .QN(n2978) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n4466), .CK(n4427), .QN(n2979) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n4467), .CK(n4427), .QN(n2980) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n4468), .CK(n4427), .QN(n2981) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n4469), .CK(n4427), .QN(n2982) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n4470), .CK(n4427), .QN(n2983) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n4471), .CK(n4427), .QN(n2984) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n4472), .CK(n4427), .QN(n2985) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n4473), .CK(n4427), .QN(n2986) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n4474), .CK(n4427), .QN(n2987) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n4475), .CK(n4427), .QN(n2988) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n4476), .CK(n4427), .QN(n2989) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n4477), .CK(n4427), .QN(n2990) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n4478), .CK(n4427), .QN(n2991) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n4479), .CK(n4427), .QN(n2992) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n4480), .CK(n4427), .QN(n2993) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n4481), .CK(n4427), .QN(n2994) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n4482), .CK(n4427), .QN(n2995) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n4483), .CK(n4427), .QN(n2996) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n4484), .CK(n4427), .QN(n2997) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n4485), .CK(n4427), .QN(n2998) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n4486), .CK(n4427), .QN(n2999) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n4455), .CK(n4428), .QN(n3000) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n4456), .CK(n4428), .QN(n3001) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n4457), .CK(n4428), .QN(n3002) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n4458), .CK(n4428), .QN(n3003) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n4459), .CK(n4428), .QN(n3004) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n4460), .CK(n4428), .QN(n3005) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n4461), .CK(n4428), .QN(n3006) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n4462), .CK(n4428), .QN(n3007) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n4463), .CK(n4428), .QN(n3008) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n4464), .CK(n4428), .QN(n3009) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n4465), .CK(n4428), .QN(n3010) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n4466), .CK(n4428), .QN(n3011) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n4467), .CK(n4428), .QN(n3012) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n4468), .CK(n4428), .QN(n3013) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n4469), .CK(n4428), .QN(n3014) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n4470), .CK(n4428), .QN(n3015) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n4471), .CK(n4428), .QN(n3016) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n4472), .CK(n4428), .QN(n3017) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n4473), .CK(n4428), .QN(n3018) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n4474), .CK(n4428), .QN(n3019) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n4475), .CK(n4428), .QN(n3020) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n4476), .CK(n4428), .QN(n3021) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n4477), .CK(n4428), .QN(n3022) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n4478), .CK(n4428), .QN(n3023) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n4479), .CK(n4428), .QN(n3024) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n4480), .CK(n4428), .QN(n3025) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n4481), .CK(n4428), .QN(n3026) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n4482), .CK(n4428), .QN(n3027) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n4483), .CK(n4428), .QN(n3028) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n4484), .CK(n4428), .QN(n3029) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n4485), .CK(n4428), .QN(n3030) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n4486), .CK(n4428), .QN(n3031) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n4455), .CK(n4429), .QN(n3032) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n4456), .CK(n4429), .QN(n3033) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n4457), .CK(n4429), .QN(n3034) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n4458), .CK(n4429), .QN(n3035) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n4459), .CK(n4429), .QN(n3036) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n4460), .CK(n4429), .QN(n3037) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n4461), .CK(n4429), .QN(n3038) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n4462), .CK(n4429), .QN(n3039) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n4463), .CK(n4429), .QN(n3040) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n4464), .CK(n4429), .QN(n3041) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n4465), .CK(n4429), .QN(n3042) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n4466), .CK(n4429), .QN(n3043) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n4467), .CK(n4429), .QN(n3044) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n4468), .CK(n4429), .QN(n3045) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n4469), .CK(n4429), .QN(n3046) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n4470), .CK(n4429), .QN(n3047) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n4471), .CK(n4429), .QN(n3048) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n4472), .CK(n4429), .QN(n3049) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n4473), .CK(n4429), .QN(n3050) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n4474), .CK(n4429), .QN(n3051) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n4475), .CK(n4429), .QN(n3052) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n4476), .CK(n4429), .QN(n3053) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n4477), .CK(n4429), .QN(n3054) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n4478), .CK(n4429), .QN(n3055) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n4479), .CK(n4429), .QN(n3056) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n4480), .CK(n4429), .QN(n3057) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n4481), .CK(n4429), .QN(n3058) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n4482), .CK(n4429), .QN(n3059) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n4483), .CK(n4429), .QN(n3060) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n4484), .CK(n4429), .QN(n3061) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n4485), .CK(n4429), .QN(n3062) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n4486), .CK(n4429), .QN(n3063) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n4455), .CK(n4430), .QN(n3064) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n4456), .CK(n4430), .QN(n3065) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n4457), .CK(n4430), .QN(n3066) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n4458), .CK(n4430), .QN(n3067) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n4459), .CK(n4430), .QN(n3068) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n4460), .CK(n4430), .QN(n3069) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n4461), .CK(n4430), .QN(n3070) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n4462), .CK(n4430), .QN(n3071) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n4463), .CK(n4430), .QN(n3072) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n4464), .CK(n4430), .QN(n3073) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n4465), .CK(n4430), .QN(n3074) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n4466), .CK(n4430), .QN(n3075) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n4467), .CK(n4430), .QN(n3076) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n4468), .CK(n4430), .QN(n3077) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n4469), .CK(n4430), .QN(n3078) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n4470), .CK(n4430), .QN(n3079) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n4471), .CK(n4430), .QN(n3080) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n4472), .CK(n4430), .QN(n3081) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n4473), .CK(n4430), .QN(n3082) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n4474), .CK(n4430), .QN(n3083) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n4475), .CK(n4430), .QN(n3084) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n4476), .CK(n4430), .QN(n3085) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n4477), .CK(n4430), .QN(n3086) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n4478), .CK(n4430), .QN(n3087) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n4479), .CK(n4430), .QN(n3088) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n4480), .CK(n4430), .QN(n3089) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n4481), .CK(n4430), .QN(n3090) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n4482), .CK(n4430), .QN(n3091) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n4483), .CK(n4430), .QN(n3092) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n4484), .CK(n4430), .QN(n3093) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n4485), .CK(n4430), .QN(n3094) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n4486), .CK(n4430), .QN(n3095) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n4455), .CK(n4431), .QN(n3096) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n4456), .CK(n4431), .QN(n3097) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n4457), .CK(n4431), .QN(n3098) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n4458), .CK(n4431), .QN(n3099) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n4459), .CK(n4431), .QN(n3100) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n4460), .CK(n4431), .QN(n3101) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n4461), .CK(n4431), .QN(n3102) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n4462), .CK(n4431), .QN(n3103) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n4463), .CK(n4431), .QN(n3104) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n4464), .CK(n4431), .QN(n3105) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n4465), .CK(n4431), .QN(n3106) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n4466), .CK(n4431), .QN(n3107) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n4467), .CK(n4431), .QN(n3108) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n4468), .CK(n4431), .QN(n3109) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n4469), .CK(n4431), .QN(n3110) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n4470), .CK(n4431), .QN(n3111) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n4471), .CK(n4431), .QN(n3112) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n4472), .CK(n4431), .QN(n3113) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n4473), .CK(n4431), .QN(n3114) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n4474), .CK(n4431), .QN(n3115) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n4475), .CK(n4431), .QN(n3116) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n4476), .CK(n4431), .QN(n3117) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n4477), .CK(n4431), .QN(n3118) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n4478), .CK(n4431), .QN(n3119) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n4479), .CK(n4431), .QN(n3120) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n4480), .CK(n4431), .QN(n3121) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n4481), .CK(n4431), .QN(n3122) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n4482), .CK(n4431), .QN(n3123) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n4483), .CK(n4431), .QN(n3124) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n4484), .CK(n4431), .QN(n3125) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n4485), .CK(n4431), .QN(n3126) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n4486), .CK(n4431), .QN(n3127) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n4455), .CK(n4432), .QN(n3128) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n4456), .CK(n4432), .QN(n3129) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n4457), .CK(n4432), .QN(n3130) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n4458), .CK(n4432), .QN(n3131) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n4459), .CK(n4432), .QN(n3132) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n4460), .CK(n4432), .QN(n3133) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n4461), .CK(n4432), .QN(n3134) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n4462), .CK(n4432), .QN(n3135) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n4463), .CK(n4432), .QN(n3136) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n4464), .CK(n4432), .QN(n3137) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n4465), .CK(n4432), .QN(n3138) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n4466), .CK(n4432), .QN(n3139) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n4467), .CK(n4432), .QN(n3140) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n4468), .CK(n4432), .QN(n3141) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n4469), .CK(n4432), .QN(n3142) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n4470), .CK(n4432), .QN(n3143) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n4471), .CK(n4432), .QN(n3144) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n4472), .CK(n4432), .QN(n3145) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n4473), .CK(n4432), .QN(n3146) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n4474), .CK(n4432), .QN(n3147) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n4475), .CK(n4432), .QN(n3148) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n4476), .CK(n4432), .QN(n3149) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n4477), .CK(n4432), .QN(n3150) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n4478), .CK(n4432), .QN(n3151) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n4479), .CK(n4432), .QN(n3152) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n4480), .CK(n4432), .QN(n3153) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n4481), .CK(n4432), .QN(n3154) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n4482), .CK(n4432), .QN(n3155) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n4483), .CK(n4432), .QN(n3156) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n4484), .CK(n4432), .QN(n3157) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n4485), .CK(n4432), .QN(n3158) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n4486), .CK(n4432), .QN(n3159) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n4455), .CK(n4433), .QN(n3160) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n4456), .CK(n4433), .QN(n3161) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n4457), .CK(n4433), .QN(n3162) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n4458), .CK(n4433), .QN(n3163) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n4459), .CK(n4433), .QN(n3164) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n4460), .CK(n4433), .QN(n3165) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n4461), .CK(n4433), .QN(n3166) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n4462), .CK(n4433), .QN(n3167) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n4463), .CK(n4433), .QN(n3168) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n4464), .CK(n4433), .QN(n3169) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n4465), .CK(n4433), .QN(n3170) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n4466), .CK(n4433), .QN(n3171) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n4467), .CK(n4433), .QN(n3172) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n4468), .CK(n4433), .QN(n3173) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n4469), .CK(n4433), .QN(n3174) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n4470), .CK(n4433), .QN(n3175) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n4471), .CK(n4433), .QN(n3176) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n4472), .CK(n4433), .QN(n3177) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n4473), .CK(n4433), .QN(n3178) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n4474), .CK(n4433), .QN(n3179) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n4475), .CK(n4433), .QN(n3180) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n4476), .CK(n4433), .QN(n3181) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n4477), .CK(n4433), .QN(n3182) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n4478), .CK(n4433), .QN(n3183) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n4479), .CK(n4433), .QN(n3184) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n4480), .CK(n4433), .QN(n3185) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n4481), .CK(n4433), .QN(n3186) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n4482), .CK(n4433), .QN(n3187) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n4483), .CK(n4433), .QN(n3188) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n4484), .CK(n4433), .QN(n3189) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n4485), .CK(n4433), .QN(n3190) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n4486), .CK(n4433), .QN(n3191) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n4455), .CK(n4434), .QN(n3192) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n4456), .CK(n4434), .QN(n3193) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n4457), .CK(n4434), .QN(n3194) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n4458), .CK(n4434), .QN(n3195) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n4459), .CK(n4434), .QN(n3196) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n4460), .CK(n4434), .QN(n3197) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n4461), .CK(n4434), .QN(n3198) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n4462), .CK(n4434), .QN(n3199) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n4463), .CK(n4434), .QN(n3200) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n4464), .CK(n4434), .QN(n3201) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n4465), .CK(n4434), .QN(n3202) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n4466), .CK(n4434), .QN(n3203) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n4467), .CK(n4434), .QN(n3204) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n4468), .CK(n4434), .QN(n3205) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n4469), .CK(n4434), .QN(n3206) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n4470), .CK(n4434), .QN(n3207) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n4471), .CK(n4434), .QN(n3208) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n4472), .CK(n4434), .QN(n3209) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n4473), .CK(n4434), .QN(n3210) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n4474), .CK(n4434), .QN(n3211) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n4475), .CK(n4434), .QN(n3212) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n4476), .CK(n4434), .QN(n3213) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n4477), .CK(n4434), .QN(n3214) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n4478), .CK(n4434), .QN(n3215) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n4479), .CK(n4434), .QN(n3216) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n4480), .CK(n4434), .QN(n3217) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n4481), .CK(n4434), .QN(n3218) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n4482), .CK(n4434), .QN(n3219) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n4483), .CK(n4434), .QN(n3220) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n4484), .CK(n4434), .QN(n3221) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n4485), .CK(n4434), .QN(n3222) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n4486), .CK(n4434), .QN(n3223) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n4455), .CK(n4436), .QN(n3224) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n4456), .CK(n4436), .QN(n3225) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n4457), .CK(n4436), .QN(n3226) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n4458), .CK(n4436), .QN(n3227) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n4459), .CK(n4436), .QN(n3228) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n4460), .CK(n4436), .QN(n3229) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n4461), .CK(n4436), .QN(n3230) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n4462), .CK(n4436), .QN(n3231) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n4463), .CK(n4436), .QN(n3232) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n4464), .CK(n4436), .QN(n3233) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n4465), .CK(n4436), .QN(n3234) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n4466), .CK(n4436), .QN(n3235) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n4467), .CK(n4436), .QN(n3236) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n4468), .CK(n4436), .QN(n3237) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n4469), .CK(n4436), .QN(n3238) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n4470), .CK(n4436), .QN(n3239) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n4471), .CK(n4436), .QN(n3240) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n4472), .CK(n4436), .QN(n3241) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n4473), .CK(n4436), .QN(n3242) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n4474), .CK(n4436), .QN(n3243) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n4475), .CK(n4436), .QN(n3244) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n4476), .CK(n4436), .QN(n3245) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n4477), .CK(n4436), .QN(n3246) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n4478), .CK(n4436), .QN(n3247) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n4479), .CK(n4436), .QN(n3248) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n4480), .CK(n4436), .QN(n3249) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n4481), .CK(n4436), .QN(n3250) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n4482), .CK(n4436), .QN(n3251) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n4483), .CK(n4436), .QN(n3252) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n4484), .CK(n4436), .QN(n3253) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n4485), .CK(n4436), .QN(n3254) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n4486), .CK(n4436), .QN(n3255) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n4455), .CK(n4437), .QN(n3256) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n4456), .CK(n4437), .QN(n3257) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n4457), .CK(n4437), .QN(n3258) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n4458), .CK(n4437), .QN(n3259) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n4459), .CK(n4437), .QN(n3260) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n4460), .CK(n4437), .QN(n3261) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n4461), .CK(n4437), .QN(n3262) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n4462), .CK(n4437), .QN(n3263) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n4463), .CK(n4437), .QN(n3264) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n4464), .CK(n4437), .QN(n3265) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n4465), .CK(n4437), .QN(n3266) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n4466), .CK(n4437), .QN(n3267) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n4467), .CK(n4437), .QN(n3268) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n4468), .CK(n4437), .QN(n3269) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n4469), .CK(n4437), .QN(n3270) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n4470), .CK(n4437), .QN(n3271) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n4471), .CK(n4437), .QN(n3272) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n4472), .CK(n4437), .QN(n3273) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n4473), .CK(n4437), .QN(n3274) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n4474), .CK(n4437), .QN(n3275) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n4475), .CK(n4437), .QN(n3276) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n4476), .CK(n4437), .QN(n3277) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n4477), .CK(n4437), .QN(n3278) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n4478), .CK(n4437), .QN(n3279) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n4479), .CK(n4437), .QN(n3280) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n4480), .CK(n4437), .QN(n3281) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n4481), .CK(n4437), .QN(n3282) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n4482), .CK(n4437), .QN(n3283) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n4483), .CK(n4437), .QN(n3284) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n4484), .CK(n4437), .QN(n3285) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n4485), .CK(n4437), .QN(n3286) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n4486), .CK(n4437), .QN(n3287) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n4455), .CK(n4438), .QN(n3288) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n4456), .CK(n4438), .QN(n3289) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n4457), .CK(n4438), .QN(n3290) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n4458), .CK(n4438), .QN(n3291) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n4459), .CK(n4438), .QN(n3292) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n4460), .CK(n4438), .QN(n3293) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n4461), .CK(n4438), .QN(n3294) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n4462), .CK(n4438), .QN(n3295) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n4463), .CK(n4438), .QN(n3296) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n4464), .CK(n4438), .QN(n3297) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n4465), .CK(n4438), .QN(n3298) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n4466), .CK(n4438), .QN(n3299) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n4467), .CK(n4438), .QN(n3300) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n4468), .CK(n4438), .QN(n3301) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n4469), .CK(n4438), .QN(n3302) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n4470), .CK(n4438), .QN(n3303) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n4471), .CK(n4438), .QN(n3304) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n4472), .CK(n4438), .QN(n3305) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n4473), .CK(n4438), .QN(n3306) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n4474), .CK(n4438), .QN(n3307) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n4475), .CK(n4438), .QN(n3308) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n4476), .CK(n4438), .QN(n3309) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n4477), .CK(n4438), .QN(n3310) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n4478), .CK(n4438), .QN(n3311) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n4479), .CK(n4438), .QN(n3312) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n4480), .CK(n4438), .QN(n3313) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n4481), .CK(n4438), .QN(n3314) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n4482), .CK(n4438), .QN(n3315) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n4483), .CK(n4438), .QN(n3316) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n4484), .CK(n4438), .QN(n3317) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n4485), .CK(n4438), .QN(n3318) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n4486), .CK(n4438), .QN(n3319) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n4455), .CK(n4439), .QN(n3320) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n4456), .CK(n4439), .QN(n3321) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n4457), .CK(n4439), .QN(n3322) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n4458), .CK(n4439), .QN(n3323) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n4459), .CK(n4439), .QN(n3324) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n4460), .CK(n4439), .QN(n3325) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n4461), .CK(n4439), .QN(n3326) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n4462), .CK(n4439), .QN(n3327) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n4463), .CK(n4439), .QN(n3328) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n4464), .CK(n4439), .QN(n3329) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n4465), .CK(n4439), .QN(n3330) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n4466), .CK(n4439), .QN(n3331) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n4467), .CK(n4439), .QN(n3332) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n4468), .CK(n4439), .QN(n3333) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n4469), .CK(n4439), .QN(n3334) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n4470), .CK(n4439), .QN(n3335) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n4471), .CK(n4439), .QN(n3336) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n4472), .CK(n4439), .QN(n3337) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n4473), .CK(n4439), .QN(n3338) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n4474), .CK(n4439), .QN(n3339) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n4475), .CK(n4439), .QN(n3340) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n4476), .CK(n4439), .QN(n3341) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n4477), .CK(n4439), .QN(n3342) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n4478), .CK(n4439), .QN(n3343) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n4479), .CK(n4439), .QN(n3344) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n4480), .CK(n4439), .QN(n3345) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n4481), .CK(n4439), .QN(n3346) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n4482), .CK(n4439), .QN(n3347) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n4483), .CK(n4439), .QN(n3348) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n4484), .CK(n4439), .QN(n3349) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n4485), .CK(n4439), .QN(n3350) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n4486), .CK(n4439), .QN(n3351) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n4455), .CK(n4440), .QN(n3352) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n4456), .CK(n4440), .QN(n3353) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n4457), .CK(n4440), .QN(n3354) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n4458), .CK(n4440), .QN(n3355) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n4459), .CK(n4440), .QN(n3356) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n4460), .CK(n4440), .QN(n3357) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n4461), .CK(n4440), .QN(n3358) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n4462), .CK(n4440), .QN(n3359) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n4463), .CK(n4440), .QN(n3360) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n4464), .CK(n4440), .QN(n3361) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n4465), .CK(n4440), .QN(n3362) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n4466), .CK(n4440), .QN(n3363) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n4467), .CK(n4440), .QN(n3364) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n4468), .CK(n4440), .QN(n3365) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n4469), .CK(n4440), .QN(n3366) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n4470), .CK(n4440), .QN(n3367) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n4471), .CK(n4440), .QN(n3368) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n4472), .CK(n4440), .QN(n3369) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n4473), .CK(n4440), .QN(n3370) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n4474), .CK(n4440), .QN(n3371) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n4475), .CK(n4440), .QN(n3372) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n4476), .CK(n4440), .QN(n3373) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n4477), .CK(n4440), .QN(n3374) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n4478), .CK(n4440), .QN(n3375) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n4479), .CK(n4440), .QN(n3376) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n4480), .CK(n4440), .QN(n3377) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n4481), .CK(n4440), .QN(n3378) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n4482), .CK(n4440), .QN(n3379) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n4483), .CK(n4440), .QN(n3380) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n4484), .CK(n4440), .QN(n3381) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n4485), .CK(n4440), .QN(n3382) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n4486), .CK(n4440), .QN(n3383) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n4455), .CK(n4441), .QN(n3384) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n4456), .CK(n4441), .QN(n3385) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n4457), .CK(n4441), .QN(n3386) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n4458), .CK(n4441), .QN(n3387) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n4459), .CK(n4441), .QN(n3388) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n4460), .CK(n4441), .QN(n3389) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n4461), .CK(n4441), .QN(n3390) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n4462), .CK(n4441), .QN(n3391) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n4463), .CK(n4441), .QN(n3392) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n4464), .CK(n4441), .QN(n3393) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n4465), .CK(n4441), .QN(n3394) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n4466), .CK(n4441), .QN(n3395) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n4467), .CK(n4441), .QN(n3396) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n4468), .CK(n4441), .QN(n3397) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n4469), .CK(n4441), .QN(n3398) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n4470), .CK(n4441), .QN(n3399) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n4471), .CK(n4441), .QN(n3400) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n4472), .CK(n4441), .QN(n3401) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n4473), .CK(n4441), .QN(n3402) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n4474), .CK(n4441), .QN(n3403) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n4475), .CK(n4441), .QN(n3404) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n4476), .CK(n4441), .QN(n3405) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n4477), .CK(n4441), .QN(n3406) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n4478), .CK(n4441), .QN(n3407) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n4479), .CK(n4441), .QN(n3408) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n4480), .CK(n4441), .QN(n3409) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n4481), .CK(n4441), .QN(n3410) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n4482), .CK(n4441), .QN(n3411) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n4483), .CK(n4441), .QN(n3412) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n4484), .CK(n4441), .QN(n3413) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n4485), .CK(n4441), .QN(n3414) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n4486), .CK(n4441), .QN(n3415) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n4455), .CK(n4442), .QN(n3416) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n4456), .CK(n4442), .QN(n3417) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n4457), .CK(n4442), .QN(n3418) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n4458), .CK(n4442), .QN(n3419) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n4459), .CK(n4442), .QN(n3420) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n4460), .CK(n4442), .QN(n3421) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n4461), .CK(n4442), .QN(n3422) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n4462), .CK(n4442), .QN(n3423) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n4463), .CK(n4442), .QN(n3424) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n4464), .CK(n4442), .QN(n3425) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n4465), .CK(n4442), .QN(n3426) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n4466), .CK(n4442), .QN(n3427) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n4467), .CK(n4442), .QN(n3428) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n4468), .CK(n4442), .QN(n3429) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n4469), .CK(n4442), .QN(n3430) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n4470), .CK(n4442), .QN(n3431) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n4471), .CK(n4442), .QN(n3432) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n4472), .CK(n4442), .QN(n3433) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n4473), .CK(n4442), .QN(n3434) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n4474), .CK(n4442), .QN(n3435) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n4475), .CK(n4442), .QN(n3436) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n4476), .CK(n4442), .QN(n3437) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n4477), .CK(n4442), .QN(n3438) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n4478), .CK(n4442), .QN(n3439) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n4479), .CK(n4442), .QN(n3440) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n4480), .CK(n4442), .QN(n3441) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n4481), .CK(n4442), .QN(n3442) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n4482), .CK(n4442), .QN(n3443) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n4483), .CK(n4442), .QN(n3444) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n4484), .CK(n4442), .QN(n3445) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n4485), .CK(n4442), .QN(n3446) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n4486), .CK(n4442), .QN(n3447) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n4455), .CK(n4443), .QN(n3448) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n4456), .CK(n4443), .QN(n3449) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n4457), .CK(n4443), .QN(n3450) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n4458), .CK(n4443), .QN(n3451) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n4459), .CK(n4443), .QN(n3452) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n4460), .CK(n4443), .QN(n3453) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n4461), .CK(n4443), .QN(n3454) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n4462), .CK(n4443), .QN(n3455) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n4463), .CK(n4443), .QN(n3456) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n4464), .CK(n4443), .QN(n3457) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n4465), .CK(n4443), .QN(n3458) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n4466), .CK(n4443), .QN(n3459) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n4467), .CK(n4443), .QN(n3460) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n4468), .CK(n4443), .QN(n3461) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n4469), .CK(n4443), .QN(n3462) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n4470), .CK(n4443), .QN(n3463) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n4471), .CK(n4443), .QN(n3464) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n4472), .CK(n4443), .QN(n3465) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n4473), .CK(n4443), .QN(n3466) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n4474), .CK(n4443), .QN(n3467) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n4475), .CK(n4443), .QN(n3468) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n4476), .CK(n4443), .QN(n3469) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n4477), .CK(n4443), .QN(n3470) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n4478), .CK(n4443), .QN(n3471) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n4479), .CK(n4443), .QN(n3472) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n4480), .CK(n4443), .QN(n3473) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n4481), .CK(n4443), .QN(n3474) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n4482), .CK(n4443), .QN(n3475) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n4483), .CK(n4443), .QN(n3476) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n4484), .CK(n4443), .QN(n3477) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n4485), .CK(n4443), .QN(n3478) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n4486), .CK(n4443), .QN(n3479) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n4455), .CK(n4444), .QN(n3480) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n4456), .CK(n4444), .QN(n3481) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n4457), .CK(n4444), .QN(n3482) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n4458), .CK(n4444), .QN(n3483) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n4459), .CK(n4444), .QN(n3484) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n4460), .CK(n4444), .QN(n3485) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n4461), .CK(n4444), .QN(n3486) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n4462), .CK(n4444), .QN(n3487) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n4463), .CK(n4444), .QN(n3488) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n4464), .CK(n4444), .QN(n3489) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n4465), .CK(n4444), .QN(n3490) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n4466), .CK(n4444), .QN(n3491) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n4467), .CK(n4444), .QN(n3492) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n4468), .CK(n4444), .QN(n3493) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n4469), .CK(n4444), .QN(n3494) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n4470), .CK(n4444), .QN(n3495) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n4471), .CK(n4444), .QN(n3496) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n4472), .CK(n4444), .QN(n3497) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n4473), .CK(n4444), .QN(n3498) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n4474), .CK(n4444), .QN(n3499) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n4475), .CK(n4444), .QN(n3500) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n4476), .CK(n4444), .QN(n3501) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n4477), .CK(n4444), .QN(n3502) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n4478), .CK(n4444), .QN(n3503) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n4479), .CK(n4444), .QN(n3504) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n4480), .CK(n4444), .QN(n3505) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n4481), .CK(n4444), .QN(n3506) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n4482), .CK(n4444), .QN(n3507) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n4483), .CK(n4444), .QN(n3508) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n4484), .CK(n4444), .QN(n3509) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n4485), .CK(n4444), .QN(n3510) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n4486), .CK(n4444), .QN(n3511) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n4455), .CK(n4445), .QN(n3512) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n4456), .CK(n4445), .QN(n3513) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n4457), .CK(n4445), .QN(n3514) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n4458), .CK(n4445), .QN(n3515) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n4459), .CK(n4445), .QN(n3516) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n4460), .CK(n4445), .QN(n3517) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n4461), .CK(n4445), .QN(n3518) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n4462), .CK(n4445), .QN(n3519) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n4463), .CK(n4445), .QN(n3520) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n4464), .CK(n4445), .QN(n3521) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n4465), .CK(n4445), .QN(n3522) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n4466), .CK(n4445), .QN(n3523) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n4467), .CK(n4445), .QN(n3524) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n4468), .CK(n4445), .QN(n3525) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n4469), .CK(n4445), .QN(n3526) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n4470), .CK(n4445), .QN(n3527) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n4471), .CK(n4445), .QN(n3528) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n4472), .CK(n4445), .QN(n3529) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n4473), .CK(n4445), .QN(n3530) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n4474), .CK(n4445), .QN(n3531) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n4475), .CK(n4445), .QN(n3532) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n4476), .CK(n4445), .QN(n3533) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n4477), .CK(n4445), .QN(n3534) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n4478), .CK(n4445), .QN(n3535) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n4479), .CK(n4445), .QN(n3536) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n4480), .CK(n4445), .QN(n3537) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n4481), .CK(n4445), .QN(n3538) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n4482), .CK(n4445), .QN(n3539) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n4483), .CK(n4445), .QN(n3540) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n4484), .CK(n4445), .QN(n3541) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n4485), .CK(n4445), .QN(n3542) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n4486), .CK(n4445), .QN(n3543) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n4455), .CK(n4447), .QN(n3544) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n4456), .CK(n4447), .QN(n3545) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n4457), .CK(n4447), .QN(n3546) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n4458), .CK(n4447), .QN(n3547) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n4459), .CK(n4447), .QN(n3548) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n4460), .CK(n4447), .QN(n3549) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n4461), .CK(n4447), .QN(n3550) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n4462), .CK(n4447), .QN(n3551) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n4463), .CK(n4447), .QN(n3552) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n4464), .CK(n4447), .QN(n3553) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n4465), .CK(n4447), .QN(n3554) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n4466), .CK(n4447), .QN(n3555) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n4467), .CK(n4447), .QN(n3556) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n4468), .CK(n4447), .QN(n3557) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n4469), .CK(n4447), .QN(n3558) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n4470), .CK(n4447), .QN(n3559) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n4471), .CK(n4447), .QN(n3560) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n4472), .CK(n4447), .QN(n3561) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n4473), .CK(n4447), .QN(n3562) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n4474), .CK(n4447), .QN(n3563) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n4475), .CK(n4447), .QN(n3564) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n4476), .CK(n4447), .QN(n3565) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n4477), .CK(n4447), .QN(n3566) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n4478), .CK(n4447), .QN(n3567) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n4479), .CK(n4447), .QN(n3568) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n4480), .CK(n4447), .QN(n3569) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n4481), .CK(n4447), .QN(n3570) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n4482), .CK(n4447), .QN(n3571) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n4483), .CK(n4447), .QN(n3572) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n4484), .CK(n4447), .QN(n3573) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n4485), .CK(n4447), .QN(n3574) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n4486), .CK(n4447), .QN(n3575) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n4455), .CK(n4448), .QN(n3576) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n4456), .CK(n4448), .QN(n3577) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n4457), .CK(n4448), .QN(n3578) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n4458), .CK(n4448), .QN(n3579) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n4459), .CK(n4448), .QN(n3580) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n4460), .CK(n4448), .QN(n3581) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n4461), .CK(n4448), .QN(n3582) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n4462), .CK(n4448), .QN(n3583) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n4463), .CK(n4448), .QN(n3584) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n4464), .CK(n4448), .QN(n3585) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n4465), .CK(n4448), .QN(n3586) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n4466), .CK(n4448), .QN(n3587) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n4467), .CK(n4448), .QN(n3588) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n4468), .CK(n4448), .QN(n3589) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n4469), .CK(n4448), .QN(n3590) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n4470), .CK(n4448), .QN(n3591) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n4471), .CK(n4448), .QN(n3592) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n4472), .CK(n4448), .QN(n3593) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n4473), .CK(n4448), .QN(n3594) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n4474), .CK(n4448), .QN(n3595) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n4475), .CK(n4448), .QN(n3596) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n4476), .CK(n4448), .QN(n3597) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n4477), .CK(n4448), .QN(n3598) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n4478), .CK(n4448), .QN(n3599) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n4479), .CK(n4448), .QN(n3600) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n4480), .CK(n4448), .QN(n3601) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n4481), .CK(n4448), .QN(n3602) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n4482), .CK(n4448), .QN(n3603) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n4483), .CK(n4448), .QN(n3604) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n4484), .CK(n4448), .QN(n3605) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n4485), .CK(n4448), .QN(n3606) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n4486), .CK(n4448), .QN(n3607) );
  DLH_X1 \OUT1_reg[31]  ( .G(N444), .D(N410), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N444), .D(N409), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N444), .D(N408), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N444), .D(N407), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N444), .D(N406), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N444), .D(N405), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N444), .D(N404), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N444), .D(N403), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N444), .D(N402), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N444), .D(N401), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N444), .D(N400), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N444), .D(N399), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N444), .D(N398), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N444), .D(N397), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N444), .D(N396), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N444), .D(N395), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N444), .D(N394), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N444), .D(N393), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N444), .D(N392), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N444), .D(N391), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N444), .D(N390), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N444), .D(N389), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N444), .D(N388), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N444), .D(N387), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N444), .D(N386), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N444), .D(N385), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N444), .D(N384), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N444), .D(N383), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N444), .D(N382), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N444), .D(N381), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N444), .D(N380), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N444), .D(N379), .Q(OUT1[0]) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_0 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(n10), .ENCLK(n4487), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_1 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(n9), .ENCLK(n4454), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_2 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(n8), .ENCLK(n4453), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_3 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(n7), .ENCLK(n4452), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_4 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(n6), .ENCLK(n4451), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_5 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(n5), .ENCLK(n4450), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_6 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(n4), .ENCLK(n4449), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_7 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(n33), .ENCLK(n4448), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_8 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(n31), .ENCLK(n4447), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_9 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(n3), .ENCLK(n4446), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_10 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(n30), .ENCLK(n4445), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_11 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(n29), .ENCLK(n4444), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_12 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(n28), .ENCLK(n4443), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_13 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(n27), .ENCLK(n4442), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_14 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(n26), .ENCLK(n4441), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_15 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(n25), .ENCLK(n4440), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_16 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(n24), .ENCLK(n4439), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_17 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(n23), .ENCLK(n4438), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_18 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(n22), .ENCLK(n4437), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_19 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(n21), .ENCLK(n4436), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_20 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(n2), .ENCLK(n4435), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_21 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(n20), .ENCLK(n4434), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_22 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(n19), .ENCLK(n4433), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_23 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(n18), .ENCLK(n4432), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_24 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(n17), .ENCLK(n4431), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_25 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(n16), .ENCLK(n4430), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_26 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(n15), .ENCLK(n4429), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_27 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(n14), .ENCLK(n4428), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_28 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(n13), .ENCLK(n4427), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_29 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(n12), .ENCLK(n4426), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_30 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(n11), .ENCLK(n4425), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_register_file_WORD_SIZE32_ADDR_SIZE5_31 \clk_gate_REGISTERS_reg[0]  ( 
        .CLK(CLK), .EN(n1), .ENCLK(n4423), .TE(1'b0) );
  INV_X1 U3 ( .A(RESET), .ZN(n3623) );
  INV_X1 U4 ( .A(RESET), .ZN(n3669) );
  INV_X1 U5 ( .A(RESET), .ZN(n3668) );
  INV_X1 U6 ( .A(RESET), .ZN(n3616) );
  INV_X1 U7 ( .A(RESET), .ZN(n3617) );
  INV_X1 U8 ( .A(RESET), .ZN(n3663) );
  INV_X1 U9 ( .A(RESET), .ZN(n3664) );
  INV_X1 U10 ( .A(RESET), .ZN(n3618) );
  INV_X1 U11 ( .A(RESET), .ZN(n3665) );
  INV_X1 U12 ( .A(RESET), .ZN(n3619) );
  INV_X1 U13 ( .A(RESET), .ZN(n3620) );
  INV_X1 U14 ( .A(RESET), .ZN(n3671) );
  INV_X1 U15 ( .A(RESET), .ZN(n3666) );
  INV_X1 U16 ( .A(RESET), .ZN(n3621) );
  INV_X1 U17 ( .A(RESET), .ZN(n3622) );
  INV_X1 U18 ( .A(RESET), .ZN(n3667) );
  INV_X1 U19 ( .A(RESET), .ZN(n3656) );
  INV_X1 U20 ( .A(RESET), .ZN(n3657) );
  INV_X1 U21 ( .A(RESET), .ZN(n3658) );
  INV_X1 U22 ( .A(RESET), .ZN(n3659) );
  INV_X1 U23 ( .A(RESET), .ZN(n3660) );
  INV_X1 U24 ( .A(RESET), .ZN(n3661) );
  INV_X1 U25 ( .A(RESET), .ZN(n3670) );
  INV_X1 U26 ( .A(RESET), .ZN(n3662) );
  INV_X1 U27 ( .A(RESET), .ZN(n3646) );
  INV_X1 U28 ( .A(RESET), .ZN(n3645) );
  INV_X1 U29 ( .A(RESET), .ZN(n3644) );
  INV_X1 U30 ( .A(RESET), .ZN(n3643) );
  INV_X1 U31 ( .A(RESET), .ZN(n3642) );
  INV_X1 U32 ( .A(RESET), .ZN(n3636) );
  INV_X1 U33 ( .A(RESET), .ZN(n3626) );
  INV_X1 U34 ( .A(RESET), .ZN(n3637) );
  INV_X1 U35 ( .A(RESET), .ZN(n3638) );
  INV_X1 U36 ( .A(RESET), .ZN(n3635) );
  INV_X1 U37 ( .A(RESET), .ZN(n3632) );
  INV_X1 U38 ( .A(RESET), .ZN(n3633) );
  INV_X1 U39 ( .A(RESET), .ZN(n3634) );
  INV_X1 U40 ( .A(RESET), .ZN(n3631) );
  INV_X1 U41 ( .A(RESET), .ZN(n3627) );
  INV_X1 U42 ( .A(RESET), .ZN(n3628) );
  INV_X1 U43 ( .A(RESET), .ZN(n3630) );
  INV_X1 U44 ( .A(RESET), .ZN(n3625) );
  INV_X1 U45 ( .A(RESET), .ZN(n3629) );
  INV_X1 U46 ( .A(RESET), .ZN(n3655) );
  INV_X1 U47 ( .A(RESET), .ZN(n3654) );
  INV_X1 U48 ( .A(RESET), .ZN(n3641) );
  INV_X1 U49 ( .A(RESET), .ZN(n3650) );
  INV_X1 U50 ( .A(RESET), .ZN(n3647) );
  INV_X1 U51 ( .A(RESET), .ZN(n3640) );
  INV_X1 U52 ( .A(RESET), .ZN(n3639) );
  INV_X1 U53 ( .A(RESET), .ZN(n3648) );
  INV_X1 U54 ( .A(RESET), .ZN(n3649) );
  INV_X1 U55 ( .A(RESET), .ZN(n3651) );
  INV_X1 U56 ( .A(RESET), .ZN(n3652) );
  INV_X1 U57 ( .A(RESET), .ZN(n3653) );
  INV_X1 U58 ( .A(RESET), .ZN(n3624) );
  INV_X1 U59 ( .A(RESET), .ZN(n3608) );
  OAI21_X1 U60 ( .B1(n4414), .B2(n4408), .A(n3608), .ZN(n33) );
  INV_X1 U61 ( .A(RESET), .ZN(n3609) );
  OAI21_X1 U62 ( .B1(n4418), .B2(n4421), .A(n3609), .ZN(n4) );
  INV_X1 U63 ( .A(RESET), .ZN(n3610) );
  OAI21_X1 U64 ( .B1(n4417), .B2(n4421), .A(n3610), .ZN(n5) );
  INV_X1 U65 ( .A(RESET), .ZN(n3611) );
  OAI21_X1 U66 ( .B1(n4416), .B2(n4421), .A(n3611), .ZN(n6) );
  INV_X1 U67 ( .A(RESET), .ZN(n3612) );
  OAI21_X1 U68 ( .B1(n4415), .B2(n4421), .A(n3612), .ZN(n7) );
  INV_X1 U69 ( .A(RESET), .ZN(n3613) );
  OAI21_X1 U70 ( .B1(n4414), .B2(n4421), .A(n3613), .ZN(n8) );
  INV_X1 U71 ( .A(RESET), .ZN(n3614) );
  OAI21_X1 U72 ( .B1(n4422), .B2(n4410), .A(n3614), .ZN(n9) );
  INV_X1 U73 ( .A(RESET), .ZN(n3615) );
  OAI21_X1 U74 ( .B1(n4420), .B2(n4410), .A(n3615), .ZN(n10) );
  AND2_X1 U75 ( .A1(n3642), .A2(DATAIN[4]), .ZN(n4482) );
  AND2_X1 U76 ( .A1(n3643), .A2(DATAIN[3]), .ZN(n4483) );
  AND2_X1 U77 ( .A1(n3644), .A2(DATAIN[2]), .ZN(n4484) );
  AND2_X1 U78 ( .A1(n3645), .A2(DATAIN[1]), .ZN(n4485) );
  AND2_X1 U79 ( .A1(n3646), .A2(DATAIN[0]), .ZN(n4486) );
  AND2_X1 U80 ( .A1(n3647), .A2(DATAIN[23]), .ZN(n4463) );
  AND2_X1 U81 ( .A1(n3648), .A2(DATAIN[26]), .ZN(n4460) );
  AND2_X1 U82 ( .A1(n3649), .A2(DATAIN[27]), .ZN(n4459) );
  AND2_X1 U83 ( .A1(n3650), .A2(DATAIN[22]), .ZN(n4464) );
  AND2_X1 U84 ( .A1(n3651), .A2(DATAIN[28]), .ZN(n4458) );
  AND2_X1 U85 ( .A1(n3652), .A2(DATAIN[29]), .ZN(n4457) );
  AND2_X1 U86 ( .A1(n3653), .A2(DATAIN[30]), .ZN(n4456) );
  AND2_X1 U87 ( .A1(n3654), .A2(DATAIN[20]), .ZN(n4466) );
  AND2_X1 U88 ( .A1(n3655), .A2(DATAIN[19]), .ZN(n4467) );
  INV_X2 U89 ( .A(n3708), .ZN(n4391) );
  INV_X2 U90 ( .A(n3710), .ZN(n4393) );
  INV_X2 U91 ( .A(n3709), .ZN(n4390) );
  INV_X2 U92 ( .A(n3706), .ZN(n4388) );
  INV_X2 U93 ( .A(n3707), .ZN(n4389) );
  NAND2_X2 U94 ( .A1(n3673), .A2(n3701), .ZN(n4368) );
  NAND2_X2 U95 ( .A1(n3710), .A2(n3699), .ZN(n4376) );
  NAND2_X2 U96 ( .A1(n3707), .A2(n3701), .ZN(n4363) );
  NAND2_X2 U97 ( .A1(n3709), .A2(n3700), .ZN(n4375) );
  NAND2_X2 U98 ( .A1(n3707), .A2(n3700), .ZN(n4364) );
  NAND2_X2 U99 ( .A1(n3709), .A2(n3701), .ZN(n4378) );
  NAND2_X2 U100 ( .A1(n3673), .A2(n3699), .ZN(n4357) );
  NAND2_X2 U101 ( .A1(n3711), .A2(n3699), .ZN(n4377) );
  NAND2_X2 U102 ( .A1(n3707), .A2(n3699), .ZN(n4356) );
  NAND2_X2 U103 ( .A1(n3710), .A2(n3701), .ZN(n4379) );
  NAND2_X2 U104 ( .A1(n3706), .A2(n3701), .ZN(n4354) );
  NAND2_X2 U105 ( .A1(n3706), .A2(n3700), .ZN(n4351) );
  NAND2_X2 U106 ( .A1(n3710), .A2(n3700), .ZN(n4380) );
  NAND2_X2 U107 ( .A1(n3711), .A2(n3700), .ZN(n4382) );
  NAND2_X2 U108 ( .A1(n3706), .A2(n3699), .ZN(n4352) );
  INV_X2 U109 ( .A(n3673), .ZN(n3672) );
  INV_X2 U110 ( .A(n3711), .ZN(n4392) );
  AND2_X1 U111 ( .A1(ENABLE), .A2(WR), .ZN(n4413) );
  AND2_X1 U112 ( .A1(n3641), .A2(DATAIN[21]), .ZN(n4465) );
  AND2_X1 U113 ( .A1(n3640), .A2(DATAIN[24]), .ZN(n4462) );
  AND2_X1 U114 ( .A1(n3639), .A2(DATAIN[25]), .ZN(n4461) );
  AND2_X1 U115 ( .A1(n3638), .A2(DATAIN[8]), .ZN(n4478) );
  AND2_X1 U116 ( .A1(n3637), .A2(DATAIN[7]), .ZN(n4479) );
  AND2_X1 U117 ( .A1(n3636), .A2(DATAIN[5]), .ZN(n4481) );
  AND2_X1 U118 ( .A1(n3635), .A2(DATAIN[9]), .ZN(n4477) );
  AND2_X1 U119 ( .A1(n3634), .A2(DATAIN[12]), .ZN(n4474) );
  AND2_X1 U120 ( .A1(n3633), .A2(DATAIN[11]), .ZN(n4475) );
  AND2_X1 U121 ( .A1(n3632), .A2(DATAIN[10]), .ZN(n4476) );
  AND2_X1 U122 ( .A1(n3631), .A2(DATAIN[13]), .ZN(n4473) );
  AND2_X1 U123 ( .A1(n3630), .A2(DATAIN[16]), .ZN(n4470) );
  AND2_X1 U124 ( .A1(n3629), .A2(DATAIN[18]), .ZN(n4468) );
  AND2_X1 U125 ( .A1(n3628), .A2(DATAIN[15]), .ZN(n4471) );
  AND2_X1 U126 ( .A1(n3627), .A2(DATAIN[14]), .ZN(n4472) );
  AND2_X1 U127 ( .A1(n3626), .A2(DATAIN[6]), .ZN(n4480) );
  AND2_X1 U128 ( .A1(n3625), .A2(DATAIN[17]), .ZN(n4469) );
  AND2_X1 U129 ( .A1(n3624), .A2(DATAIN[31]), .ZN(n4455) );
  INV_X1 U130 ( .A(ADD_WR[2]), .ZN(n4406) );
  AND2_X1 U131 ( .A1(ENABLE), .A2(RD1), .ZN(N444) );
  BUF_X1 U132 ( .A(n4381), .Z(n3682) );
  BUF_X1 U133 ( .A(n4369), .Z(n3680) );
  BUF_X1 U134 ( .A(n4370), .Z(n3681) );
  BUF_X1 U135 ( .A(n4367), .Z(n3679) );
  BUF_X1 U136 ( .A(n4365), .Z(n3677) );
  BUF_X1 U137 ( .A(n4366), .Z(n3678) );
  BUF_X1 U138 ( .A(n4358), .Z(n3676) );
  BUF_X1 U139 ( .A(n4355), .Z(n3675) );
  BUF_X1 U140 ( .A(n4353), .Z(n3674) );
  BUF_X1 U141 ( .A(n4399), .Z(n3685) );
  NOR2_X1 U142 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[0]), .ZN(n4399) );
  AND3_X1 U143 ( .A1(n3698), .A2(n3693), .A3(ADD_RD1[2]), .ZN(n3673) );
  INV_X1 U144 ( .A(n4387), .ZN(n3684) );
  INV_X1 U145 ( .A(ADD_RD1[3]), .ZN(n3698) );
  NOR2_X1 U146 ( .A1(ADD_RD1[1]), .A2(n3687), .ZN(n3701) );
  NOR2_X1 U147 ( .A1(ADD_RD1[0]), .A2(n3686), .ZN(n3700) );
  NOR2_X1 U148 ( .A1(n3686), .A2(n3687), .ZN(n3699) );
  INV_X1 U149 ( .A(n3684), .ZN(n3683) );
  NAND2_X1 U151 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[2]), .ZN(n3688) );
  INV_X1 U152 ( .A(ADD_RD1[4]), .ZN(n3693) );
  NOR2_X1 U153 ( .A1(n3688), .A2(n3693), .ZN(n3706) );
  INV_X1 U154 ( .A(ADD_RD1[1]), .ZN(n3686) );
  INV_X1 U155 ( .A(ADD_RD1[0]), .ZN(n3687) );
  OAI22_X1 U156 ( .A1(n3607), .A2(n4352), .B1(n3575), .B2(n4351), .ZN(n3692)
         );
  NAND3_X1 U157 ( .A1(n3698), .A2(ADD_RD1[2]), .A3(ADD_RD1[4]), .ZN(n4387) );
  NAND2_X1 U158 ( .A1(n3684), .A2(n3699), .ZN(n4353) );
  OAI22_X1 U159 ( .A1(n3543), .A2(n4354), .B1(n3351), .B2(n3674), .ZN(n3691)
         );
  NOR2_X1 U160 ( .A1(ADD_RD1[4]), .A2(n3688), .ZN(n3707) );
  NAND2_X1 U161 ( .A1(n3684), .A2(n3700), .ZN(n4355) );
  OAI22_X1 U162 ( .A1(n3095), .A2(n4356), .B1(n3319), .B2(n3675), .ZN(n3690)
         );
  NAND2_X1 U163 ( .A1(n3684), .A2(n3701), .ZN(n4358) );
  OAI22_X1 U164 ( .A1(n3287), .A2(n3676), .B1(n2839), .B2(n4357), .ZN(n3689)
         );
  NOR4_X1 U165 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3720) );
  OAI22_X1 U166 ( .A1(n3063), .A2(n4364), .B1(n3031), .B2(n4363), .ZN(n3697)
         );
  NOR3_X1 U167 ( .A1(ADD_RD1[2]), .A2(n3698), .A3(n3693), .ZN(n3708) );
  NAND2_X1 U168 ( .A1(n3708), .A2(n3699), .ZN(n4366) );
  NAND2_X1 U169 ( .A1(n3673), .A2(n3700), .ZN(n4365) );
  OAI22_X1 U170 ( .A1(n3479), .A2(n3678), .B1(n2807), .B2(n3677), .ZN(n3696)
         );
  NOR3_X1 U171 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[2]), .A3(n3693), .ZN(n3709) );
  NAND2_X1 U172 ( .A1(n3709), .A2(n3699), .ZN(n4367) );
  OAI22_X1 U173 ( .A1(n2775), .A2(n4368), .B1(n3223), .B2(n3679), .ZN(n3695)
         );
  NAND2_X1 U174 ( .A1(n3708), .A2(n3700), .ZN(n4370) );
  NAND2_X1 U175 ( .A1(n3708), .A2(n3701), .ZN(n4369) );
  OAI22_X1 U176 ( .A1(n3447), .A2(n3681), .B1(n3415), .B2(n3680), .ZN(n3694)
         );
  NOR4_X1 U177 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3719) );
  NOR3_X1 U178 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[4]), .A3(n3698), .ZN(n3710) );
  OAI22_X1 U179 ( .A1(n2967), .A2(n4376), .B1(n3191), .B2(n4375), .ZN(n3705)
         );
  NOR3_X1 U180 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[2]), .A3(ADD_RD1[4]), .ZN(n3711)
         );
  OAI22_X1 U181 ( .A1(n3159), .A2(n4378), .B1(n2711), .B2(n4377), .ZN(n3704)
         );
  OAI22_X1 U182 ( .A1(n2935), .A2(n4380), .B1(n2903), .B2(n4379), .ZN(n3703)
         );
  NAND2_X1 U183 ( .A1(n3711), .A2(n3701), .ZN(n4381) );
  OAI22_X1 U184 ( .A1(n2679), .A2(n4382), .B1(n2647), .B2(n3682), .ZN(n3702)
         );
  NOR4_X1 U185 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3718) );
  OAI22_X1 U186 ( .A1(n3511), .A2(n4388), .B1(n3255), .B2(n4387), .ZN(n3715)
         );
  OAI22_X1 U187 ( .A1(n2999), .A2(n4389), .B1(n2743), .B2(n3672), .ZN(n3714)
         );
  OAI22_X1 U188 ( .A1(n3383), .A2(n4391), .B1(n3127), .B2(n4390), .ZN(n3713)
         );
  OAI22_X1 U189 ( .A1(n2871), .A2(n4393), .B1(n2615), .B2(n4392), .ZN(n3712)
         );
  OR4_X1 U190 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716) );
  NAND2_X1 U191 ( .A1(n3685), .A2(n3716), .ZN(n3717) );
  NAND4_X1 U192 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(N379) );
  OAI22_X1 U193 ( .A1(n3606), .A2(n4352), .B1(n3574), .B2(n4351), .ZN(n3724)
         );
  OAI22_X1 U194 ( .A1(n3542), .A2(n4354), .B1(n3350), .B2(n4353), .ZN(n3723)
         );
  OAI22_X1 U195 ( .A1(n3094), .A2(n4356), .B1(n3318), .B2(n4355), .ZN(n3722)
         );
  OAI22_X1 U196 ( .A1(n3286), .A2(n4358), .B1(n2838), .B2(n4357), .ZN(n3721)
         );
  NOR4_X1 U197 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3741) );
  OAI22_X1 U198 ( .A1(n3062), .A2(n4364), .B1(n3030), .B2(n4363), .ZN(n3728)
         );
  OAI22_X1 U199 ( .A1(n3478), .A2(n4366), .B1(n2806), .B2(n4365), .ZN(n3727)
         );
  OAI22_X1 U200 ( .A1(n2774), .A2(n4368), .B1(n3222), .B2(n4367), .ZN(n3726)
         );
  OAI22_X1 U201 ( .A1(n3446), .A2(n4370), .B1(n3414), .B2(n4369), .ZN(n3725)
         );
  NOR4_X1 U202 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3740) );
  OAI22_X1 U203 ( .A1(n2966), .A2(n4376), .B1(n3190), .B2(n4375), .ZN(n3732)
         );
  OAI22_X1 U204 ( .A1(n3158), .A2(n4378), .B1(n2710), .B2(n4377), .ZN(n3731)
         );
  OAI22_X1 U205 ( .A1(n2934), .A2(n4380), .B1(n2902), .B2(n4379), .ZN(n3730)
         );
  OAI22_X1 U206 ( .A1(n2678), .A2(n4382), .B1(n2646), .B2(n4381), .ZN(n3729)
         );
  NOR4_X1 U207 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3739) );
  OAI22_X1 U208 ( .A1(n3510), .A2(n4388), .B1(n3254), .B2(n3683), .ZN(n3736)
         );
  OAI22_X1 U209 ( .A1(n2998), .A2(n4389), .B1(n2742), .B2(n3672), .ZN(n3735)
         );
  OAI22_X1 U210 ( .A1(n3382), .A2(n4391), .B1(n3126), .B2(n4390), .ZN(n3734)
         );
  OAI22_X1 U211 ( .A1(n2870), .A2(n4393), .B1(n2614), .B2(n4392), .ZN(n3733)
         );
  OR4_X1 U212 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3737) );
  NAND2_X1 U213 ( .A1(n4399), .A2(n3737), .ZN(n3738) );
  NAND4_X1 U214 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(N380) );
  OAI22_X1 U215 ( .A1(n3605), .A2(n4352), .B1(n3573), .B2(n4351), .ZN(n3745)
         );
  OAI22_X1 U216 ( .A1(n3541), .A2(n4354), .B1(n3349), .B2(n3674), .ZN(n3744)
         );
  OAI22_X1 U217 ( .A1(n3093), .A2(n4356), .B1(n3317), .B2(n3675), .ZN(n3743)
         );
  OAI22_X1 U218 ( .A1(n3285), .A2(n3676), .B1(n2837), .B2(n4357), .ZN(n3742)
         );
  NOR4_X1 U219 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3762) );
  OAI22_X1 U220 ( .A1(n3061), .A2(n4364), .B1(n3029), .B2(n4363), .ZN(n3749)
         );
  OAI22_X1 U221 ( .A1(n3477), .A2(n3678), .B1(n2805), .B2(n3677), .ZN(n3748)
         );
  OAI22_X1 U222 ( .A1(n2773), .A2(n4368), .B1(n3221), .B2(n3679), .ZN(n3747)
         );
  OAI22_X1 U223 ( .A1(n3445), .A2(n3681), .B1(n3413), .B2(n3680), .ZN(n3746)
         );
  NOR4_X1 U224 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3761) );
  OAI22_X1 U225 ( .A1(n2965), .A2(n4376), .B1(n3189), .B2(n4375), .ZN(n3753)
         );
  OAI22_X1 U226 ( .A1(n3157), .A2(n4378), .B1(n2709), .B2(n4377), .ZN(n3752)
         );
  OAI22_X1 U227 ( .A1(n2933), .A2(n4380), .B1(n2901), .B2(n4379), .ZN(n3751)
         );
  OAI22_X1 U228 ( .A1(n2677), .A2(n4382), .B1(n2645), .B2(n3682), .ZN(n3750)
         );
  NOR4_X1 U229 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3760) );
  OAI22_X1 U230 ( .A1(n3509), .A2(n4388), .B1(n3253), .B2(n4387), .ZN(n3757)
         );
  OAI22_X1 U231 ( .A1(n2997), .A2(n4389), .B1(n2741), .B2(n3672), .ZN(n3756)
         );
  OAI22_X1 U232 ( .A1(n3381), .A2(n4391), .B1(n3125), .B2(n4390), .ZN(n3755)
         );
  OAI22_X1 U233 ( .A1(n2869), .A2(n4393), .B1(n2613), .B2(n4392), .ZN(n3754)
         );
  OR4_X1 U234 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758) );
  NAND2_X1 U235 ( .A1(n3685), .A2(n3758), .ZN(n3759) );
  NAND4_X1 U236 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(N381) );
  OAI22_X1 U237 ( .A1(n3604), .A2(n4352), .B1(n3572), .B2(n4351), .ZN(n3766)
         );
  OAI22_X1 U238 ( .A1(n3540), .A2(n4354), .B1(n3348), .B2(n4353), .ZN(n3765)
         );
  OAI22_X1 U239 ( .A1(n3092), .A2(n4356), .B1(n3316), .B2(n4355), .ZN(n3764)
         );
  OAI22_X1 U240 ( .A1(n3284), .A2(n4358), .B1(n2836), .B2(n4357), .ZN(n3763)
         );
  NOR4_X1 U241 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3783) );
  OAI22_X1 U242 ( .A1(n3060), .A2(n4364), .B1(n3028), .B2(n4363), .ZN(n3770)
         );
  OAI22_X1 U243 ( .A1(n3476), .A2(n4366), .B1(n2804), .B2(n4365), .ZN(n3769)
         );
  OAI22_X1 U244 ( .A1(n2772), .A2(n4368), .B1(n3220), .B2(n4367), .ZN(n3768)
         );
  OAI22_X1 U245 ( .A1(n3444), .A2(n4370), .B1(n3412), .B2(n4369), .ZN(n3767)
         );
  NOR4_X1 U246 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3782) );
  OAI22_X1 U247 ( .A1(n2964), .A2(n4376), .B1(n3188), .B2(n4375), .ZN(n3774)
         );
  OAI22_X1 U248 ( .A1(n3156), .A2(n4378), .B1(n2708), .B2(n4377), .ZN(n3773)
         );
  OAI22_X1 U249 ( .A1(n2932), .A2(n4380), .B1(n2900), .B2(n4379), .ZN(n3772)
         );
  OAI22_X1 U250 ( .A1(n2676), .A2(n4382), .B1(n2644), .B2(n4381), .ZN(n3771)
         );
  NOR4_X1 U251 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3781) );
  OAI22_X1 U252 ( .A1(n3508), .A2(n4388), .B1(n3252), .B2(n3683), .ZN(n3778)
         );
  OAI22_X1 U253 ( .A1(n2996), .A2(n4389), .B1(n2740), .B2(n3672), .ZN(n3777)
         );
  OAI22_X1 U254 ( .A1(n3380), .A2(n4391), .B1(n3124), .B2(n4390), .ZN(n3776)
         );
  OAI22_X1 U255 ( .A1(n2868), .A2(n4393), .B1(n2612), .B2(n4392), .ZN(n3775)
         );
  OR4_X1 U256 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779) );
  NAND2_X1 U257 ( .A1(n4399), .A2(n3779), .ZN(n3780) );
  NAND4_X1 U258 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(N382) );
  OAI22_X1 U259 ( .A1(n3603), .A2(n4352), .B1(n3571), .B2(n4351), .ZN(n3787)
         );
  OAI22_X1 U260 ( .A1(n3539), .A2(n4354), .B1(n3347), .B2(n3674), .ZN(n3786)
         );
  OAI22_X1 U261 ( .A1(n3091), .A2(n4356), .B1(n3315), .B2(n3675), .ZN(n3785)
         );
  OAI22_X1 U262 ( .A1(n3283), .A2(n3676), .B1(n2835), .B2(n4357), .ZN(n3784)
         );
  NOR4_X1 U263 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3804) );
  OAI22_X1 U264 ( .A1(n3059), .A2(n4364), .B1(n3027), .B2(n4363), .ZN(n3791)
         );
  OAI22_X1 U265 ( .A1(n3475), .A2(n3678), .B1(n2803), .B2(n3677), .ZN(n3790)
         );
  OAI22_X1 U266 ( .A1(n2771), .A2(n4368), .B1(n3219), .B2(n3679), .ZN(n3789)
         );
  OAI22_X1 U267 ( .A1(n3443), .A2(n3681), .B1(n3411), .B2(n3680), .ZN(n3788)
         );
  NOR4_X1 U268 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3803) );
  OAI22_X1 U269 ( .A1(n2963), .A2(n4376), .B1(n3187), .B2(n4375), .ZN(n3795)
         );
  OAI22_X1 U270 ( .A1(n3155), .A2(n4378), .B1(n2707), .B2(n4377), .ZN(n3794)
         );
  OAI22_X1 U271 ( .A1(n2931), .A2(n4380), .B1(n2899), .B2(n4379), .ZN(n3793)
         );
  OAI22_X1 U272 ( .A1(n2675), .A2(n4382), .B1(n2643), .B2(n3682), .ZN(n3792)
         );
  NOR4_X1 U273 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3802) );
  OAI22_X1 U274 ( .A1(n3507), .A2(n4388), .B1(n3251), .B2(n4387), .ZN(n3799)
         );
  OAI22_X1 U275 ( .A1(n2995), .A2(n4389), .B1(n2739), .B2(n3672), .ZN(n3798)
         );
  OAI22_X1 U276 ( .A1(n3379), .A2(n4391), .B1(n3123), .B2(n4390), .ZN(n3797)
         );
  OAI22_X1 U277 ( .A1(n2867), .A2(n4393), .B1(n2611), .B2(n4392), .ZN(n3796)
         );
  OR4_X1 U278 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800) );
  NAND2_X1 U279 ( .A1(n3685), .A2(n3800), .ZN(n3801) );
  NAND4_X1 U280 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(N383) );
  OAI22_X1 U281 ( .A1(n3602), .A2(n4352), .B1(n3570), .B2(n4351), .ZN(n3808)
         );
  OAI22_X1 U282 ( .A1(n3538), .A2(n4354), .B1(n3346), .B2(n4353), .ZN(n3807)
         );
  OAI22_X1 U283 ( .A1(n3090), .A2(n4356), .B1(n3314), .B2(n4355), .ZN(n3806)
         );
  OAI22_X1 U284 ( .A1(n3282), .A2(n4358), .B1(n2834), .B2(n4357), .ZN(n3805)
         );
  NOR4_X1 U285 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3825) );
  OAI22_X1 U286 ( .A1(n3058), .A2(n4364), .B1(n3026), .B2(n4363), .ZN(n3812)
         );
  OAI22_X1 U287 ( .A1(n3474), .A2(n4366), .B1(n2802), .B2(n4365), .ZN(n3811)
         );
  OAI22_X1 U288 ( .A1(n2770), .A2(n4368), .B1(n3218), .B2(n4367), .ZN(n3810)
         );
  OAI22_X1 U289 ( .A1(n3442), .A2(n4370), .B1(n3410), .B2(n4369), .ZN(n3809)
         );
  NOR4_X1 U290 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3824) );
  OAI22_X1 U291 ( .A1(n2962), .A2(n4376), .B1(n3186), .B2(n4375), .ZN(n3816)
         );
  OAI22_X1 U292 ( .A1(n3154), .A2(n4378), .B1(n2706), .B2(n4377), .ZN(n3815)
         );
  OAI22_X1 U293 ( .A1(n2930), .A2(n4380), .B1(n2898), .B2(n4379), .ZN(n3814)
         );
  OAI22_X1 U294 ( .A1(n2674), .A2(n4382), .B1(n2642), .B2(n4381), .ZN(n3813)
         );
  NOR4_X1 U295 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3823) );
  OAI22_X1 U296 ( .A1(n3506), .A2(n4388), .B1(n3250), .B2(n3683), .ZN(n3820)
         );
  OAI22_X1 U297 ( .A1(n2994), .A2(n4389), .B1(n2738), .B2(n3672), .ZN(n3819)
         );
  OAI22_X1 U298 ( .A1(n3378), .A2(n4391), .B1(n3122), .B2(n4390), .ZN(n3818)
         );
  OAI22_X1 U299 ( .A1(n2866), .A2(n4393), .B1(n2610), .B2(n4392), .ZN(n3817)
         );
  OR4_X1 U300 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821) );
  NAND2_X1 U301 ( .A1(n4399), .A2(n3821), .ZN(n3822) );
  NAND4_X1 U302 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(N384) );
  OAI22_X1 U303 ( .A1(n3601), .A2(n4352), .B1(n3569), .B2(n4351), .ZN(n3829)
         );
  OAI22_X1 U304 ( .A1(n3537), .A2(n4354), .B1(n3345), .B2(n4353), .ZN(n3828)
         );
  OAI22_X1 U305 ( .A1(n3089), .A2(n4356), .B1(n3313), .B2(n4355), .ZN(n3827)
         );
  OAI22_X1 U306 ( .A1(n3281), .A2(n4358), .B1(n2833), .B2(n4357), .ZN(n3826)
         );
  NOR4_X1 U307 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3846) );
  OAI22_X1 U308 ( .A1(n3057), .A2(n4364), .B1(n3025), .B2(n4363), .ZN(n3833)
         );
  OAI22_X1 U309 ( .A1(n3473), .A2(n4366), .B1(n2801), .B2(n4365), .ZN(n3832)
         );
  OAI22_X1 U310 ( .A1(n2769), .A2(n4368), .B1(n3217), .B2(n4367), .ZN(n3831)
         );
  OAI22_X1 U311 ( .A1(n3441), .A2(n4370), .B1(n3409), .B2(n4369), .ZN(n3830)
         );
  NOR4_X1 U312 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3845) );
  OAI22_X1 U313 ( .A1(n2961), .A2(n4376), .B1(n3185), .B2(n4375), .ZN(n3837)
         );
  OAI22_X1 U314 ( .A1(n3153), .A2(n4378), .B1(n2705), .B2(n4377), .ZN(n3836)
         );
  OAI22_X1 U315 ( .A1(n2929), .A2(n4380), .B1(n2897), .B2(n4379), .ZN(n3835)
         );
  OAI22_X1 U316 ( .A1(n2673), .A2(n4382), .B1(n2641), .B2(n4381), .ZN(n3834)
         );
  NOR4_X1 U317 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3844) );
  OAI22_X1 U318 ( .A1(n3505), .A2(n4388), .B1(n3249), .B2(n4387), .ZN(n3841)
         );
  OAI22_X1 U319 ( .A1(n2993), .A2(n4389), .B1(n2737), .B2(n3672), .ZN(n3840)
         );
  OAI22_X1 U320 ( .A1(n3377), .A2(n4391), .B1(n3121), .B2(n4390), .ZN(n3839)
         );
  OAI22_X1 U321 ( .A1(n2865), .A2(n4393), .B1(n2609), .B2(n4392), .ZN(n3838)
         );
  OR4_X1 U322 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842) );
  NAND2_X1 U323 ( .A1(n4399), .A2(n3842), .ZN(n3843) );
  NAND4_X1 U324 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(N385) );
  OAI22_X1 U325 ( .A1(n3600), .A2(n4352), .B1(n3568), .B2(n4351), .ZN(n3850)
         );
  OAI22_X1 U326 ( .A1(n3536), .A2(n4354), .B1(n3344), .B2(n4353), .ZN(n3849)
         );
  OAI22_X1 U327 ( .A1(n3088), .A2(n4356), .B1(n3312), .B2(n4355), .ZN(n3848)
         );
  OAI22_X1 U328 ( .A1(n3280), .A2(n4358), .B1(n2832), .B2(n4357), .ZN(n3847)
         );
  NOR4_X1 U329 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3867) );
  OAI22_X1 U330 ( .A1(n3056), .A2(n4364), .B1(n3024), .B2(n4363), .ZN(n3854)
         );
  OAI22_X1 U331 ( .A1(n3472), .A2(n4366), .B1(n2800), .B2(n4365), .ZN(n3853)
         );
  OAI22_X1 U332 ( .A1(n2768), .A2(n4368), .B1(n3216), .B2(n4367), .ZN(n3852)
         );
  OAI22_X1 U333 ( .A1(n3440), .A2(n4370), .B1(n3408), .B2(n4369), .ZN(n3851)
         );
  NOR4_X1 U334 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3866) );
  OAI22_X1 U335 ( .A1(n2960), .A2(n4376), .B1(n3184), .B2(n4375), .ZN(n3858)
         );
  OAI22_X1 U336 ( .A1(n3152), .A2(n4378), .B1(n2704), .B2(n4377), .ZN(n3857)
         );
  OAI22_X1 U337 ( .A1(n2928), .A2(n4380), .B1(n2896), .B2(n4379), .ZN(n3856)
         );
  OAI22_X1 U338 ( .A1(n2672), .A2(n4382), .B1(n2640), .B2(n4381), .ZN(n3855)
         );
  NOR4_X1 U339 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3865) );
  OAI22_X1 U340 ( .A1(n3504), .A2(n4388), .B1(n3248), .B2(n3683), .ZN(n3862)
         );
  OAI22_X1 U341 ( .A1(n2992), .A2(n4389), .B1(n2736), .B2(n3672), .ZN(n3861)
         );
  OAI22_X1 U342 ( .A1(n3376), .A2(n4391), .B1(n3120), .B2(n4390), .ZN(n3860)
         );
  OAI22_X1 U343 ( .A1(n2864), .A2(n4393), .B1(n2608), .B2(n4392), .ZN(n3859)
         );
  OR4_X1 U344 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863) );
  NAND2_X1 U345 ( .A1(n4399), .A2(n3863), .ZN(n3864) );
  NAND4_X1 U346 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(N386) );
  OAI22_X1 U347 ( .A1(n3599), .A2(n4352), .B1(n3567), .B2(n4351), .ZN(n3871)
         );
  OAI22_X1 U348 ( .A1(n3535), .A2(n4354), .B1(n3343), .B2(n4353), .ZN(n3870)
         );
  OAI22_X1 U349 ( .A1(n3087), .A2(n4356), .B1(n3311), .B2(n4355), .ZN(n3869)
         );
  OAI22_X1 U350 ( .A1(n3279), .A2(n4358), .B1(n2831), .B2(n4357), .ZN(n3868)
         );
  NOR4_X1 U351 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3888) );
  OAI22_X1 U352 ( .A1(n3055), .A2(n4364), .B1(n3023), .B2(n4363), .ZN(n3875)
         );
  OAI22_X1 U353 ( .A1(n3471), .A2(n4366), .B1(n2799), .B2(n4365), .ZN(n3874)
         );
  OAI22_X1 U354 ( .A1(n2767), .A2(n4368), .B1(n3215), .B2(n4367), .ZN(n3873)
         );
  OAI22_X1 U355 ( .A1(n3439), .A2(n4370), .B1(n3407), .B2(n4369), .ZN(n3872)
         );
  NOR4_X1 U356 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3887) );
  OAI22_X1 U357 ( .A1(n2959), .A2(n4376), .B1(n3183), .B2(n4375), .ZN(n3879)
         );
  OAI22_X1 U358 ( .A1(n3151), .A2(n4378), .B1(n2703), .B2(n4377), .ZN(n3878)
         );
  OAI22_X1 U359 ( .A1(n2927), .A2(n4380), .B1(n2895), .B2(n4379), .ZN(n3877)
         );
  OAI22_X1 U360 ( .A1(n2671), .A2(n4382), .B1(n2639), .B2(n4381), .ZN(n3876)
         );
  NOR4_X1 U361 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3886) );
  OAI22_X1 U362 ( .A1(n3503), .A2(n4388), .B1(n3247), .B2(n4387), .ZN(n3883)
         );
  OAI22_X1 U363 ( .A1(n2991), .A2(n4389), .B1(n2735), .B2(n3672), .ZN(n3882)
         );
  OAI22_X1 U364 ( .A1(n3375), .A2(n4391), .B1(n3119), .B2(n4390), .ZN(n3881)
         );
  OAI22_X1 U365 ( .A1(n2863), .A2(n4393), .B1(n2607), .B2(n4392), .ZN(n3880)
         );
  OR4_X1 U366 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884) );
  NAND2_X1 U367 ( .A1(n4399), .A2(n3884), .ZN(n3885) );
  NAND4_X1 U368 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(N387) );
  OAI22_X1 U369 ( .A1(n3598), .A2(n4352), .B1(n3566), .B2(n4351), .ZN(n3892)
         );
  OAI22_X1 U370 ( .A1(n3534), .A2(n4354), .B1(n3342), .B2(n4353), .ZN(n3891)
         );
  OAI22_X1 U371 ( .A1(n3086), .A2(n4356), .B1(n3310), .B2(n4355), .ZN(n3890)
         );
  OAI22_X1 U372 ( .A1(n3278), .A2(n4358), .B1(n2830), .B2(n4357), .ZN(n3889)
         );
  NOR4_X1 U373 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3909) );
  OAI22_X1 U374 ( .A1(n3054), .A2(n4364), .B1(n3022), .B2(n4363), .ZN(n3896)
         );
  OAI22_X1 U375 ( .A1(n3470), .A2(n4366), .B1(n2798), .B2(n4365), .ZN(n3895)
         );
  OAI22_X1 U376 ( .A1(n2766), .A2(n4368), .B1(n3214), .B2(n4367), .ZN(n3894)
         );
  OAI22_X1 U377 ( .A1(n3438), .A2(n4370), .B1(n3406), .B2(n4369), .ZN(n3893)
         );
  NOR4_X1 U378 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3908) );
  OAI22_X1 U379 ( .A1(n2958), .A2(n4376), .B1(n3182), .B2(n4375), .ZN(n3900)
         );
  OAI22_X1 U380 ( .A1(n3150), .A2(n4378), .B1(n2702), .B2(n4377), .ZN(n3899)
         );
  OAI22_X1 U381 ( .A1(n2926), .A2(n4380), .B1(n2894), .B2(n4379), .ZN(n3898)
         );
  OAI22_X1 U382 ( .A1(n2670), .A2(n4382), .B1(n2638), .B2(n4381), .ZN(n3897)
         );
  NOR4_X1 U383 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3907) );
  OAI22_X1 U384 ( .A1(n3502), .A2(n4388), .B1(n3246), .B2(n3683), .ZN(n3904)
         );
  OAI22_X1 U385 ( .A1(n2990), .A2(n4389), .B1(n2734), .B2(n3672), .ZN(n3903)
         );
  OAI22_X1 U386 ( .A1(n3374), .A2(n4391), .B1(n3118), .B2(n4390), .ZN(n3902)
         );
  OAI22_X1 U387 ( .A1(n2862), .A2(n4393), .B1(n2606), .B2(n4392), .ZN(n3901)
         );
  OR4_X1 U388 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905) );
  NAND2_X1 U389 ( .A1(n4399), .A2(n3905), .ZN(n3906) );
  NAND4_X1 U390 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(N388) );
  OAI22_X1 U391 ( .A1(n3597), .A2(n4352), .B1(n3565), .B2(n4351), .ZN(n3913)
         );
  OAI22_X1 U392 ( .A1(n3533), .A2(n4354), .B1(n3341), .B2(n4353), .ZN(n3912)
         );
  OAI22_X1 U393 ( .A1(n3085), .A2(n4356), .B1(n3309), .B2(n4355), .ZN(n3911)
         );
  OAI22_X1 U394 ( .A1(n3277), .A2(n4358), .B1(n2829), .B2(n4357), .ZN(n3910)
         );
  NOR4_X1 U395 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3930) );
  OAI22_X1 U396 ( .A1(n3053), .A2(n4364), .B1(n3021), .B2(n4363), .ZN(n3917)
         );
  OAI22_X1 U397 ( .A1(n3469), .A2(n4366), .B1(n2797), .B2(n4365), .ZN(n3916)
         );
  OAI22_X1 U398 ( .A1(n2765), .A2(n4368), .B1(n3213), .B2(n4367), .ZN(n3915)
         );
  OAI22_X1 U399 ( .A1(n3437), .A2(n4370), .B1(n3405), .B2(n4369), .ZN(n3914)
         );
  NOR4_X1 U400 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3929) );
  OAI22_X1 U401 ( .A1(n2957), .A2(n4376), .B1(n3181), .B2(n4375), .ZN(n3921)
         );
  OAI22_X1 U402 ( .A1(n3149), .A2(n4378), .B1(n2701), .B2(n4377), .ZN(n3920)
         );
  OAI22_X1 U403 ( .A1(n2925), .A2(n4380), .B1(n2893), .B2(n4379), .ZN(n3919)
         );
  OAI22_X1 U404 ( .A1(n2669), .A2(n4382), .B1(n2637), .B2(n4381), .ZN(n3918)
         );
  NOR4_X1 U405 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3928) );
  OAI22_X1 U406 ( .A1(n3501), .A2(n4388), .B1(n3245), .B2(n4387), .ZN(n3925)
         );
  OAI22_X1 U407 ( .A1(n2989), .A2(n4389), .B1(n2733), .B2(n3672), .ZN(n3924)
         );
  OAI22_X1 U408 ( .A1(n3373), .A2(n4391), .B1(n3117), .B2(n4390), .ZN(n3923)
         );
  OAI22_X1 U409 ( .A1(n2861), .A2(n4393), .B1(n2605), .B2(n4392), .ZN(n3922)
         );
  OR4_X1 U410 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3926) );
  NAND2_X1 U411 ( .A1(n4399), .A2(n3926), .ZN(n3927) );
  NAND4_X1 U412 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(N389) );
  OAI22_X1 U413 ( .A1(n3596), .A2(n4352), .B1(n3564), .B2(n4351), .ZN(n3934)
         );
  OAI22_X1 U414 ( .A1(n3532), .A2(n4354), .B1(n3340), .B2(n4353), .ZN(n3933)
         );
  OAI22_X1 U415 ( .A1(n3084), .A2(n4356), .B1(n3308), .B2(n4355), .ZN(n3932)
         );
  OAI22_X1 U416 ( .A1(n3276), .A2(n4358), .B1(n2828), .B2(n4357), .ZN(n3931)
         );
  NOR4_X1 U417 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3951) );
  OAI22_X1 U418 ( .A1(n3052), .A2(n4364), .B1(n3020), .B2(n4363), .ZN(n3938)
         );
  OAI22_X1 U419 ( .A1(n3468), .A2(n4366), .B1(n2796), .B2(n4365), .ZN(n3937)
         );
  OAI22_X1 U420 ( .A1(n2764), .A2(n4368), .B1(n3212), .B2(n4367), .ZN(n3936)
         );
  OAI22_X1 U421 ( .A1(n3436), .A2(n4370), .B1(n3404), .B2(n4369), .ZN(n3935)
         );
  NOR4_X1 U422 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3950) );
  OAI22_X1 U423 ( .A1(n2956), .A2(n4376), .B1(n3180), .B2(n4375), .ZN(n3942)
         );
  OAI22_X1 U424 ( .A1(n3148), .A2(n4378), .B1(n2700), .B2(n4377), .ZN(n3941)
         );
  OAI22_X1 U425 ( .A1(n2924), .A2(n4380), .B1(n2892), .B2(n4379), .ZN(n3940)
         );
  OAI22_X1 U426 ( .A1(n2668), .A2(n4382), .B1(n2636), .B2(n4381), .ZN(n3939)
         );
  NOR4_X1 U427 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3949) );
  OAI22_X1 U428 ( .A1(n3500), .A2(n4388), .B1(n3244), .B2(n4387), .ZN(n3946)
         );
  OAI22_X1 U429 ( .A1(n2988), .A2(n4389), .B1(n2732), .B2(n3672), .ZN(n3945)
         );
  OAI22_X1 U430 ( .A1(n3372), .A2(n4391), .B1(n3116), .B2(n4390), .ZN(n3944)
         );
  OAI22_X1 U431 ( .A1(n2860), .A2(n4393), .B1(n2604), .B2(n4392), .ZN(n3943)
         );
  OR4_X1 U432 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947) );
  NAND2_X1 U433 ( .A1(n4399), .A2(n3947), .ZN(n3948) );
  NAND4_X1 U434 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(N390) );
  OAI22_X1 U435 ( .A1(n3595), .A2(n4352), .B1(n3563), .B2(n4351), .ZN(n3955)
         );
  OAI22_X1 U436 ( .A1(n3531), .A2(n4354), .B1(n3339), .B2(n4353), .ZN(n3954)
         );
  OAI22_X1 U437 ( .A1(n3083), .A2(n4356), .B1(n3307), .B2(n4355), .ZN(n3953)
         );
  OAI22_X1 U438 ( .A1(n3275), .A2(n4358), .B1(n2827), .B2(n4357), .ZN(n3952)
         );
  NOR4_X1 U439 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3972) );
  OAI22_X1 U440 ( .A1(n3051), .A2(n4364), .B1(n3019), .B2(n4363), .ZN(n3959)
         );
  OAI22_X1 U441 ( .A1(n3467), .A2(n4366), .B1(n2795), .B2(n4365), .ZN(n3958)
         );
  OAI22_X1 U442 ( .A1(n2763), .A2(n4368), .B1(n3211), .B2(n4367), .ZN(n3957)
         );
  OAI22_X1 U443 ( .A1(n3435), .A2(n4370), .B1(n3403), .B2(n4369), .ZN(n3956)
         );
  NOR4_X1 U444 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3971) );
  OAI22_X1 U445 ( .A1(n2955), .A2(n4376), .B1(n3179), .B2(n4375), .ZN(n3963)
         );
  OAI22_X1 U446 ( .A1(n3147), .A2(n4378), .B1(n2699), .B2(n4377), .ZN(n3962)
         );
  OAI22_X1 U447 ( .A1(n2923), .A2(n4380), .B1(n2891), .B2(n4379), .ZN(n3961)
         );
  OAI22_X1 U448 ( .A1(n2667), .A2(n4382), .B1(n2635), .B2(n4381), .ZN(n3960)
         );
  NOR4_X1 U449 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3970) );
  OAI22_X1 U450 ( .A1(n3499), .A2(n4388), .B1(n3243), .B2(n3683), .ZN(n3967)
         );
  OAI22_X1 U451 ( .A1(n2987), .A2(n4389), .B1(n2731), .B2(n3672), .ZN(n3966)
         );
  OAI22_X1 U452 ( .A1(n3371), .A2(n4391), .B1(n3115), .B2(n4390), .ZN(n3965)
         );
  OAI22_X1 U453 ( .A1(n2859), .A2(n4393), .B1(n2603), .B2(n4392), .ZN(n3964)
         );
  OR4_X1 U454 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3968) );
  NAND2_X1 U455 ( .A1(n3685), .A2(n3968), .ZN(n3969) );
  NAND4_X1 U456 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(N391) );
  OAI22_X1 U457 ( .A1(n3594), .A2(n4352), .B1(n3562), .B2(n4351), .ZN(n3976)
         );
  OAI22_X1 U458 ( .A1(n3530), .A2(n4354), .B1(n3338), .B2(n3674), .ZN(n3975)
         );
  OAI22_X1 U459 ( .A1(n3082), .A2(n4356), .B1(n3306), .B2(n3675), .ZN(n3974)
         );
  OAI22_X1 U460 ( .A1(n3274), .A2(n3676), .B1(n2826), .B2(n4357), .ZN(n3973)
         );
  NOR4_X1 U461 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3993) );
  OAI22_X1 U462 ( .A1(n3050), .A2(n4364), .B1(n3018), .B2(n4363), .ZN(n3980)
         );
  OAI22_X1 U463 ( .A1(n3466), .A2(n3678), .B1(n2794), .B2(n3677), .ZN(n3979)
         );
  OAI22_X1 U464 ( .A1(n2762), .A2(n4368), .B1(n3210), .B2(n3679), .ZN(n3978)
         );
  OAI22_X1 U465 ( .A1(n3434), .A2(n3681), .B1(n3402), .B2(n3680), .ZN(n3977)
         );
  NOR4_X1 U466 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3992) );
  OAI22_X1 U467 ( .A1(n2954), .A2(n4376), .B1(n3178), .B2(n4375), .ZN(n3984)
         );
  OAI22_X1 U468 ( .A1(n3146), .A2(n4378), .B1(n2698), .B2(n4377), .ZN(n3983)
         );
  OAI22_X1 U469 ( .A1(n2922), .A2(n4380), .B1(n2890), .B2(n4379), .ZN(n3982)
         );
  OAI22_X1 U470 ( .A1(n2666), .A2(n4382), .B1(n2634), .B2(n3682), .ZN(n3981)
         );
  NOR4_X1 U471 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3991) );
  OAI22_X1 U472 ( .A1(n3498), .A2(n4388), .B1(n3242), .B2(n3683), .ZN(n3988)
         );
  OAI22_X1 U473 ( .A1(n2986), .A2(n4389), .B1(n2730), .B2(n3672), .ZN(n3987)
         );
  OAI22_X1 U474 ( .A1(n3370), .A2(n4391), .B1(n3114), .B2(n4390), .ZN(n3986)
         );
  OAI22_X1 U475 ( .A1(n2858), .A2(n4393), .B1(n2602), .B2(n4392), .ZN(n3985)
         );
  OR4_X1 U476 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989) );
  NAND2_X1 U477 ( .A1(n3685), .A2(n3989), .ZN(n3990) );
  NAND4_X1 U478 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(N392) );
  OAI22_X1 U479 ( .A1(n3593), .A2(n4352), .B1(n3561), .B2(n4351), .ZN(n3997)
         );
  OAI22_X1 U480 ( .A1(n3529), .A2(n4354), .B1(n3337), .B2(n4353), .ZN(n3996)
         );
  OAI22_X1 U481 ( .A1(n3081), .A2(n4356), .B1(n3305), .B2(n4355), .ZN(n3995)
         );
  OAI22_X1 U482 ( .A1(n3273), .A2(n4358), .B1(n2825), .B2(n4357), .ZN(n3994)
         );
  NOR4_X1 U483 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4014) );
  OAI22_X1 U484 ( .A1(n3049), .A2(n4364), .B1(n3017), .B2(n4363), .ZN(n4001)
         );
  OAI22_X1 U485 ( .A1(n3465), .A2(n4366), .B1(n2793), .B2(n4365), .ZN(n4000)
         );
  OAI22_X1 U486 ( .A1(n2761), .A2(n4368), .B1(n3209), .B2(n4367), .ZN(n3999)
         );
  OAI22_X1 U487 ( .A1(n3433), .A2(n4370), .B1(n3401), .B2(n4369), .ZN(n3998)
         );
  NOR4_X1 U488 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4013) );
  OAI22_X1 U489 ( .A1(n2953), .A2(n4376), .B1(n3177), .B2(n4375), .ZN(n4005)
         );
  OAI22_X1 U490 ( .A1(n3145), .A2(n4378), .B1(n2697), .B2(n4377), .ZN(n4004)
         );
  OAI22_X1 U491 ( .A1(n2921), .A2(n4380), .B1(n2889), .B2(n4379), .ZN(n4003)
         );
  OAI22_X1 U492 ( .A1(n2665), .A2(n4382), .B1(n2633), .B2(n4381), .ZN(n4002)
         );
  NOR4_X1 U493 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4012) );
  OAI22_X1 U494 ( .A1(n3497), .A2(n4388), .B1(n3241), .B2(n3683), .ZN(n4009)
         );
  OAI22_X1 U495 ( .A1(n2985), .A2(n4389), .B1(n2729), .B2(n3672), .ZN(n4008)
         );
  OAI22_X1 U496 ( .A1(n3369), .A2(n4391), .B1(n3113), .B2(n4390), .ZN(n4007)
         );
  OAI22_X1 U497 ( .A1(n2857), .A2(n4393), .B1(n2601), .B2(n4392), .ZN(n4006)
         );
  OR4_X1 U498 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010) );
  NAND2_X1 U499 ( .A1(n3685), .A2(n4010), .ZN(n4011) );
  NAND4_X1 U500 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(N393) );
  OAI22_X1 U501 ( .A1(n3592), .A2(n4352), .B1(n3560), .B2(n4351), .ZN(n4018)
         );
  OAI22_X1 U502 ( .A1(n3528), .A2(n4354), .B1(n3336), .B2(n3674), .ZN(n4017)
         );
  OAI22_X1 U503 ( .A1(n3080), .A2(n4356), .B1(n3304), .B2(n3675), .ZN(n4016)
         );
  OAI22_X1 U504 ( .A1(n3272), .A2(n3676), .B1(n2824), .B2(n4357), .ZN(n4015)
         );
  NOR4_X1 U505 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4035) );
  OAI22_X1 U506 ( .A1(n3048), .A2(n4364), .B1(n3016), .B2(n4363), .ZN(n4022)
         );
  OAI22_X1 U507 ( .A1(n3464), .A2(n3678), .B1(n2792), .B2(n3677), .ZN(n4021)
         );
  OAI22_X1 U508 ( .A1(n2760), .A2(n4368), .B1(n3208), .B2(n3679), .ZN(n4020)
         );
  OAI22_X1 U509 ( .A1(n3432), .A2(n3681), .B1(n3400), .B2(n3680), .ZN(n4019)
         );
  NOR4_X1 U510 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4034) );
  OAI22_X1 U511 ( .A1(n2952), .A2(n4376), .B1(n3176), .B2(n4375), .ZN(n4026)
         );
  OAI22_X1 U512 ( .A1(n3144), .A2(n4378), .B1(n2696), .B2(n4377), .ZN(n4025)
         );
  OAI22_X1 U513 ( .A1(n2920), .A2(n4380), .B1(n2888), .B2(n4379), .ZN(n4024)
         );
  OAI22_X1 U514 ( .A1(n2664), .A2(n4382), .B1(n2632), .B2(n3682), .ZN(n4023)
         );
  NOR4_X1 U515 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4033) );
  OAI22_X1 U516 ( .A1(n3496), .A2(n4388), .B1(n3240), .B2(n3683), .ZN(n4030)
         );
  OAI22_X1 U517 ( .A1(n2984), .A2(n4389), .B1(n2728), .B2(n3672), .ZN(n4029)
         );
  OAI22_X1 U518 ( .A1(n3368), .A2(n4391), .B1(n3112), .B2(n4390), .ZN(n4028)
         );
  OAI22_X1 U519 ( .A1(n2856), .A2(n4393), .B1(n2600), .B2(n4392), .ZN(n4027)
         );
  OR4_X1 U520 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4031) );
  NAND2_X1 U521 ( .A1(n3685), .A2(n4031), .ZN(n4032) );
  NAND4_X1 U522 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(N394) );
  OAI22_X1 U523 ( .A1(n3591), .A2(n4352), .B1(n3559), .B2(n4351), .ZN(n4039)
         );
  OAI22_X1 U524 ( .A1(n3527), .A2(n4354), .B1(n3335), .B2(n4353), .ZN(n4038)
         );
  OAI22_X1 U525 ( .A1(n3079), .A2(n4356), .B1(n3303), .B2(n4355), .ZN(n4037)
         );
  OAI22_X1 U526 ( .A1(n3271), .A2(n4358), .B1(n2823), .B2(n4357), .ZN(n4036)
         );
  NOR4_X1 U527 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4056) );
  OAI22_X1 U528 ( .A1(n3047), .A2(n4364), .B1(n3015), .B2(n4363), .ZN(n4043)
         );
  OAI22_X1 U529 ( .A1(n3463), .A2(n4366), .B1(n2791), .B2(n4365), .ZN(n4042)
         );
  OAI22_X1 U530 ( .A1(n2759), .A2(n4368), .B1(n3207), .B2(n4367), .ZN(n4041)
         );
  OAI22_X1 U531 ( .A1(n3431), .A2(n4370), .B1(n3399), .B2(n4369), .ZN(n4040)
         );
  NOR4_X1 U532 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4055) );
  OAI22_X1 U533 ( .A1(n2951), .A2(n4376), .B1(n3175), .B2(n4375), .ZN(n4047)
         );
  OAI22_X1 U534 ( .A1(n3143), .A2(n4378), .B1(n2695), .B2(n4377), .ZN(n4046)
         );
  OAI22_X1 U535 ( .A1(n2919), .A2(n4380), .B1(n2887), .B2(n4379), .ZN(n4045)
         );
  OAI22_X1 U536 ( .A1(n2663), .A2(n4382), .B1(n2631), .B2(n4381), .ZN(n4044)
         );
  NOR4_X1 U537 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4054) );
  OAI22_X1 U538 ( .A1(n3495), .A2(n4388), .B1(n3239), .B2(n3683), .ZN(n4051)
         );
  OAI22_X1 U539 ( .A1(n2983), .A2(n4389), .B1(n2727), .B2(n3672), .ZN(n4050)
         );
  OAI22_X1 U540 ( .A1(n3367), .A2(n4391), .B1(n3111), .B2(n4390), .ZN(n4049)
         );
  OAI22_X1 U541 ( .A1(n2855), .A2(n4393), .B1(n2599), .B2(n4392), .ZN(n4048)
         );
  OR4_X1 U542 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4052) );
  NAND2_X1 U543 ( .A1(n3685), .A2(n4052), .ZN(n4053) );
  NAND4_X1 U544 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(N395) );
  OAI22_X1 U545 ( .A1(n3590), .A2(n4352), .B1(n3558), .B2(n4351), .ZN(n4060)
         );
  OAI22_X1 U546 ( .A1(n3526), .A2(n4354), .B1(n3334), .B2(n3674), .ZN(n4059)
         );
  OAI22_X1 U547 ( .A1(n3078), .A2(n4356), .B1(n3302), .B2(n3675), .ZN(n4058)
         );
  OAI22_X1 U548 ( .A1(n3270), .A2(n3676), .B1(n2822), .B2(n4357), .ZN(n4057)
         );
  NOR4_X1 U549 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4077) );
  OAI22_X1 U550 ( .A1(n3046), .A2(n4364), .B1(n3014), .B2(n4363), .ZN(n4064)
         );
  OAI22_X1 U551 ( .A1(n3462), .A2(n3678), .B1(n2790), .B2(n3677), .ZN(n4063)
         );
  OAI22_X1 U552 ( .A1(n2758), .A2(n4368), .B1(n3206), .B2(n3679), .ZN(n4062)
         );
  OAI22_X1 U553 ( .A1(n3430), .A2(n3681), .B1(n3398), .B2(n3680), .ZN(n4061)
         );
  NOR4_X1 U554 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4076) );
  OAI22_X1 U555 ( .A1(n2950), .A2(n4376), .B1(n3174), .B2(n4375), .ZN(n4068)
         );
  OAI22_X1 U556 ( .A1(n3142), .A2(n4378), .B1(n2694), .B2(n4377), .ZN(n4067)
         );
  OAI22_X1 U557 ( .A1(n2918), .A2(n4380), .B1(n2886), .B2(n4379), .ZN(n4066)
         );
  OAI22_X1 U558 ( .A1(n2662), .A2(n4382), .B1(n2630), .B2(n3682), .ZN(n4065)
         );
  NOR4_X1 U559 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4075) );
  OAI22_X1 U560 ( .A1(n3494), .A2(n4388), .B1(n3238), .B2(n3683), .ZN(n4072)
         );
  OAI22_X1 U561 ( .A1(n2982), .A2(n4389), .B1(n2726), .B2(n3672), .ZN(n4071)
         );
  OAI22_X1 U562 ( .A1(n3366), .A2(n4391), .B1(n3110), .B2(n4390), .ZN(n4070)
         );
  OAI22_X1 U563 ( .A1(n2854), .A2(n4393), .B1(n2598), .B2(n4392), .ZN(n4069)
         );
  OR4_X1 U564 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4073) );
  NAND2_X1 U565 ( .A1(n3685), .A2(n4073), .ZN(n4074) );
  NAND4_X1 U566 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(N396) );
  OAI22_X1 U567 ( .A1(n3589), .A2(n4352), .B1(n3557), .B2(n4351), .ZN(n4081)
         );
  OAI22_X1 U568 ( .A1(n3525), .A2(n4354), .B1(n3333), .B2(n4353), .ZN(n4080)
         );
  OAI22_X1 U569 ( .A1(n3077), .A2(n4356), .B1(n3301), .B2(n4355), .ZN(n4079)
         );
  OAI22_X1 U570 ( .A1(n3269), .A2(n4358), .B1(n2821), .B2(n4357), .ZN(n4078)
         );
  NOR4_X1 U571 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .ZN(n4098) );
  OAI22_X1 U572 ( .A1(n3045), .A2(n4364), .B1(n3013), .B2(n4363), .ZN(n4085)
         );
  OAI22_X1 U573 ( .A1(n3461), .A2(n4366), .B1(n2789), .B2(n4365), .ZN(n4084)
         );
  OAI22_X1 U574 ( .A1(n2757), .A2(n4368), .B1(n3205), .B2(n4367), .ZN(n4083)
         );
  OAI22_X1 U575 ( .A1(n3429), .A2(n4370), .B1(n3397), .B2(n4369), .ZN(n4082)
         );
  NOR4_X1 U576 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4097) );
  OAI22_X1 U577 ( .A1(n2949), .A2(n4376), .B1(n3173), .B2(n4375), .ZN(n4089)
         );
  OAI22_X1 U578 ( .A1(n3141), .A2(n4378), .B1(n2693), .B2(n4377), .ZN(n4088)
         );
  OAI22_X1 U579 ( .A1(n2917), .A2(n4380), .B1(n2885), .B2(n4379), .ZN(n4087)
         );
  OAI22_X1 U580 ( .A1(n2661), .A2(n4382), .B1(n2629), .B2(n4381), .ZN(n4086)
         );
  NOR4_X1 U581 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4096) );
  OAI22_X1 U582 ( .A1(n3493), .A2(n4388), .B1(n3237), .B2(n3683), .ZN(n4093)
         );
  OAI22_X1 U583 ( .A1(n2981), .A2(n4389), .B1(n2725), .B2(n3672), .ZN(n4092)
         );
  OAI22_X1 U584 ( .A1(n3365), .A2(n4391), .B1(n3109), .B2(n4390), .ZN(n4091)
         );
  OAI22_X1 U585 ( .A1(n2853), .A2(n4393), .B1(n2597), .B2(n4392), .ZN(n4090)
         );
  OR4_X1 U586 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4094) );
  NAND2_X1 U587 ( .A1(n3685), .A2(n4094), .ZN(n4095) );
  NAND4_X1 U588 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(N397) );
  OAI22_X1 U589 ( .A1(n3588), .A2(n4352), .B1(n3556), .B2(n4351), .ZN(n4102)
         );
  OAI22_X1 U590 ( .A1(n3524), .A2(n4354), .B1(n3332), .B2(n3674), .ZN(n4101)
         );
  OAI22_X1 U591 ( .A1(n3076), .A2(n4356), .B1(n3300), .B2(n3675), .ZN(n4100)
         );
  OAI22_X1 U592 ( .A1(n3268), .A2(n3676), .B1(n2820), .B2(n4357), .ZN(n4099)
         );
  NOR4_X1 U593 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4119) );
  OAI22_X1 U594 ( .A1(n3044), .A2(n4364), .B1(n3012), .B2(n4363), .ZN(n4106)
         );
  OAI22_X1 U595 ( .A1(n3460), .A2(n3678), .B1(n2788), .B2(n3677), .ZN(n4105)
         );
  OAI22_X1 U596 ( .A1(n2756), .A2(n4368), .B1(n3204), .B2(n3679), .ZN(n4104)
         );
  OAI22_X1 U597 ( .A1(n3428), .A2(n3681), .B1(n3396), .B2(n3680), .ZN(n4103)
         );
  NOR4_X1 U598 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4118) );
  OAI22_X1 U599 ( .A1(n2948), .A2(n4376), .B1(n3172), .B2(n4375), .ZN(n4110)
         );
  OAI22_X1 U600 ( .A1(n3140), .A2(n4378), .B1(n2692), .B2(n4377), .ZN(n4109)
         );
  OAI22_X1 U601 ( .A1(n2916), .A2(n4380), .B1(n2884), .B2(n4379), .ZN(n4108)
         );
  OAI22_X1 U602 ( .A1(n2660), .A2(n4382), .B1(n2628), .B2(n3682), .ZN(n4107)
         );
  NOR4_X1 U603 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4117) );
  OAI22_X1 U604 ( .A1(n3492), .A2(n4388), .B1(n3236), .B2(n3683), .ZN(n4114)
         );
  OAI22_X1 U605 ( .A1(n2980), .A2(n4389), .B1(n2724), .B2(n3672), .ZN(n4113)
         );
  OAI22_X1 U606 ( .A1(n3364), .A2(n4391), .B1(n3108), .B2(n4390), .ZN(n4112)
         );
  OAI22_X1 U607 ( .A1(n2852), .A2(n4393), .B1(n2596), .B2(n4392), .ZN(n4111)
         );
  OR4_X1 U608 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4115) );
  NAND2_X1 U609 ( .A1(n3685), .A2(n4115), .ZN(n4116) );
  NAND4_X1 U610 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(N398) );
  OAI22_X1 U611 ( .A1(n3587), .A2(n4352), .B1(n3555), .B2(n4351), .ZN(n4123)
         );
  OAI22_X1 U612 ( .A1(n3523), .A2(n4354), .B1(n3331), .B2(n4353), .ZN(n4122)
         );
  OAI22_X1 U613 ( .A1(n3075), .A2(n4356), .B1(n3299), .B2(n4355), .ZN(n4121)
         );
  OAI22_X1 U614 ( .A1(n3267), .A2(n4358), .B1(n2819), .B2(n4357), .ZN(n4120)
         );
  NOR4_X1 U615 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4140) );
  OAI22_X1 U616 ( .A1(n3043), .A2(n4364), .B1(n3011), .B2(n4363), .ZN(n4127)
         );
  OAI22_X1 U617 ( .A1(n3459), .A2(n4366), .B1(n2787), .B2(n4365), .ZN(n4126)
         );
  OAI22_X1 U618 ( .A1(n2755), .A2(n4368), .B1(n3203), .B2(n4367), .ZN(n4125)
         );
  OAI22_X1 U619 ( .A1(n3427), .A2(n4370), .B1(n3395), .B2(n4369), .ZN(n4124)
         );
  NOR4_X1 U620 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4139) );
  OAI22_X1 U621 ( .A1(n2947), .A2(n4376), .B1(n3171), .B2(n4375), .ZN(n4131)
         );
  OAI22_X1 U622 ( .A1(n3139), .A2(n4378), .B1(n2691), .B2(n4377), .ZN(n4130)
         );
  OAI22_X1 U623 ( .A1(n2915), .A2(n4380), .B1(n2883), .B2(n4379), .ZN(n4129)
         );
  OAI22_X1 U624 ( .A1(n2659), .A2(n4382), .B1(n2627), .B2(n4381), .ZN(n4128)
         );
  NOR4_X1 U625 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4138) );
  OAI22_X1 U626 ( .A1(n3491), .A2(n4388), .B1(n3235), .B2(n3683), .ZN(n4135)
         );
  OAI22_X1 U627 ( .A1(n2979), .A2(n4389), .B1(n2723), .B2(n3672), .ZN(n4134)
         );
  OAI22_X1 U628 ( .A1(n3363), .A2(n4391), .B1(n3107), .B2(n4390), .ZN(n4133)
         );
  OAI22_X1 U629 ( .A1(n2851), .A2(n4393), .B1(n2595), .B2(n4392), .ZN(n4132)
         );
  OR4_X1 U630 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4136) );
  NAND2_X1 U631 ( .A1(n3685), .A2(n4136), .ZN(n4137) );
  NAND4_X1 U632 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(N399) );
  OAI22_X1 U633 ( .A1(n3586), .A2(n4352), .B1(n3554), .B2(n4351), .ZN(n4144)
         );
  OAI22_X1 U634 ( .A1(n3522), .A2(n4354), .B1(n3330), .B2(n3674), .ZN(n4143)
         );
  OAI22_X1 U635 ( .A1(n3074), .A2(n4356), .B1(n3298), .B2(n3675), .ZN(n4142)
         );
  OAI22_X1 U636 ( .A1(n3266), .A2(n3676), .B1(n2818), .B2(n4357), .ZN(n4141)
         );
  NOR4_X1 U637 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4161) );
  OAI22_X1 U638 ( .A1(n3042), .A2(n4364), .B1(n3010), .B2(n4363), .ZN(n4148)
         );
  OAI22_X1 U639 ( .A1(n3458), .A2(n3678), .B1(n2786), .B2(n3677), .ZN(n4147)
         );
  OAI22_X1 U640 ( .A1(n2754), .A2(n4368), .B1(n3202), .B2(n3679), .ZN(n4146)
         );
  OAI22_X1 U641 ( .A1(n3426), .A2(n3681), .B1(n3394), .B2(n3680), .ZN(n4145)
         );
  NOR4_X1 U642 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4160) );
  OAI22_X1 U643 ( .A1(n2946), .A2(n4376), .B1(n3170), .B2(n4375), .ZN(n4152)
         );
  OAI22_X1 U644 ( .A1(n3138), .A2(n4378), .B1(n2690), .B2(n4377), .ZN(n4151)
         );
  OAI22_X1 U645 ( .A1(n2914), .A2(n4380), .B1(n2882), .B2(n4379), .ZN(n4150)
         );
  OAI22_X1 U646 ( .A1(n2658), .A2(n4382), .B1(n2626), .B2(n3682), .ZN(n4149)
         );
  NOR4_X1 U647 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4159) );
  OAI22_X1 U648 ( .A1(n3490), .A2(n4388), .B1(n3234), .B2(n3683), .ZN(n4156)
         );
  OAI22_X1 U649 ( .A1(n2978), .A2(n4389), .B1(n2722), .B2(n3672), .ZN(n4155)
         );
  OAI22_X1 U650 ( .A1(n3362), .A2(n4391), .B1(n3106), .B2(n4390), .ZN(n4154)
         );
  OAI22_X1 U651 ( .A1(n2850), .A2(n4393), .B1(n2594), .B2(n4392), .ZN(n4153)
         );
  OR4_X1 U652 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157) );
  NAND2_X1 U653 ( .A1(n3685), .A2(n4157), .ZN(n4158) );
  NAND4_X1 U654 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(N400) );
  OAI22_X1 U655 ( .A1(n3585), .A2(n4352), .B1(n3553), .B2(n4351), .ZN(n4165)
         );
  OAI22_X1 U656 ( .A1(n3521), .A2(n4354), .B1(n3329), .B2(n4353), .ZN(n4164)
         );
  OAI22_X1 U657 ( .A1(n3073), .A2(n4356), .B1(n3297), .B2(n4355), .ZN(n4163)
         );
  OAI22_X1 U658 ( .A1(n3265), .A2(n4358), .B1(n2817), .B2(n4357), .ZN(n4162)
         );
  NOR4_X1 U659 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4182) );
  OAI22_X1 U660 ( .A1(n3041), .A2(n4364), .B1(n3009), .B2(n4363), .ZN(n4169)
         );
  OAI22_X1 U661 ( .A1(n3457), .A2(n4366), .B1(n2785), .B2(n4365), .ZN(n4168)
         );
  OAI22_X1 U662 ( .A1(n2753), .A2(n4368), .B1(n3201), .B2(n4367), .ZN(n4167)
         );
  OAI22_X1 U663 ( .A1(n3425), .A2(n4370), .B1(n3393), .B2(n4369), .ZN(n4166)
         );
  NOR4_X1 U664 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4181) );
  OAI22_X1 U665 ( .A1(n2945), .A2(n4376), .B1(n3169), .B2(n4375), .ZN(n4173)
         );
  OAI22_X1 U666 ( .A1(n3137), .A2(n4378), .B1(n2689), .B2(n4377), .ZN(n4172)
         );
  OAI22_X1 U667 ( .A1(n2913), .A2(n4380), .B1(n2881), .B2(n4379), .ZN(n4171)
         );
  OAI22_X1 U668 ( .A1(n2657), .A2(n4382), .B1(n2625), .B2(n4381), .ZN(n4170)
         );
  NOR4_X1 U669 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4180) );
  OAI22_X1 U670 ( .A1(n3489), .A2(n4388), .B1(n3233), .B2(n3683), .ZN(n4177)
         );
  OAI22_X1 U671 ( .A1(n2977), .A2(n4389), .B1(n2721), .B2(n3672), .ZN(n4176)
         );
  OAI22_X1 U672 ( .A1(n3361), .A2(n4391), .B1(n3105), .B2(n4390), .ZN(n4175)
         );
  OAI22_X1 U673 ( .A1(n2849), .A2(n4393), .B1(n2593), .B2(n4392), .ZN(n4174)
         );
  OR4_X1 U674 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4178) );
  NAND2_X1 U675 ( .A1(n4399), .A2(n4178), .ZN(n4179) );
  NAND4_X1 U676 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(N401) );
  OAI22_X1 U677 ( .A1(n3584), .A2(n4352), .B1(n3552), .B2(n4351), .ZN(n4186)
         );
  OAI22_X1 U678 ( .A1(n3520), .A2(n4354), .B1(n3328), .B2(n4353), .ZN(n4185)
         );
  OAI22_X1 U679 ( .A1(n3072), .A2(n4356), .B1(n3296), .B2(n4355), .ZN(n4184)
         );
  OAI22_X1 U680 ( .A1(n3264), .A2(n4358), .B1(n2816), .B2(n4357), .ZN(n4183)
         );
  NOR4_X1 U681 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4203) );
  OAI22_X1 U682 ( .A1(n3040), .A2(n4364), .B1(n3008), .B2(n4363), .ZN(n4190)
         );
  OAI22_X1 U683 ( .A1(n3456), .A2(n4366), .B1(n2784), .B2(n4365), .ZN(n4189)
         );
  OAI22_X1 U684 ( .A1(n2752), .A2(n4368), .B1(n3200), .B2(n4367), .ZN(n4188)
         );
  OAI22_X1 U685 ( .A1(n3424), .A2(n4370), .B1(n3392), .B2(n4369), .ZN(n4187)
         );
  NOR4_X1 U686 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4202) );
  OAI22_X1 U687 ( .A1(n2944), .A2(n4376), .B1(n3168), .B2(n4375), .ZN(n4194)
         );
  OAI22_X1 U688 ( .A1(n3136), .A2(n4378), .B1(n2688), .B2(n4377), .ZN(n4193)
         );
  OAI22_X1 U689 ( .A1(n2912), .A2(n4380), .B1(n2880), .B2(n4379), .ZN(n4192)
         );
  OAI22_X1 U690 ( .A1(n2656), .A2(n4382), .B1(n2624), .B2(n4381), .ZN(n4191)
         );
  NOR4_X1 U691 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4201) );
  OAI22_X1 U692 ( .A1(n3488), .A2(n4388), .B1(n3232), .B2(n3683), .ZN(n4198)
         );
  OAI22_X1 U693 ( .A1(n2976), .A2(n4389), .B1(n2720), .B2(n3672), .ZN(n4197)
         );
  OAI22_X1 U694 ( .A1(n3360), .A2(n4391), .B1(n3104), .B2(n4390), .ZN(n4196)
         );
  OAI22_X1 U695 ( .A1(n2848), .A2(n4393), .B1(n2592), .B2(n4392), .ZN(n4195)
         );
  OR4_X1 U696 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4199) );
  NAND2_X1 U697 ( .A1(n4399), .A2(n4199), .ZN(n4200) );
  NAND4_X1 U698 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(N402) );
  OAI22_X1 U699 ( .A1(n3583), .A2(n4352), .B1(n3551), .B2(n4351), .ZN(n4207)
         );
  OAI22_X1 U700 ( .A1(n3519), .A2(n4354), .B1(n3327), .B2(n3674), .ZN(n4206)
         );
  OAI22_X1 U701 ( .A1(n3071), .A2(n4356), .B1(n3295), .B2(n3675), .ZN(n4205)
         );
  OAI22_X1 U702 ( .A1(n3263), .A2(n3676), .B1(n2815), .B2(n4357), .ZN(n4204)
         );
  NOR4_X1 U703 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4224) );
  OAI22_X1 U704 ( .A1(n3039), .A2(n4364), .B1(n3007), .B2(n4363), .ZN(n4211)
         );
  OAI22_X1 U705 ( .A1(n3455), .A2(n3678), .B1(n2783), .B2(n3677), .ZN(n4210)
         );
  OAI22_X1 U706 ( .A1(n2751), .A2(n4368), .B1(n3199), .B2(n3679), .ZN(n4209)
         );
  OAI22_X1 U707 ( .A1(n3423), .A2(n3681), .B1(n3391), .B2(n3680), .ZN(n4208)
         );
  NOR4_X1 U708 ( .A1(n4211), .A2(n4210), .A3(n4209), .A4(n4208), .ZN(n4223) );
  OAI22_X1 U709 ( .A1(n2943), .A2(n4376), .B1(n3167), .B2(n4375), .ZN(n4215)
         );
  OAI22_X1 U710 ( .A1(n3135), .A2(n4378), .B1(n2687), .B2(n4377), .ZN(n4214)
         );
  OAI22_X1 U711 ( .A1(n2911), .A2(n4380), .B1(n2879), .B2(n4379), .ZN(n4213)
         );
  OAI22_X1 U712 ( .A1(n2655), .A2(n4382), .B1(n2623), .B2(n3682), .ZN(n4212)
         );
  NOR4_X1 U713 ( .A1(n4215), .A2(n4214), .A3(n4213), .A4(n4212), .ZN(n4222) );
  OAI22_X1 U714 ( .A1(n3487), .A2(n4388), .B1(n3231), .B2(n4387), .ZN(n4219)
         );
  OAI22_X1 U715 ( .A1(n2975), .A2(n4389), .B1(n2719), .B2(n3672), .ZN(n4218)
         );
  OAI22_X1 U716 ( .A1(n3359), .A2(n4391), .B1(n3103), .B2(n4390), .ZN(n4217)
         );
  OAI22_X1 U717 ( .A1(n2847), .A2(n4393), .B1(n2591), .B2(n4392), .ZN(n4216)
         );
  OR4_X1 U718 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4220) );
  NAND2_X1 U719 ( .A1(n3685), .A2(n4220), .ZN(n4221) );
  NAND4_X1 U720 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(N403) );
  OAI22_X1 U721 ( .A1(n3582), .A2(n4352), .B1(n3550), .B2(n4351), .ZN(n4228)
         );
  OAI22_X1 U722 ( .A1(n3518), .A2(n4354), .B1(n3326), .B2(n3674), .ZN(n4227)
         );
  OAI22_X1 U723 ( .A1(n3070), .A2(n4356), .B1(n3294), .B2(n3675), .ZN(n4226)
         );
  OAI22_X1 U724 ( .A1(n3262), .A2(n3676), .B1(n2814), .B2(n4357), .ZN(n4225)
         );
  NOR4_X1 U725 ( .A1(n4228), .A2(n4227), .A3(n4226), .A4(n4225), .ZN(n4245) );
  OAI22_X1 U726 ( .A1(n3038), .A2(n4364), .B1(n3006), .B2(n4363), .ZN(n4232)
         );
  OAI22_X1 U727 ( .A1(n3454), .A2(n3678), .B1(n2782), .B2(n3677), .ZN(n4231)
         );
  OAI22_X1 U728 ( .A1(n2750), .A2(n4368), .B1(n3198), .B2(n3679), .ZN(n4230)
         );
  OAI22_X1 U729 ( .A1(n3422), .A2(n3681), .B1(n3390), .B2(n3680), .ZN(n4229)
         );
  NOR4_X1 U730 ( .A1(n4232), .A2(n4231), .A3(n4230), .A4(n4229), .ZN(n4244) );
  OAI22_X1 U731 ( .A1(n2942), .A2(n4376), .B1(n3166), .B2(n4375), .ZN(n4236)
         );
  OAI22_X1 U732 ( .A1(n3134), .A2(n4378), .B1(n2686), .B2(n4377), .ZN(n4235)
         );
  OAI22_X1 U733 ( .A1(n2910), .A2(n4380), .B1(n2878), .B2(n4379), .ZN(n4234)
         );
  OAI22_X1 U734 ( .A1(n2654), .A2(n4382), .B1(n2622), .B2(n3682), .ZN(n4233)
         );
  NOR4_X1 U735 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4243) );
  OAI22_X1 U736 ( .A1(n3486), .A2(n4388), .B1(n3230), .B2(n4387), .ZN(n4240)
         );
  OAI22_X1 U737 ( .A1(n2974), .A2(n4389), .B1(n2718), .B2(n3672), .ZN(n4239)
         );
  OAI22_X1 U738 ( .A1(n3358), .A2(n4391), .B1(n3102), .B2(n4390), .ZN(n4238)
         );
  OAI22_X1 U739 ( .A1(n2846), .A2(n4393), .B1(n2590), .B2(n4392), .ZN(n4237)
         );
  OR4_X1 U740 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4241) );
  NAND2_X1 U741 ( .A1(n3685), .A2(n4241), .ZN(n4242) );
  NAND4_X1 U742 ( .A1(n4245), .A2(n4244), .A3(n4243), .A4(n4242), .ZN(N404) );
  OAI22_X1 U743 ( .A1(n3581), .A2(n4352), .B1(n3549), .B2(n4351), .ZN(n4249)
         );
  OAI22_X1 U744 ( .A1(n3517), .A2(n4354), .B1(n3325), .B2(n3674), .ZN(n4248)
         );
  OAI22_X1 U745 ( .A1(n3069), .A2(n4356), .B1(n3293), .B2(n3675), .ZN(n4247)
         );
  OAI22_X1 U746 ( .A1(n3261), .A2(n3676), .B1(n2813), .B2(n4357), .ZN(n4246)
         );
  NOR4_X1 U747 ( .A1(n4249), .A2(n4248), .A3(n4247), .A4(n4246), .ZN(n4266) );
  OAI22_X1 U748 ( .A1(n3037), .A2(n4364), .B1(n3005), .B2(n4363), .ZN(n4253)
         );
  OAI22_X1 U749 ( .A1(n3453), .A2(n3678), .B1(n2781), .B2(n3677), .ZN(n4252)
         );
  OAI22_X1 U750 ( .A1(n2749), .A2(n4368), .B1(n3197), .B2(n3679), .ZN(n4251)
         );
  OAI22_X1 U751 ( .A1(n3421), .A2(n3681), .B1(n3389), .B2(n3680), .ZN(n4250)
         );
  NOR4_X1 U752 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4250), .ZN(n4265) );
  OAI22_X1 U753 ( .A1(n2941), .A2(n4376), .B1(n3165), .B2(n4375), .ZN(n4257)
         );
  OAI22_X1 U754 ( .A1(n3133), .A2(n4378), .B1(n2685), .B2(n4377), .ZN(n4256)
         );
  OAI22_X1 U755 ( .A1(n2909), .A2(n4380), .B1(n2877), .B2(n4379), .ZN(n4255)
         );
  OAI22_X1 U756 ( .A1(n2653), .A2(n4382), .B1(n2621), .B2(n3682), .ZN(n4254)
         );
  NOR4_X1 U757 ( .A1(n4257), .A2(n4256), .A3(n4255), .A4(n4254), .ZN(n4264) );
  OAI22_X1 U758 ( .A1(n3485), .A2(n4388), .B1(n3229), .B2(n4387), .ZN(n4261)
         );
  OAI22_X1 U759 ( .A1(n2973), .A2(n4389), .B1(n2717), .B2(n3672), .ZN(n4260)
         );
  OAI22_X1 U760 ( .A1(n3357), .A2(n4391), .B1(n3101), .B2(n4390), .ZN(n4259)
         );
  OAI22_X1 U761 ( .A1(n2845), .A2(n4393), .B1(n2589), .B2(n4392), .ZN(n4258)
         );
  OR4_X1 U762 ( .A1(n4261), .A2(n4260), .A3(n4259), .A4(n4258), .ZN(n4262) );
  NAND2_X1 U763 ( .A1(n3685), .A2(n4262), .ZN(n4263) );
  NAND4_X1 U764 ( .A1(n4266), .A2(n4265), .A3(n4264), .A4(n4263), .ZN(N405) );
  OAI22_X1 U765 ( .A1(n3580), .A2(n4352), .B1(n3548), .B2(n4351), .ZN(n4270)
         );
  OAI22_X1 U766 ( .A1(n3516), .A2(n4354), .B1(n3324), .B2(n3674), .ZN(n4269)
         );
  OAI22_X1 U767 ( .A1(n3068), .A2(n4356), .B1(n3292), .B2(n3675), .ZN(n4268)
         );
  OAI22_X1 U768 ( .A1(n3260), .A2(n3676), .B1(n2812), .B2(n4357), .ZN(n4267)
         );
  NOR4_X1 U769 ( .A1(n4270), .A2(n4269), .A3(n4268), .A4(n4267), .ZN(n4287) );
  OAI22_X1 U770 ( .A1(n3036), .A2(n4364), .B1(n3004), .B2(n4363), .ZN(n4274)
         );
  OAI22_X1 U771 ( .A1(n3452), .A2(n3678), .B1(n2780), .B2(n3677), .ZN(n4273)
         );
  OAI22_X1 U772 ( .A1(n2748), .A2(n4368), .B1(n3196), .B2(n3679), .ZN(n4272)
         );
  OAI22_X1 U773 ( .A1(n3420), .A2(n3681), .B1(n3388), .B2(n3680), .ZN(n4271)
         );
  NOR4_X1 U774 ( .A1(n4274), .A2(n4273), .A3(n4272), .A4(n4271), .ZN(n4286) );
  OAI22_X1 U775 ( .A1(n2940), .A2(n4376), .B1(n3164), .B2(n4375), .ZN(n4278)
         );
  OAI22_X1 U776 ( .A1(n3132), .A2(n4378), .B1(n2684), .B2(n4377), .ZN(n4277)
         );
  OAI22_X1 U777 ( .A1(n2908), .A2(n4380), .B1(n2876), .B2(n4379), .ZN(n4276)
         );
  OAI22_X1 U778 ( .A1(n2652), .A2(n4382), .B1(n2620), .B2(n3682), .ZN(n4275)
         );
  NOR4_X1 U779 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(n4285) );
  OAI22_X1 U780 ( .A1(n3484), .A2(n4388), .B1(n3228), .B2(n4387), .ZN(n4282)
         );
  OAI22_X1 U781 ( .A1(n2972), .A2(n4389), .B1(n2716), .B2(n3672), .ZN(n4281)
         );
  OAI22_X1 U782 ( .A1(n3356), .A2(n4391), .B1(n3100), .B2(n4390), .ZN(n4280)
         );
  OAI22_X1 U783 ( .A1(n2844), .A2(n4393), .B1(n2588), .B2(n4392), .ZN(n4279)
         );
  OR4_X1 U784 ( .A1(n4282), .A2(n4281), .A3(n4280), .A4(n4279), .ZN(n4283) );
  NAND2_X1 U785 ( .A1(n3685), .A2(n4283), .ZN(n4284) );
  NAND4_X1 U786 ( .A1(n4287), .A2(n4286), .A3(n4285), .A4(n4284), .ZN(N406) );
  OAI22_X1 U787 ( .A1(n3579), .A2(n4352), .B1(n3547), .B2(n4351), .ZN(n4291)
         );
  OAI22_X1 U788 ( .A1(n3515), .A2(n4354), .B1(n3323), .B2(n3674), .ZN(n4290)
         );
  OAI22_X1 U789 ( .A1(n3067), .A2(n4356), .B1(n3291), .B2(n3675), .ZN(n4289)
         );
  OAI22_X1 U790 ( .A1(n3259), .A2(n3676), .B1(n2811), .B2(n4357), .ZN(n4288)
         );
  NOR4_X1 U791 ( .A1(n4291), .A2(n4290), .A3(n4289), .A4(n4288), .ZN(n4308) );
  OAI22_X1 U792 ( .A1(n3035), .A2(n4364), .B1(n3003), .B2(n4363), .ZN(n4295)
         );
  OAI22_X1 U793 ( .A1(n3451), .A2(n3678), .B1(n2779), .B2(n3677), .ZN(n4294)
         );
  OAI22_X1 U794 ( .A1(n2747), .A2(n4368), .B1(n3195), .B2(n3679), .ZN(n4293)
         );
  OAI22_X1 U795 ( .A1(n3419), .A2(n3681), .B1(n3387), .B2(n3680), .ZN(n4292)
         );
  NOR4_X1 U796 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4307) );
  OAI22_X1 U797 ( .A1(n2939), .A2(n4376), .B1(n3163), .B2(n4375), .ZN(n4299)
         );
  OAI22_X1 U798 ( .A1(n3131), .A2(n4378), .B1(n2683), .B2(n4377), .ZN(n4298)
         );
  OAI22_X1 U799 ( .A1(n2907), .A2(n4380), .B1(n2875), .B2(n4379), .ZN(n4297)
         );
  OAI22_X1 U800 ( .A1(n2651), .A2(n4382), .B1(n2619), .B2(n3682), .ZN(n4296)
         );
  NOR4_X1 U801 ( .A1(n4299), .A2(n4298), .A3(n4297), .A4(n4296), .ZN(n4306) );
  OAI22_X1 U802 ( .A1(n3483), .A2(n4388), .B1(n3227), .B2(n4387), .ZN(n4303)
         );
  OAI22_X1 U803 ( .A1(n2971), .A2(n4389), .B1(n2715), .B2(n3672), .ZN(n4302)
         );
  OAI22_X1 U804 ( .A1(n3355), .A2(n4391), .B1(n3099), .B2(n4390), .ZN(n4301)
         );
  OAI22_X1 U805 ( .A1(n2843), .A2(n4393), .B1(n2587), .B2(n4392), .ZN(n4300)
         );
  OR4_X1 U806 ( .A1(n4303), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(n4304) );
  NAND2_X1 U807 ( .A1(n3685), .A2(n4304), .ZN(n4305) );
  NAND4_X1 U808 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), .ZN(N407) );
  OAI22_X1 U809 ( .A1(n3578), .A2(n4352), .B1(n3546), .B2(n4351), .ZN(n4312)
         );
  OAI22_X1 U810 ( .A1(n3514), .A2(n4354), .B1(n3322), .B2(n3674), .ZN(n4311)
         );
  OAI22_X1 U811 ( .A1(n3066), .A2(n4356), .B1(n3290), .B2(n3675), .ZN(n4310)
         );
  OAI22_X1 U812 ( .A1(n3258), .A2(n3676), .B1(n2810), .B2(n4357), .ZN(n4309)
         );
  NOR4_X1 U813 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4329) );
  OAI22_X1 U814 ( .A1(n3034), .A2(n4364), .B1(n3002), .B2(n4363), .ZN(n4316)
         );
  OAI22_X1 U815 ( .A1(n3450), .A2(n3678), .B1(n2778), .B2(n3677), .ZN(n4315)
         );
  OAI22_X1 U816 ( .A1(n2746), .A2(n4368), .B1(n3194), .B2(n3679), .ZN(n4314)
         );
  OAI22_X1 U817 ( .A1(n3418), .A2(n3681), .B1(n3386), .B2(n3680), .ZN(n4313)
         );
  NOR4_X1 U818 ( .A1(n4316), .A2(n4315), .A3(n4314), .A4(n4313), .ZN(n4328) );
  OAI22_X1 U819 ( .A1(n2938), .A2(n4376), .B1(n3162), .B2(n4375), .ZN(n4320)
         );
  OAI22_X1 U820 ( .A1(n3130), .A2(n4378), .B1(n2682), .B2(n4377), .ZN(n4319)
         );
  OAI22_X1 U821 ( .A1(n2906), .A2(n4380), .B1(n2874), .B2(n4379), .ZN(n4318)
         );
  OAI22_X1 U822 ( .A1(n2650), .A2(n4382), .B1(n2618), .B2(n3682), .ZN(n4317)
         );
  NOR4_X1 U823 ( .A1(n4320), .A2(n4319), .A3(n4318), .A4(n4317), .ZN(n4327) );
  OAI22_X1 U824 ( .A1(n3482), .A2(n4388), .B1(n3226), .B2(n4387), .ZN(n4324)
         );
  OAI22_X1 U825 ( .A1(n2970), .A2(n4389), .B1(n2714), .B2(n3672), .ZN(n4323)
         );
  OAI22_X1 U826 ( .A1(n3354), .A2(n4391), .B1(n3098), .B2(n4390), .ZN(n4322)
         );
  OAI22_X1 U827 ( .A1(n2842), .A2(n4393), .B1(n2586), .B2(n4392), .ZN(n4321)
         );
  OR4_X1 U828 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(n4325) );
  NAND2_X1 U829 ( .A1(n3685), .A2(n4325), .ZN(n4326) );
  NAND4_X1 U830 ( .A1(n4329), .A2(n4328), .A3(n4327), .A4(n4326), .ZN(N408) );
  OAI22_X1 U831 ( .A1(n3577), .A2(n4352), .B1(n3545), .B2(n4351), .ZN(n4333)
         );
  OAI22_X1 U832 ( .A1(n3513), .A2(n4354), .B1(n3321), .B2(n3674), .ZN(n4332)
         );
  OAI22_X1 U833 ( .A1(n3065), .A2(n4356), .B1(n3289), .B2(n3675), .ZN(n4331)
         );
  OAI22_X1 U834 ( .A1(n3257), .A2(n3676), .B1(n2809), .B2(n4357), .ZN(n4330)
         );
  NOR4_X1 U835 ( .A1(n4333), .A2(n4332), .A3(n4331), .A4(n4330), .ZN(n4350) );
  OAI22_X1 U836 ( .A1(n3033), .A2(n4364), .B1(n3001), .B2(n4363), .ZN(n4337)
         );
  OAI22_X1 U837 ( .A1(n3449), .A2(n3678), .B1(n2777), .B2(n3677), .ZN(n4336)
         );
  OAI22_X1 U838 ( .A1(n2745), .A2(n4368), .B1(n3193), .B2(n3679), .ZN(n4335)
         );
  OAI22_X1 U839 ( .A1(n3417), .A2(n3681), .B1(n3385), .B2(n3680), .ZN(n4334)
         );
  NOR4_X1 U840 ( .A1(n4337), .A2(n4336), .A3(n4335), .A4(n4334), .ZN(n4349) );
  OAI22_X1 U841 ( .A1(n2937), .A2(n4376), .B1(n3161), .B2(n4375), .ZN(n4341)
         );
  OAI22_X1 U842 ( .A1(n3129), .A2(n4378), .B1(n2681), .B2(n4377), .ZN(n4340)
         );
  OAI22_X1 U843 ( .A1(n2905), .A2(n4380), .B1(n2873), .B2(n4379), .ZN(n4339)
         );
  OAI22_X1 U844 ( .A1(n2649), .A2(n4382), .B1(n2617), .B2(n3682), .ZN(n4338)
         );
  NOR4_X1 U845 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4348) );
  OAI22_X1 U846 ( .A1(n3481), .A2(n4388), .B1(n3225), .B2(n4387), .ZN(n4345)
         );
  OAI22_X1 U847 ( .A1(n2969), .A2(n4389), .B1(n2713), .B2(n3672), .ZN(n4344)
         );
  OAI22_X1 U848 ( .A1(n3353), .A2(n4391), .B1(n3097), .B2(n4390), .ZN(n4343)
         );
  OAI22_X1 U849 ( .A1(n2841), .A2(n4393), .B1(n2585), .B2(n4392), .ZN(n4342)
         );
  OR4_X1 U850 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4346) );
  NAND2_X1 U851 ( .A1(n3685), .A2(n4346), .ZN(n4347) );
  NAND4_X1 U852 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(N409) );
  OAI22_X1 U853 ( .A1(n3576), .A2(n4352), .B1(n3544), .B2(n4351), .ZN(n4362)
         );
  OAI22_X1 U854 ( .A1(n3512), .A2(n4354), .B1(n3320), .B2(n3674), .ZN(n4361)
         );
  OAI22_X1 U855 ( .A1(n3064), .A2(n4356), .B1(n3288), .B2(n3675), .ZN(n4360)
         );
  OAI22_X1 U856 ( .A1(n3256), .A2(n3676), .B1(n2808), .B2(n4357), .ZN(n4359)
         );
  NOR4_X1 U857 ( .A1(n4362), .A2(n4361), .A3(n4360), .A4(n4359), .ZN(n4403) );
  OAI22_X1 U858 ( .A1(n3032), .A2(n4364), .B1(n3000), .B2(n4363), .ZN(n4374)
         );
  OAI22_X1 U859 ( .A1(n3448), .A2(n3678), .B1(n2776), .B2(n3677), .ZN(n4373)
         );
  OAI22_X1 U860 ( .A1(n2744), .A2(n4368), .B1(n3192), .B2(n3679), .ZN(n4372)
         );
  OAI22_X1 U861 ( .A1(n3416), .A2(n3681), .B1(n3384), .B2(n3680), .ZN(n4371)
         );
  NOR4_X1 U862 ( .A1(n4374), .A2(n4373), .A3(n4372), .A4(n4371), .ZN(n4402) );
  OAI22_X1 U863 ( .A1(n2936), .A2(n4376), .B1(n3160), .B2(n4375), .ZN(n4386)
         );
  OAI22_X1 U864 ( .A1(n3128), .A2(n4378), .B1(n2680), .B2(n4377), .ZN(n4385)
         );
  OAI22_X1 U865 ( .A1(n2904), .A2(n4380), .B1(n2872), .B2(n4379), .ZN(n4384)
         );
  OAI22_X1 U866 ( .A1(n2648), .A2(n4382), .B1(n2616), .B2(n3682), .ZN(n4383)
         );
  NOR4_X1 U867 ( .A1(n4386), .A2(n4385), .A3(n4384), .A4(n4383), .ZN(n4401) );
  OAI22_X1 U868 ( .A1(n3480), .A2(n4388), .B1(n3224), .B2(n4387), .ZN(n4397)
         );
  OAI22_X1 U869 ( .A1(n2968), .A2(n4389), .B1(n2712), .B2(n3672), .ZN(n4396)
         );
  OAI22_X1 U870 ( .A1(n3352), .A2(n4391), .B1(n3096), .B2(n4390), .ZN(n4395)
         );
  OAI22_X1 U871 ( .A1(n2840), .A2(n4393), .B1(n2584), .B2(n4392), .ZN(n4394)
         );
  OR4_X1 U872 ( .A1(n4397), .A2(n4396), .A3(n4395), .A4(n4394), .ZN(n4398) );
  NAND2_X1 U873 ( .A1(n3685), .A2(n4398), .ZN(n4400) );
  NAND4_X1 U874 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(N410) );
  NAND3_X1 U875 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(ADD_WR[1]), .ZN(n4414)
         );
  NAND3_X1 U876 ( .A1(n4413), .A2(ADD_WR[4]), .A3(ADD_WR[3]), .ZN(n4408) );
  INV_X1 U877 ( .A(ADD_WR[0]), .ZN(n4404) );
  NAND3_X1 U878 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .A3(n4404), .ZN(n4415) );
  OAI21_X1 U879 ( .B1(n4408), .B2(n4415), .A(n3662), .ZN(n31) );
  NOR2_X1 U880 ( .A1(ADD_WR[1]), .A2(n4404), .ZN(n4405) );
  NAND2_X1 U881 ( .A1(ADD_WR[2]), .A2(n4405), .ZN(n4416) );
  OAI21_X1 U882 ( .B1(n4408), .B2(n4416), .A(n3661), .ZN(n30) );
  NOR2_X1 U883 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .ZN(n4407) );
  NAND2_X1 U884 ( .A1(ADD_WR[2]), .A2(n4407), .ZN(n4417) );
  OAI21_X1 U885 ( .B1(n4408), .B2(n4417), .A(n3660), .ZN(n29) );
  NAND3_X1 U886 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n4406), .ZN(n4418) );
  OAI21_X1 U887 ( .B1(n4408), .B2(n4418), .A(n3659), .ZN(n28) );
  NAND3_X1 U888 ( .A1(ADD_WR[1]), .A2(n4406), .A3(n4404), .ZN(n4419) );
  OAI21_X1 U889 ( .B1(n4408), .B2(n4419), .A(n3658), .ZN(n27) );
  NAND2_X1 U890 ( .A1(n4405), .A2(n4406), .ZN(n4420) );
  OAI21_X1 U891 ( .B1(n4408), .B2(n4420), .A(n3657), .ZN(n26) );
  NAND2_X1 U892 ( .A1(n4407), .A2(n4406), .ZN(n4422) );
  OAI21_X1 U893 ( .B1(n4408), .B2(n4422), .A(n3656), .ZN(n25) );
  INV_X1 U894 ( .A(ADD_WR[3]), .ZN(n4411) );
  NAND3_X1 U895 ( .A1(ADD_WR[4]), .A2(n4413), .A3(n4411), .ZN(n4409) );
  OAI21_X1 U896 ( .B1(n4414), .B2(n4409), .A(n3667), .ZN(n24) );
  OAI21_X1 U897 ( .B1(n4415), .B2(n4409), .A(n3622), .ZN(n23) );
  OAI21_X1 U898 ( .B1(n4416), .B2(n4409), .A(n3621), .ZN(n22) );
  OAI21_X1 U899 ( .B1(n4417), .B2(n4409), .A(n3666), .ZN(n21) );
  OAI21_X1 U900 ( .B1(n4418), .B2(n4409), .A(n3620), .ZN(n20) );
  OAI21_X1 U901 ( .B1(n4419), .B2(n4409), .A(n3619), .ZN(n19) );
  OAI21_X1 U902 ( .B1(n4420), .B2(n4409), .A(n3665), .ZN(n18) );
  OAI21_X1 U903 ( .B1(n4422), .B2(n4409), .A(n3618), .ZN(n17) );
  INV_X1 U904 ( .A(ADD_WR[4]), .ZN(n4412) );
  NAND3_X1 U905 ( .A1(n4413), .A2(ADD_WR[3]), .A3(n4412), .ZN(n4410) );
  OAI21_X1 U906 ( .B1(n4414), .B2(n4410), .A(n3664), .ZN(n16) );
  OAI21_X1 U907 ( .B1(n4415), .B2(n4410), .A(n3663), .ZN(n15) );
  OAI21_X1 U908 ( .B1(n4416), .B2(n4410), .A(n3617), .ZN(n14) );
  OAI21_X1 U909 ( .B1(n4417), .B2(n4410), .A(n3616), .ZN(n13) );
  OAI21_X1 U910 ( .B1(n4418), .B2(n4410), .A(n3668), .ZN(n12) );
  OAI21_X1 U911 ( .B1(n4419), .B2(n4410), .A(n3669), .ZN(n11) );
  NAND3_X1 U912 ( .A1(n4413), .A2(n4412), .A3(n4411), .ZN(n4421) );
  OAI21_X1 U913 ( .B1(n4419), .B2(n4421), .A(n3670), .ZN(n3) );
  OAI21_X1 U914 ( .B1(n4420), .B2(n4421), .A(n3671), .ZN(n2) );
  OAI21_X1 U915 ( .B1(n4422), .B2(n4421), .A(n3623), .ZN(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net79314, n2, n3;
  assign net79314 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net79314), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net79314, n2, n3;
  assign net79314 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net79314), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net79314, n2, n3;
  assign net79314 = EN;

  AND2_X1 main_gate ( .A1(n2), .A2(CLK), .ZN(ENCLK) );
  OR2_X1 U1 ( .A1(TE), .A2(net79314), .ZN(n3) );
  DLL_X1 U2 ( .D(n3), .GN(CLK), .Q(n2) );
endmodule


module dlx ( RST, CLK );
  input RST, CLK;
  wire   \cw_dec[2] , \cw_mem[4] , \unit_control/n153 , \unit_control/n152 ,
         \unit_control/cw2delay[4] , \unit_control/cw2delay[3] ,
         \unit_control/cw1delay[17] , \unit_control/cw1delay[14] ,
         \unit_control/cw1delay[13] , \unit_control/cw1delay[12] ,
         \unit_control/cw1delay[10] , \unit_control/cw1delay[9] ,
         \unit_control/cw1delay[4] , \unit_control/cw1delay[3] ,
         \unit_control/next_state[1] , \unit_control/next_state[0] ,
         \unit_fetch/adder_out[31] , \unit_fetch/adder_out[30] ,
         \unit_fetch/adder_out[29] , \unit_fetch/adder_out[28] ,
         \unit_fetch/adder_out[27] , \unit_fetch/adder_out[26] ,
         \unit_fetch/adder_out[25] , \unit_fetch/adder_out[24] ,
         \unit_fetch/adder_out[23] , \unit_fetch/adder_out[22] ,
         \unit_fetch/adder_out[21] , \unit_fetch/adder_out[20] ,
         \unit_fetch/adder_out[19] , \unit_fetch/adder_out[18] ,
         \unit_fetch/adder_out[17] , \unit_fetch/adder_out[16] ,
         \unit_fetch/adder_out[15] , \unit_fetch/adder_out[14] ,
         \unit_fetch/adder_out[13] , \unit_fetch/adder_out[12] ,
         \unit_fetch/adder_out[11] , \unit_fetch/adder_out[10] ,
         \unit_fetch/adder_out[9] , \unit_fetch/adder_out[8] ,
         \unit_fetch/adder_out[7] , \unit_fetch/adder_out[6] ,
         \unit_fetch/adder_out[5] , \unit_fetch/adder_out[4] ,
         \unit_fetch/adder_out[3] , \unit_fetch/pc_regout[0] ,
         \unit_fetch/pc_regout[1] , \unit_fetch/pc_regout[2] ,
         \unit_fetch/pc_regout[3] , \unit_fetch/pc_regout[4] ,
         \unit_fetch/pc_regout[5] , \unit_fetch/pc_regout[6] ,
         \unit_fetch/pc_regout[7] , \unit_fetch/pc_regout[8] ,
         \unit_fetch/pc_regout[9] , \unit_fetch/pc_regout[10] ,
         \unit_fetch/pc_regout[11] , \unit_fetch/pc_regout[12] ,
         \unit_fetch/pc_regout[13] , \unit_fetch/pc_regout[14] ,
         \unit_fetch/pc_regout[15] , \unit_fetch/pc_regout[16] ,
         \unit_fetch/pc_regout[17] , \unit_fetch/pc_regout[18] ,
         \unit_fetch/pc_regout[19] , \unit_fetch/pc_regout[21] ,
         \unit_fetch/pc_regout[22] , \unit_fetch/pc_regout[23] ,
         \unit_fetch/pc_regout[24] , \unit_fetch/pc_regout[25] ,
         \unit_fetch/pc_regout[26] , \unit_fetch/pc_regout[27] ,
         \unit_fetch/pc_regout[28] , \unit_fetch/pc_regout[29] ,
         \unit_fetch/pc_regout[30] , \unit_decode/registerA[31] ,
         \unit_decode/registerA[30] , \unit_decode/registerA[29] ,
         \unit_decode/registerA[28] , \unit_decode/registerA[27] ,
         \unit_decode/registerA[26] , \unit_decode/registerA[25] ,
         \unit_decode/registerA[24] , \unit_decode/registerA[23] ,
         \unit_decode/registerA[22] , \unit_decode/registerA[21] ,
         \unit_decode/registerA[20] , \unit_decode/registerA[19] ,
         \unit_decode/registerA[18] , \unit_decode/registerA[17] ,
         \unit_decode/registerA[16] , \unit_decode/registerA[15] ,
         \unit_decode/registerA[14] , \unit_decode/registerA[13] ,
         \unit_decode/registerA[12] , \unit_decode/registerA[11] ,
         \unit_decode/registerA[10] , \unit_decode/registerA[9] ,
         \unit_decode/registerA[8] , \unit_decode/registerA[7] ,
         \unit_decode/registerA[6] , \unit_decode/registerA[5] ,
         \unit_decode/registerA[4] , \unit_decode/registerA[3] ,
         \unit_decode/registerA[2] , \unit_decode/registerA[1] ,
         \unit_decode/registerA[0] , \unit_decode/RS1s[4] ,
         \unit_decode/RS1s[3] , \unit_decode/RS1s[2] , \unit_decode/RS1s[1] ,
         \unit_fetch/unit_instructionRegister/n98 ,
         \unit_fetch/unit_instructionRegister/n97 ,
         \unit_fetch/unit_instructionRegister/n96 ,
         \unit_fetch/unit_instructionRegister/n95 ,
         \unit_fetch/unit_instructionRegister/n94 ,
         \unit_fetch/unit_instructionRegister/n93 ,
         \unit_fetch/unit_instructionRegister/n91 ,
         \unit_fetch/unit_instructionRegister/n90 ,
         \unit_fetch/unit_instructionRegister/n89 ,
         \unit_fetch/unit_instructionRegister/n88 ,
         \unit_fetch/unit_instructionRegister/n87 ,
         \unit_fetch/unit_instructionRegister/n86 ,
         \unit_fetch/unit_instructionRegister/n85 ,
         \unit_fetch/unit_instructionRegister/n83 ,
         \unit_fetch/unit_instructionRegister/n82 ,
         \unit_fetch/unit_instructionRegister/n81 ,
         \unit_fetch/unit_instructionRegister/n80 ,
         \unit_fetch/unit_instructionRegister/n79 ,
         \unit_fetch/unit_instructionRegister/n78 ,
         \unit_fetch/unit_instructionRegister/n77 ,
         \unit_fetch/unit_instructionRegister/n75 ,
         \unit_fetch/unit_instructionRegister/n74 ,
         \unit_fetch/unit_instructionRegister/n73 ,
         \unit_fetch/unit_instructionRegister/n72 ,
         \unit_fetch/unit_instructionRegister/n71 ,
         \unit_fetch/unit_instructionRegister/n70 ,
         \unit_fetch/unit_instructionRegister/n68 ,
         \unit_fetch/unit_instructionRegister/n67 ,
         \unit_fetch/unit_instructionRegister/n66 ,
         \unit_fetch/unit_instructionRegister/n65 ,
         \unit_fetch/unit_instructionRegister/n64 ,
         \unit_fetch/unit_instructionRegister/n63 ,
         \unit_fetch/unit_instructionRegister/n62 ,
         \unit_fetch/unit_instructionRegister/n61 ,
         \unit_fetch/unit_instructionRegister/n60 ,
         \unit_fetch/unit_instructionRegister/n59 ,
         \unit_fetch/unit_instructionRegister/n57 ,
         \unit_fetch/unit_instructionRegister/n56 ,
         \unit_fetch/unit_instructionRegister/n55 ,
         \unit_fetch/unit_instructionRegister/n54 ,
         \unit_fetch/unit_instructionRegister/n53 ,
         \unit_fetch/unit_instructionRegister/n51 ,
         \unit_fetch/unit_instructionRegister/n50 ,
         \unit_fetch/unit_instructionRegister/n49 ,
         \unit_fetch/unit_instructionRegister/n48 ,
         \unit_fetch/unit_instructionRegister/n47 ,
         \unit_fetch/unit_instructionRegister/n46 ,
         \unit_fetch/unit_instructionRegister/n45 ,
         \unit_fetch/unit_instructionRegister/n43 ,
         \unit_fetch/unit_instructionRegister/n42 ,
         \unit_fetch/unit_instructionRegister/n41 ,
         \unit_fetch/unit_instructionRegister/n40 ,
         \unit_fetch/unit_instructionRegister/n39 ,
         \unit_fetch/unit_instructionRegister/n38 ,
         \unit_control/uut_second_stage/ffi_24/n3 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_0/n5 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_1/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_2/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_3/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_4/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_5/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_6/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_7/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_8/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_9/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_10/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_11/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_12/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_13/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_14/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_15/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_16/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_17/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_18/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_19/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_20/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_21/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_22/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_23/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_24/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_25/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_26/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_27/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_28/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_29/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_30/n4 ,
         \unit_execution/COMP_REGN_ALUOUT/ffi_31/n4 ,
         \unit_execution/COMP_NPC2/ffi_0/n4 ,
         \unit_execution/COMP_NPC2/ffi_1/n4 ,
         \unit_execution/COMP_NPC2/ffi_2/n4 ,
         \unit_execution/COMP_NPC2/ffi_3/n4 ,
         \unit_execution/COMP_NPC2/ffi_4/n4 ,
         \unit_execution/COMP_NPC2/ffi_5/n4 ,
         \unit_execution/COMP_NPC2/ffi_6/n4 ,
         \unit_execution/COMP_NPC2/ffi_7/n4 ,
         \unit_execution/COMP_NPC2/ffi_8/n4 ,
         \unit_execution/COMP_NPC2/ffi_9/n4 ,
         \unit_execution/COMP_NPC2/ffi_10/n4 ,
         \unit_execution/COMP_NPC2/ffi_11/n4 ,
         \unit_execution/COMP_NPC2/ffi_12/n4 ,
         \unit_execution/COMP_NPC2/ffi_13/n4 ,
         \unit_execution/COMP_NPC2/ffi_14/n4 ,
         \unit_execution/COMP_NPC2/ffi_15/n4 ,
         \unit_execution/COMP_NPC2/ffi_16/n4 ,
         \unit_execution/COMP_NPC2/ffi_17/n4 ,
         \unit_execution/COMP_NPC2/ffi_18/n4 ,
         \unit_execution/COMP_NPC2/ffi_19/n4 ,
         \unit_execution/COMP_NPC2/ffi_20/n4 ,
         \unit_execution/COMP_NPC2/ffi_21/n4 ,
         \unit_execution/COMP_NPC2/ffi_22/n4 ,
         \unit_execution/COMP_NPC2/ffi_23/n4 ,
         \unit_execution/COMP_NPC2/ffi_24/n4 ,
         \unit_execution/COMP_NPC2/ffi_25/n4 ,
         \unit_execution/COMP_NPC2/ffi_26/n4 ,
         \unit_execution/COMP_NPC2/ffi_27/n4 ,
         \unit_execution/COMP_NPC2/ffi_28/n4 ,
         \unit_execution/COMP_NPC2/ffi_29/n4 ,
         \unit_execution/COMP_NPC2/ffi_30/n4 ,
         \unit_execution/COMP_NPC2/ffi_31/n4 , \unit_decode/RD1reg/ffi_0/n4 ,
         \unit_decode/RD1reg/ffi_1/n4 , \unit_decode/RD1reg/ffi_2/n4 ,
         \unit_decode/RD1reg/ffi_3/n4 , \unit_decode/RD1reg/ffi_4/n4 ,
         \unit_decode/IMMreg/ffi_0/n4 , \unit_decode/IMMreg/ffi_2/n4 ,
         \unit_decode/IMMreg/ffi_3/n4 , \unit_decode/IMMreg/ffi_5/n4 ,
         \unit_decode/IMMreg/ffi_6/n4 , \unit_decode/IMMreg/ffi_7/n4 ,
         \unit_decode/IMMreg/ffi_8/n4 , \unit_decode/IMMreg/ffi_9/n4 ,
         \unit_decode/IMMreg/ffi_11/n4 , \unit_decode/IMMreg/ffi_13/n4 ,
         \unit_decode/IMMreg/ffi_14/n4 , \unit_decode/IMMreg/ffi_15/n4 ,
         \unit_decode/IMMreg/ffi_16/n5 , \unit_decode/IMMreg/ffi_16/n4 ,
         \unit_decode/IMMreg/ffi_17/n5 , \unit_decode/IMMreg/ffi_17/n4 ,
         \unit_decode/IMMreg/ffi_18/n5 , \unit_decode/IMMreg/ffi_18/n4 ,
         \unit_decode/IMMreg/ffi_19/n5 , \unit_decode/IMMreg/ffi_19/n4 ,
         \unit_decode/IMMreg/ffi_20/n5 , \unit_decode/IMMreg/ffi_20/n4 ,
         \unit_decode/IMMreg/ffi_21/n5 , \unit_decode/IMMreg/ffi_21/n4 ,
         \unit_decode/IMMreg/ffi_22/n5 , \unit_decode/IMMreg/ffi_22/n4 ,
         \unit_decode/IMMreg/ffi_23/n5 , \unit_decode/IMMreg/ffi_23/n4 ,
         \unit_decode/IMMreg/ffi_24/n5 , \unit_decode/IMMreg/ffi_24/n4 ,
         \unit_decode/IMMreg/ffi_25/n5 , \unit_decode/IMMreg/ffi_25/n4 ,
         \unit_decode/IMMreg/ffi_31/n4 , \unit_decode/Areg/ffi_0/n4 ,
         \unit_decode/Areg/ffi_1/n4 , \unit_decode/Areg/ffi_2/n4 ,
         \unit_decode/Areg/ffi_3/n4 , \unit_decode/Areg/ffi_4/n4 ,
         \unit_decode/Areg/ffi_5/n4 , \unit_decode/Areg/ffi_6/n4 ,
         \unit_decode/Areg/ffi_7/n4 , \unit_decode/Areg/ffi_9/n4 ,
         \unit_decode/Areg/ffi_10/n4 , \unit_decode/Areg/ffi_11/n4 ,
         \unit_decode/Areg/ffi_12/n4 , \unit_decode/Areg/ffi_13/n4 ,
         \unit_decode/Areg/ffi_14/n4 , \unit_decode/Areg/ffi_15/n4 ,
         \unit_decode/Areg/ffi_16/n4 , \unit_decode/Areg/ffi_17/n4 ,
         \unit_decode/Areg/ffi_18/n4 , \unit_decode/Areg/ffi_20/n4 ,
         \unit_decode/Areg/ffi_21/n4 , \unit_decode/Areg/ffi_22/n4 ,
         \unit_decode/Areg/ffi_23/n4 , \unit_decode/Areg/ffi_24/n4 ,
         \unit_decode/Areg/ffi_25/n4 , \unit_decode/Areg/ffi_26/n4 ,
         \unit_decode/Areg/ffi_27/n4 , \unit_decode/Areg/ffi_28/n4 ,
         \unit_decode/Areg/ffi_29/n4 , \unit_decode/Areg/ffi_30/n4 ,
         \unit_decode/Areg/ffi_31/n4 , \unit_decode/NPC1reg/ffi_0/n4 ,
         \unit_decode/NPC1reg/ffi_1/n4 , \unit_decode/NPC1reg/ffi_2/n4 ,
         \unit_decode/NPC1reg/ffi_3/n4 , \unit_decode/NPC1reg/ffi_4/n4 ,
         \unit_decode/NPC1reg/ffi_5/n4 , \unit_decode/NPC1reg/ffi_6/n4 ,
         \unit_decode/NPC1reg/ffi_7/n4 , \unit_decode/NPC1reg/ffi_8/n4 ,
         \unit_decode/NPC1reg/ffi_9/n4 , \unit_decode/NPC1reg/ffi_10/n4 ,
         \unit_decode/NPC1reg/ffi_11/n4 , \unit_decode/NPC1reg/ffi_12/n4 ,
         \unit_decode/NPC1reg/ffi_13/n4 , \unit_decode/NPC1reg/ffi_14/n4 ,
         \unit_decode/NPC1reg/ffi_15/n4 , \unit_decode/NPC1reg/ffi_16/n4 ,
         \unit_decode/NPC1reg/ffi_17/n4 , \unit_decode/NPC1reg/ffi_18/n4 ,
         \unit_decode/NPC1reg/ffi_19/n4 , \unit_decode/NPC1reg/ffi_20/n4 ,
         \unit_decode/NPC1reg/ffi_21/n4 , \unit_decode/NPC1reg/ffi_22/n4 ,
         \unit_decode/NPC1reg/ffi_23/n4 , \unit_decode/NPC1reg/ffi_24/n4 ,
         \unit_decode/NPC1reg/ffi_25/n4 , \unit_decode/NPC1reg/ffi_26/n4 ,
         \unit_decode/NPC1reg/ffi_27/n4 , \unit_decode/NPC1reg/ffi_28/n4 ,
         \unit_decode/NPC1reg/ffi_29/n4 , \unit_decode/NPC1reg/ffi_30/n4 ,
         \unit_decode/NPC1reg/ffi_31/n4 ,
         \unit_fetch/unit_npcregister/ffi_0/n5 ,
         \unit_fetch/unit_npcregister/ffi_0/n4 ,
         \unit_fetch/unit_npcregister/ffi_1/n5 ,
         \unit_fetch/unit_npcregister/ffi_1/n4 ,
         \unit_fetch/unit_npcregister/ffi_2/n5 ,
         \unit_fetch/unit_npcregister/ffi_2/n4 ,
         \unit_fetch/unit_npcregister/ffi_3/n5 ,
         \unit_fetch/unit_npcregister/ffi_3/n4 ,
         \unit_fetch/unit_npcregister/ffi_4/n5 ,
         \unit_fetch/unit_npcregister/ffi_4/n4 ,
         \unit_fetch/unit_npcregister/ffi_5/n5 ,
         \unit_fetch/unit_npcregister/ffi_5/n4 ,
         \unit_fetch/unit_npcregister/ffi_6/n5 ,
         \unit_fetch/unit_npcregister/ffi_6/n4 ,
         \unit_fetch/unit_npcregister/ffi_7/n5 ,
         \unit_fetch/unit_npcregister/ffi_7/n4 ,
         \unit_fetch/unit_npcregister/ffi_8/n5 ,
         \unit_fetch/unit_npcregister/ffi_8/n4 ,
         \unit_fetch/unit_npcregister/ffi_9/n5 ,
         \unit_fetch/unit_npcregister/ffi_9/n4 ,
         \unit_fetch/unit_npcregister/ffi_10/n5 ,
         \unit_fetch/unit_npcregister/ffi_10/n4 ,
         \unit_fetch/unit_npcregister/ffi_11/n5 ,
         \unit_fetch/unit_npcregister/ffi_11/n4 ,
         \unit_fetch/unit_npcregister/ffi_12/n5 ,
         \unit_fetch/unit_npcregister/ffi_12/n4 ,
         \unit_fetch/unit_npcregister/ffi_13/n5 ,
         \unit_fetch/unit_npcregister/ffi_13/n4 ,
         \unit_fetch/unit_npcregister/ffi_14/n5 ,
         \unit_fetch/unit_npcregister/ffi_14/n4 ,
         \unit_fetch/unit_npcregister/ffi_15/n5 ,
         \unit_fetch/unit_npcregister/ffi_15/n4 ,
         \unit_fetch/unit_npcregister/ffi_16/n5 ,
         \unit_fetch/unit_npcregister/ffi_16/n4 ,
         \unit_fetch/unit_npcregister/ffi_17/n5 ,
         \unit_fetch/unit_npcregister/ffi_17/n4 ,
         \unit_fetch/unit_npcregister/ffi_18/n5 ,
         \unit_fetch/unit_npcregister/ffi_18/n4 ,
         \unit_fetch/unit_npcregister/ffi_19/n5 ,
         \unit_fetch/unit_npcregister/ffi_19/n4 ,
         \unit_fetch/unit_npcregister/ffi_20/n5 ,
         \unit_fetch/unit_npcregister/ffi_20/n4 ,
         \unit_fetch/unit_npcregister/ffi_21/n5 ,
         \unit_fetch/unit_npcregister/ffi_21/n4 ,
         \unit_fetch/unit_npcregister/ffi_22/n5 ,
         \unit_fetch/unit_npcregister/ffi_22/n4 ,
         \unit_fetch/unit_npcregister/ffi_23/n5 ,
         \unit_fetch/unit_npcregister/ffi_23/n4 ,
         \unit_fetch/unit_npcregister/ffi_24/n5 ,
         \unit_fetch/unit_npcregister/ffi_24/n4 ,
         \unit_fetch/unit_npcregister/ffi_25/n5 ,
         \unit_fetch/unit_npcregister/ffi_25/n4 ,
         \unit_fetch/unit_npcregister/ffi_26/n5 ,
         \unit_fetch/unit_npcregister/ffi_26/n4 ,
         \unit_fetch/unit_npcregister/ffi_27/n5 ,
         \unit_fetch/unit_npcregister/ffi_27/n4 ,
         \unit_fetch/unit_npcregister/ffi_28/n5 ,
         \unit_fetch/unit_npcregister/ffi_28/n4 ,
         \unit_fetch/unit_npcregister/ffi_29/n5 ,
         \unit_fetch/unit_npcregister/ffi_29/n4 ,
         \unit_fetch/unit_npcregister/ffi_30/n5 ,
         \unit_fetch/unit_npcregister/ffi_30/n4 ,
         \unit_fetch/unit_npcregister/ffi_31/n5 ,
         \unit_fetch/unit_npcregister/ffi_31/n4 ,
         \unit_fetch/unit_programCounter/ffi_0/n5 ,
         \unit_fetch/unit_programCounter/ffi_0/n4 ,
         \unit_fetch/unit_programCounter/ffi_1/n5 ,
         \unit_fetch/unit_programCounter/ffi_1/n4 ,
         \unit_fetch/unit_programCounter/ffi_2/n5 ,
         \unit_fetch/unit_programCounter/ffi_2/n4 ,
         \unit_fetch/unit_programCounter/ffi_3/n5 ,
         \unit_fetch/unit_programCounter/ffi_3/n4 ,
         \unit_fetch/unit_programCounter/ffi_4/n5 ,
         \unit_fetch/unit_programCounter/ffi_4/n4 ,
         \unit_fetch/unit_programCounter/ffi_5/n5 ,
         \unit_fetch/unit_programCounter/ffi_5/n4 ,
         \unit_fetch/unit_programCounter/ffi_6/n5 ,
         \unit_fetch/unit_programCounter/ffi_6/n4 ,
         \unit_fetch/unit_programCounter/ffi_7/n5 ,
         \unit_fetch/unit_programCounter/ffi_7/n4 ,
         \unit_fetch/unit_programCounter/ffi_8/n5 ,
         \unit_fetch/unit_programCounter/ffi_8/n4 ,
         \unit_fetch/unit_programCounter/ffi_9/n5 ,
         \unit_fetch/unit_programCounter/ffi_9/n4 ,
         \unit_fetch/unit_programCounter/ffi_10/n5 ,
         \unit_fetch/unit_programCounter/ffi_10/n4 ,
         \unit_fetch/unit_programCounter/ffi_11/n5 ,
         \unit_fetch/unit_programCounter/ffi_11/n4 ,
         \unit_fetch/unit_programCounter/ffi_12/n5 ,
         \unit_fetch/unit_programCounter/ffi_12/n4 ,
         \unit_fetch/unit_programCounter/ffi_13/n5 ,
         \unit_fetch/unit_programCounter/ffi_14/n5 ,
         \unit_fetch/unit_programCounter/ffi_14/n4 ,
         \unit_fetch/unit_programCounter/ffi_15/n5 ,
         \unit_fetch/unit_programCounter/ffi_15/n4 ,
         \unit_fetch/unit_programCounter/ffi_16/n5 ,
         \unit_fetch/unit_programCounter/ffi_16/n4 ,
         \unit_fetch/unit_programCounter/ffi_17/n5 ,
         \unit_fetch/unit_programCounter/ffi_17/n4 ,
         \unit_fetch/unit_programCounter/ffi_18/n5 ,
         \unit_fetch/unit_programCounter/ffi_18/n4 ,
         \unit_fetch/unit_programCounter/ffi_19/n5 ,
         \unit_fetch/unit_programCounter/ffi_19/n4 ,
         \unit_fetch/unit_programCounter/ffi_20/n5 ,
         \unit_fetch/unit_programCounter/ffi_20/n4 ,
         \unit_fetch/unit_programCounter/ffi_21/n5 ,
         \unit_fetch/unit_programCounter/ffi_21/n4 ,
         \unit_fetch/unit_programCounter/ffi_22/n5 ,
         \unit_fetch/unit_programCounter/ffi_22/n4 ,
         \unit_fetch/unit_programCounter/ffi_23/n5 ,
         \unit_fetch/unit_programCounter/ffi_23/n4 ,
         \unit_fetch/unit_programCounter/ffi_24/n5 ,
         \unit_fetch/unit_programCounter/ffi_24/n4 ,
         \unit_fetch/unit_programCounter/ffi_25/n5 ,
         \unit_fetch/unit_programCounter/ffi_25/n4 ,
         \unit_fetch/unit_programCounter/ffi_26/n5 ,
         \unit_fetch/unit_programCounter/ffi_26/n4 ,
         \unit_fetch/unit_programCounter/ffi_27/n5 ,
         \unit_fetch/unit_programCounter/ffi_27/n4 ,
         \unit_fetch/unit_programCounter/ffi_28/n5 ,
         \unit_fetch/unit_programCounter/ffi_28/n4 ,
         \unit_fetch/unit_programCounter/ffi_29/n5 ,
         \unit_fetch/unit_programCounter/ffi_29/n4 ,
         \unit_fetch/unit_programCounter/ffi_30/n5 ,
         \unit_fetch/unit_programCounter/ffi_30/n4 ,
         \unit_fetch/unit_programCounter/ffi_31/n5 ,
         \unit_control/uut_fourth_stage/ffi_3/n6 ,
         \unit_control/uut_fourth_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_3/n5 ,
         \unit_control/uut_third_stage/ffi_4/n5 ,
         \unit_control/uut_third_stage/ffi_9/n6 ,
         \unit_control/uut_third_stage/ffi_9/n5 ,
         \unit_control/uut_third_stage/ffi_10/n5 ,
         \unit_control/uut_third_stage/ffi_12/n5 ,
         \unit_control/uut_third_stage/ffi_13/n5 ,
         \unit_control/uut_third_stage/ffi_14/n5 ,
         \unit_control/uut_third_stage/ffi_15/n5 ,
         \unit_control/uut_third_stage/ffi_17/n6 ,
         \unit_control/uut_third_stage/ffi_17/n5 ,
         \unit_control/uut_third_stage/ffi_19/n5 ,
         \unit_control/uut_second_stage/ffi_3/n5 ,
         \unit_control/uut_second_stage/ffi_10/n5 ,
         \unit_control/uut_second_stage/ffi_12/n5 ,
         \unit_control/uut_second_stage/ffi_13/n5 ,
         \unit_control/uut_second_stage/ffi_14/n5 ,
         \unit_control/uut_second_stage/ffi_17/n5 ,
         \unit_control/uut_second_stage/ffi_21/n5 , n4, n6, n471, n1330, n1331,
         n1333, n1336, n1337, n1338, n1340, n1341, n1342,
         \unit_fetch/unit_adder/add_19/n89 ,
         \unit_fetch/unit_adder/add_19/n86 ,
         \unit_fetch/unit_adder/add_19/n85 ,
         \unit_fetch/unit_adder/add_19/n84 ,
         \unit_fetch/unit_adder/add_19/n82 ,
         \unit_fetch/unit_adder/add_19/n81 ,
         \unit_fetch/unit_adder/add_19/n79 ,
         \unit_fetch/unit_adder/add_19/n78 ,
         \unit_fetch/unit_adder/add_19/n77 ,
         \unit_fetch/unit_adder/add_19/n73 ,
         \unit_fetch/unit_adder/add_19/n70 ,
         \unit_fetch/unit_adder/add_19/n69 ,
         \unit_fetch/unit_adder/add_19/n66 ,
         \unit_fetch/unit_adder/add_19/n63 ,
         \unit_fetch/unit_adder/add_19/n57 ,
         \unit_fetch/unit_adder/add_19/n54 ,
         \unit_fetch/unit_adder/add_19/n53 ,
         \unit_fetch/unit_adder/add_19/n52 ,
         \unit_fetch/unit_adder/add_19/n48 ,
         \unit_fetch/unit_adder/add_19/n47 ,
         \unit_fetch/unit_adder/add_19/n45 ,
         \unit_fetch/unit_adder/add_19/n44 ,
         \unit_fetch/unit_adder/add_19/n43 ,
         \unit_fetch/unit_adder/add_19/n42 ,
         \unit_fetch/unit_adder/add_19/n41 ,
         \unit_fetch/unit_adder/add_19/n38 ,
         \unit_fetch/unit_adder/add_19/n37 ,
         \unit_fetch/unit_adder/add_19/n35 ,
         \unit_fetch/unit_adder/add_19/n34 ,
         \unit_fetch/unit_adder/add_19/n33 ,
         \unit_fetch/unit_adder/add_19/n32 ,
         \unit_fetch/unit_adder/add_19/n29 ,
         \unit_fetch/unit_adder/add_19/n28 ,
         \unit_fetch/unit_adder/add_19/n18 ,
         \unit_fetch/unit_adder/add_19/n17 ,
         \unit_fetch/unit_adder/add_19/n15 ,
         \unit_fetch/unit_adder/add_19/n14 ,
         \unit_fetch/unit_adder/add_19/n12 , \unit_fetch/unit_adder/add_19/n9 ,
         \unit_fetch/unit_adder/add_19/n8 , \unit_fetch/unit_adder/add_19/n7 ,
         \unit_fetch/unit_adder/add_19/n6 , \unit_fetch/unit_adder/add_19/n5 ,
         \unit_fetch/unit_adder/add_19/n4 , \unit_fetch/unit_adder/add_19/n3 ,
         \unit_fetch/unit_adder/add_19/n2 , \unit_fetch/unit_adder/add_19/n1 ,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087;
  wire   [4:0] wr_address;
  wire   [31:0] wr_data;

  DFFR_X1 \unit_control/current_state_reg[1]  ( .D(
        \unit_control/next_state[1] ), .CK(CLK), .RN(n1942), .Q(
        \unit_control/n152 ) );
  DFFR_X1 \unit_control/current_state_reg[0]  ( .D(
        \unit_control/next_state[0] ), .CK(CLK), .RN(n1942), .Q(
        \unit_control/n153 ) );
  register_file_WORD_SIZE32_ADDR_SIZE5 \unit_decode/RegisterFile  ( .CLK(CLK), 
        .ENABLE(\cw_dec[2] ), .RD1(\unit_control/cw1delay[9] ), .RD2(1'b0), 
        .WR(\cw_mem[4] ), .ADD_WR(wr_address), .ADD_RD1({\unit_decode/RS1s[4] , 
        \unit_decode/RS1s[3] , \unit_decode/RS1s[2] , \unit_decode/RS1s[1] , 
        n1707}), .ADD_RD2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATAIN(wr_data), 
        .OUT1({\unit_decode/registerA[31] , \unit_decode/registerA[30] , 
        \unit_decode/registerA[29] , \unit_decode/registerA[28] , 
        \unit_decode/registerA[27] , \unit_decode/registerA[26] , 
        \unit_decode/registerA[25] , \unit_decode/registerA[24] , 
        \unit_decode/registerA[23] , \unit_decode/registerA[22] , 
        \unit_decode/registerA[21] , \unit_decode/registerA[20] , 
        \unit_decode/registerA[19] , \unit_decode/registerA[18] , 
        \unit_decode/registerA[17] , \unit_decode/registerA[16] , 
        \unit_decode/registerA[15] , \unit_decode/registerA[14] , 
        \unit_decode/registerA[13] , \unit_decode/registerA[12] , 
        \unit_decode/registerA[11] , \unit_decode/registerA[10] , 
        \unit_decode/registerA[9] , \unit_decode/registerA[8] , 
        \unit_decode/registerA[7] , \unit_decode/registerA[6] , 
        \unit_decode/registerA[5] , \unit_decode/registerA[4] , 
        \unit_decode/registerA[3] , \unit_decode/registerA[2] , 
        \unit_decode/registerA[1] , \unit_decode/registerA[0] }), .RESET(RST)
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[0]  ( .D(
        \unit_fetch/unit_instructionRegister/n98 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n38 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[1]  ( .D(
        \unit_fetch/unit_instructionRegister/n97 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n39 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[2]  ( .D(
        \unit_fetch/unit_instructionRegister/n96 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n40 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[3]  ( .D(
        \unit_fetch/unit_instructionRegister/n95 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n41 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[4]  ( .D(
        \unit_fetch/unit_instructionRegister/n94 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n42 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[5]  ( .D(
        \unit_fetch/unit_instructionRegister/n93 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n43 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[7]  ( .D(
        \unit_fetch/unit_instructionRegister/n91 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n45 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[8]  ( .D(
        \unit_fetch/unit_instructionRegister/n90 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n46 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[10]  ( .D(
        \unit_fetch/unit_instructionRegister/n88 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n48 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[11]  ( .D(
        \unit_fetch/unit_instructionRegister/n87 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n49 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[12]  ( .D(
        \unit_fetch/unit_instructionRegister/n86 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n50 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[13]  ( .D(
        \unit_fetch/unit_instructionRegister/n85 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n51 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[15]  ( .D(
        \unit_fetch/unit_instructionRegister/n83 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n53 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[16]  ( .D(
        \unit_fetch/unit_instructionRegister/n82 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n54 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[18]  ( .D(
        \unit_fetch/unit_instructionRegister/n80 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n56 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[19]  ( .D(
        \unit_fetch/unit_instructionRegister/n79 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n57 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[21]  ( .D(
        \unit_fetch/unit_instructionRegister/n77 ), .CK(CLK), .Q(n1707), .QN(
        \unit_fetch/unit_instructionRegister/n59 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[23]  ( .D(
        \unit_fetch/unit_instructionRegister/n67 ), .CK(CLK), .Q(
        \unit_decode/RS1s[2] ), .QN(\unit_fetch/unit_instructionRegister/n61 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[24]  ( .D(
        \unit_fetch/unit_instructionRegister/n75 ), .CK(CLK), .Q(
        \unit_decode/RS1s[3] ), .QN(\unit_fetch/unit_instructionRegister/n62 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[25]  ( .D(
        \unit_fetch/unit_instructionRegister/n74 ), .CK(CLK), .Q(
        \unit_decode/RS1s[4] ), .QN(\unit_fetch/unit_instructionRegister/n63 )
         );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[26]  ( .D(
        \unit_fetch/unit_instructionRegister/n68 ), .CK(CLK), .QN(n1333) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[27]  ( .D(
        \unit_fetch/unit_instructionRegister/n73 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n64 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[28]  ( .D(
        \unit_fetch/unit_instructionRegister/n70 ), .CK(CLK), .QN(n1331) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[29]  ( .D(
        \unit_fetch/unit_instructionRegister/n72 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n65 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[31]  ( .D(
        \unit_fetch/unit_instructionRegister/n71 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n66 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_0/Q_reg  ( .D(n2940), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_0/n5 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_2/Q_reg  ( .D(n2942), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_2/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_3/Q_reg  ( .D(n2943), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_3/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_4/Q_reg  ( .D(n2944), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_4/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_5/Q_reg  ( .D(n2945), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_5/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_6/Q_reg  ( .D(n2946), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_6/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_7/Q_reg  ( .D(n2947), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_7/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_8/Q_reg  ( .D(n2948), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_8/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_9/Q_reg  ( .D(n2949), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_9/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_10/Q_reg  ( .D(n2950), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_10/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_11/Q_reg  ( .D(n2951), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_11/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_12/Q_reg  ( .D(n2952), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_12/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_13/Q_reg  ( .D(n2953), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_13/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_14/Q_reg  ( .D(n2954), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_14/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_15/Q_reg  ( .D(n2955), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_15/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_16/Q_reg  ( .D(n2956), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_16/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_17/Q_reg  ( .D(n2957), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_17/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_18/Q_reg  ( .D(n2958), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_18/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_19/Q_reg  ( .D(n2959), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_19/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_20/Q_reg  ( .D(n2960), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_20/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_21/Q_reg  ( .D(n2961), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_21/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_22/Q_reg  ( .D(n2962), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_22/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_23/Q_reg  ( .D(n2963), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_23/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_24/Q_reg  ( .D(n2964), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_24/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_25/Q_reg  ( .D(n2965), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_25/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_26/Q_reg  ( .D(n2966), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_26/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_27/Q_reg  ( .D(n2967), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_27/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_28/Q_reg  ( .D(n2968), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_28/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_29/Q_reg  ( .D(n2969), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_29/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_30/Q_reg  ( .D(n2970), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_30/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_31/Q_reg  ( .D(n2971), .CK(n3004), .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_31/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_0/Q_reg  ( .D(n2972), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_0/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_1/Q_reg  ( .D(n2973), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_1/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_2/Q_reg  ( .D(n2974), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_2/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_3/Q_reg  ( .D(n2975), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_3/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_4/Q_reg  ( .D(n2976), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_4/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_5/Q_reg  ( .D(n2977), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_5/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_6/Q_reg  ( .D(n2978), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_6/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_7/Q_reg  ( .D(n2979), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_7/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_8/Q_reg  ( .D(n2980), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_8/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_9/Q_reg  ( .D(n2981), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_9/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_10/Q_reg  ( .D(n2982), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_10/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_11/Q_reg  ( .D(n2983), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_11/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_12/Q_reg  ( .D(n2984), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_12/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_13/Q_reg  ( .D(n2985), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_13/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_14/Q_reg  ( .D(n2986), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_14/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_15/Q_reg  ( .D(n2987), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_15/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_16/Q_reg  ( .D(n2988), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_16/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_17/Q_reg  ( .D(n2989), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_17/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_18/Q_reg  ( .D(n2990), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_18/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_19/Q_reg  ( .D(n2991), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_19/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_20/Q_reg  ( .D(n2992), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_20/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_21/Q_reg  ( .D(n2993), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_21/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_22/Q_reg  ( .D(n2994), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_22/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_23/Q_reg  ( .D(n2995), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_23/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_24/Q_reg  ( .D(n2996), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_24/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_25/Q_reg  ( .D(n2997), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_25/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_26/Q_reg  ( .D(n2998), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_26/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_27/Q_reg  ( .D(n2999), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_27/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_28/Q_reg  ( .D(n3000), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_28/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_29/Q_reg  ( .D(n3001), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_29/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_30/Q_reg  ( .D(n3002), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_30/n4 ) );
  DFF_X1 \unit_execution/COMP_NPC2/ffi_31/Q_reg  ( .D(n3003), .CK(n3004), .QN(
        \unit_execution/COMP_NPC2/ffi_31/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_0/Q_reg  ( .D(n3005), .CK(n3087), .QN(
        \unit_decode/RD1reg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_1/Q_reg  ( .D(n3006), .CK(n3087), .QN(
        \unit_decode/RD1reg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_2/Q_reg  ( .D(n3007), .CK(n3087), .QN(
        \unit_decode/RD1reg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_3/Q_reg  ( .D(n3008), .CK(n3087), .Q(n1683), 
        .QN(\unit_decode/RD1reg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/RD1reg/ffi_4/Q_reg  ( .D(n3009), .CK(n3087), .Q(n1654), 
        .QN(\unit_decode/RD1reg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_5/Q_reg  ( .D(n3014), .CK(n3087), .Q(n1680), 
        .QN(\unit_decode/IMMreg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_6/Q_reg  ( .D(n3013), .CK(n3087), .Q(n1652), 
        .QN(\unit_decode/IMMreg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_7/Q_reg  ( .D(n3015), .CK(n3087), .Q(n1556), 
        .QN(\unit_decode/IMMreg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_8/Q_reg  ( .D(n3016), .CK(n3087), .Q(n1681), 
        .QN(\unit_decode/IMMreg/ffi_8/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_9/Q_reg  ( .D(n3017), .CK(n3087), .Q(n1684), 
        .QN(\unit_decode/IMMreg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_11/Q_reg  ( .D(n3019), .CK(n3087), .QN(
        \unit_decode/IMMreg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_13/Q_reg  ( .D(n3021), .CK(n3087), .Q(n1672), 
        .QN(\unit_decode/IMMreg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_14/Q_reg  ( .D(n3020), .CK(n3087), .Q(n1663), 
        .QN(\unit_decode/IMMreg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_15/Q_reg  ( .D(n3022), .CK(n3087), .Q(n1669), 
        .QN(\unit_decode/IMMreg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_16/Q_reg  ( .D(\unit_decode/IMMreg/ffi_16/n5 ), .CK(n3087), .Q(n1668), .QN(\unit_decode/IMMreg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_17/Q_reg  ( .D(\unit_decode/IMMreg/ffi_17/n5 ), .CK(n3087), .Q(n1666), .QN(\unit_decode/IMMreg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_18/Q_reg  ( .D(\unit_decode/IMMreg/ffi_18/n5 ), .CK(n3087), .Q(n1679), .QN(\unit_decode/IMMreg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_19/Q_reg  ( .D(\unit_decode/IMMreg/ffi_19/n5 ), .CK(n3087), .Q(n1675), .QN(\unit_decode/IMMreg/ffi_19/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_20/Q_reg  ( .D(\unit_decode/IMMreg/ffi_20/n5 ), .CK(n3087), .Q(n1678), .QN(\unit_decode/IMMreg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_21/Q_reg  ( .D(\unit_decode/IMMreg/ffi_21/n5 ), .CK(n3087), .Q(n1682), .QN(\unit_decode/IMMreg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_22/Q_reg  ( .D(\unit_decode/IMMreg/ffi_22/n5 ), .CK(n3087), .QN(\unit_decode/IMMreg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_23/Q_reg  ( .D(\unit_decode/IMMreg/ffi_23/n5 ), .CK(n3087), .Q(n1674), .QN(\unit_decode/IMMreg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/IMMreg/ffi_24/Q_reg  ( .D(\unit_decode/IMMreg/ffi_24/n5 ), .CK(n3087), .Q(n1670), .QN(\unit_decode/IMMreg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_0/Q_reg  ( .D(n3023), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_1/Q_reg  ( .D(n3024), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_2/Q_reg  ( .D(n3025), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_3/Q_reg  ( .D(n3026), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_4/Q_reg  ( .D(n3027), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_5/Q_reg  ( .D(n3028), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_6/Q_reg  ( .D(n3029), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_7/Q_reg  ( .D(n3030), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_9/Q_reg  ( .D(n3032), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_10/Q_reg  ( .D(n3033), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_10/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_11/Q_reg  ( .D(n3034), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_12/Q_reg  ( .D(n3035), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_12/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_13/Q_reg  ( .D(n3036), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_14/Q_reg  ( .D(n3037), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_15/Q_reg  ( .D(n3038), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_16/Q_reg  ( .D(n3039), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_17/Q_reg  ( .D(n3040), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_18/Q_reg  ( .D(n3041), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_20/Q_reg  ( .D(n3043), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_21/Q_reg  ( .D(n3044), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_22/Q_reg  ( .D(n3045), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_23/Q_reg  ( .D(n3046), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_24/Q_reg  ( .D(n3047), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_25/Q_reg  ( .D(n3048), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_25/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_26/Q_reg  ( .D(n3049), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_26/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_27/Q_reg  ( .D(n3050), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_27/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_28/Q_reg  ( .D(n3051), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_28/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_29/Q_reg  ( .D(n3052), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_29/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_30/Q_reg  ( .D(n3053), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_30/n4 ) );
  DFF_X1 \unit_decode/Areg/ffi_31/Q_reg  ( .D(n3054), .CK(n3087), .QN(
        \unit_decode/Areg/ffi_31/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_0/Q_reg  ( .D(n3055), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_0/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_1/Q_reg  ( .D(n3056), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_1/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_2/Q_reg  ( .D(n3057), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_2/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_3/Q_reg  ( .D(n3058), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_3/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_4/Q_reg  ( .D(n3059), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_4/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_5/Q_reg  ( .D(n3060), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_5/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_6/Q_reg  ( .D(n3061), .CK(n3087), .Q(n1513), 
        .QN(\unit_decode/NPC1reg/ffi_6/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_7/Q_reg  ( .D(n3062), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_7/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_8/Q_reg  ( .D(n3063), .CK(n3087), .Q(n1648), 
        .QN(\unit_decode/NPC1reg/ffi_8/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_9/Q_reg  ( .D(n3064), .CK(n3087), .Q(n1515), 
        .QN(\unit_decode/NPC1reg/ffi_9/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_10/Q_reg  ( .D(n3065), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_10/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_11/Q_reg  ( .D(n3066), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_11/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_12/Q_reg  ( .D(n3067), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_12/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_13/Q_reg  ( .D(n3068), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_13/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_14/Q_reg  ( .D(n3069), .CK(n3087), .Q(n1514), 
        .QN(\unit_decode/NPC1reg/ffi_14/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_15/Q_reg  ( .D(n3070), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_15/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_16/Q_reg  ( .D(n3071), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_16/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_17/Q_reg  ( .D(n3072), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_17/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_18/Q_reg  ( .D(n3073), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_18/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_19/Q_reg  ( .D(n3074), .CK(n3087), .Q(n1644), 
        .QN(\unit_decode/NPC1reg/ffi_19/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_20/Q_reg  ( .D(n3075), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_20/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_21/Q_reg  ( .D(n3076), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_21/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_22/Q_reg  ( .D(n3077), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_22/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_23/Q_reg  ( .D(n3078), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_23/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_24/Q_reg  ( .D(n3079), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_24/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_25/Q_reg  ( .D(n3080), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_25/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_26/Q_reg  ( .D(n3081), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_26/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_27/Q_reg  ( .D(n3082), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_27/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_28/Q_reg  ( .D(n3083), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_28/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_29/Q_reg  ( .D(n3084), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_29/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_30/Q_reg  ( .D(n3085), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_30/n4 ) );
  DFF_X1 \unit_decode/NPC1reg/ffi_31/Q_reg  ( .D(n3086), .CK(n3087), .QN(
        \unit_decode/NPC1reg/ffi_31/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_1/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_1/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_1/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_2/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_2/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_2/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_3/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_3/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_3/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_4/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_4/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_4/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_5/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_5/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_5/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_6/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_6/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_6/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_7/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_7/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_7/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_8/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_8/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_8/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_9/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_9/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_9/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_10/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_10/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_10/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_11/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_11/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_11/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_12/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_12/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_12/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_13/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_13/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_13/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_14/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_14/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_14/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_15/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_15/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_15/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_16/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_16/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_16/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_17/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_17/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_17/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_18/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_18/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_18/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_20/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_20/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_20/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_21/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_21/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_21/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_22/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_22/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_22/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_23/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_23/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_23/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_24/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_24/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_24/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_25/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_25/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_25/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_26/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_26/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_26/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_27/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_27/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_27/n4 ) );
  DFF_X1 \unit_fetch/unit_npcregister/ffi_30/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_30/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_npcregister/ffi_30/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_1/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_1/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[1] ), .QN(
        \unit_fetch/unit_programCounter/ffi_1/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_3/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_3/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[3] ), .QN(
        \unit_fetch/unit_programCounter/ffi_3/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_4/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_4/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[4] ), .QN(
        \unit_fetch/unit_programCounter/ffi_4/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_5/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_5/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[5] ), .QN(
        \unit_fetch/unit_programCounter/ffi_5/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_7/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_7/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[7] ), .QN(
        \unit_fetch/unit_programCounter/ffi_7/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_8/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_8/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[8] ), .QN(
        \unit_fetch/unit_programCounter/ffi_8/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_9/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_9/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[9] ), .QN(
        \unit_fetch/unit_programCounter/ffi_9/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_10/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_10/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[10] ), .QN(
        \unit_fetch/unit_programCounter/ffi_10/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_11/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_11/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[11] ), .QN(
        \unit_fetch/unit_programCounter/ffi_11/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_12/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_12/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[12] ), .QN(
        \unit_fetch/unit_programCounter/ffi_12/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_14/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_14/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[14] ), .QN(
        \unit_fetch/unit_programCounter/ffi_14/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_15/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_15/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[15] ), .QN(
        \unit_fetch/unit_programCounter/ffi_15/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_16/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_16/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[16] ), .QN(
        \unit_fetch/unit_programCounter/ffi_16/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_17/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_17/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[17] ), .QN(
        \unit_fetch/unit_programCounter/ffi_17/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_18/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_18/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[18] ), .QN(
        \unit_fetch/unit_programCounter/ffi_18/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_19/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_19/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[19] ), .QN(
        \unit_fetch/unit_programCounter/ffi_19/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_20/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_20/n5 ), .CK(n2933), .QN(
        \unit_fetch/unit_programCounter/ffi_20/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_21/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_21/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[21] ), .QN(
        \unit_fetch/unit_programCounter/ffi_21/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_22/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_22/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[22] ), .QN(
        \unit_fetch/unit_programCounter/ffi_22/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_23/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_23/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[23] ), .QN(
        \unit_fetch/unit_programCounter/ffi_23/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_24/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_24/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[24] ), .QN(
        \unit_fetch/unit_programCounter/ffi_24/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_25/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_25/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[25] ), .QN(
        \unit_fetch/unit_programCounter/ffi_25/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_26/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_26/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[26] ), .QN(
        \unit_fetch/unit_programCounter/ffi_26/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_27/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_27/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[27] ), .QN(
        \unit_fetch/unit_programCounter/ffi_27/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_28/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_28/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[28] ), .QN(
        \unit_fetch/unit_programCounter/ffi_28/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_29/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_29/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[29] ), .QN(
        \unit_fetch/unit_programCounter/ffi_29/n4 ) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_30/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_30/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[30] ), .QN(
        \unit_fetch/unit_programCounter/ffi_30/n4 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_9/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_9/n6 ), .CK(CLK), .Q(n1915), .QN(
        \unit_control/uut_third_stage/ffi_9/n5 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_17/n6 ), .CK(CLK), .QN(
        \unit_control/uut_third_stage/ffi_17/n5 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_19/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_15/n5 ), .CK(CLK), .Q(n1913), .QN(
        \unit_control/uut_third_stage/ffi_19/n5 ) );
  SNPS_CLOCK_GATE_HIGH_dlx_0 \clk_gate_unit_decode/NPC1reg/ffi_31/Q_reg  ( 
        .CLK(CLK), .EN(n2932), .ENCLK(n3087), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dlx_1 \clk_gate_unit_execution/COMP_NPC2/ffi_31/Q_reg  ( 
        .CLK(CLK), .EN(n471), .ENCLK(n3004), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dlx_3 \clk_gate_unit_fetch/unit_programCounter/ffi_9/Q_reg  ( 
        .CLK(CLK), .EN(n1923), .ENCLK(n2933), .TE(1'b0) );
  DFF_X2 \unit_decode/IMMreg/ffi_3/Q_reg  ( .D(n3012), .CK(n3087), .Q(n1662), 
        .QN(\unit_decode/IMMreg/ffi_3/n4 ) );
  DFF_X2 \unit_decode/IMMreg/ffi_31/Q_reg  ( .D(n2934), .CK(n3087), .Q(n1660), 
        .QN(\unit_decode/IMMreg/ffi_31/n4 ) );
  DFF_X2 \unit_decode/IMMreg/ffi_0/Q_reg  ( .D(n3010), .CK(n3087), .Q(n1653), 
        .QN(\unit_decode/IMMreg/ffi_0/n4 ) );
  DFF_X1 \unit_execution/COMP_REGN_ALUOUT/ffi_1/Q_reg  ( .D(n2941), .CK(n3004), 
        .QN(\unit_execution/COMP_REGN_ALUOUT/ffi_1/n4 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[17]  ( .D(
        \unit_fetch/unit_instructionRegister/n81 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n55 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[22]  ( .D(
        \unit_fetch/unit_instructionRegister/n78 ), .CK(CLK), .Q(
        \unit_decode/RS1s[1] ), .QN(\unit_fetch/unit_instructionRegister/n60 )
         );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U69  ( .A(n1642), .B(
        \unit_fetch/unit_programCounter/ffi_10/n4 ), .ZN(
        \unit_fetch/adder_out[10] ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U13  ( .A(
        \unit_fetch/unit_adder/add_19/n14 ), .B(
        \unit_fetch/unit_programCounter/ffi_20/n4 ), .ZN(
        \unit_fetch/adder_out[20] ) );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U18  ( .A1(n1641), .A2(
        \unit_fetch/unit_adder/add_19/n15 ), .ZN(
        \unit_fetch/unit_adder/add_19/n14 ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U89  ( .A(
        \unit_fetch/unit_adder/add_19/n77 ), .B(
        \unit_fetch/unit_programCounter/ffi_6/n4 ), .Z(
        \unit_fetch/adder_out[6] ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U104  ( .A(
        \unit_fetch/unit_programCounter/ffi_3/n4 ), .B(n1603), .ZN(
        \unit_fetch/adder_out[3] ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U94  ( .A(
        \unit_fetch/unit_adder/add_19/n82 ), .B(
        \unit_fetch/unit_adder/add_19/n81 ), .Z(\unit_fetch/adder_out[5] ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U101  ( .A1(
        \unit_fetch/unit_adder/add_19/n85 ), .A2(\unit_fetch/pc_regout[4] ), 
        .ZN(\unit_fetch/unit_adder/add_19/n82 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U100  ( .A(
        \unit_fetch/unit_adder/add_19/n84 ), .B(
        \unit_fetch/unit_adder/add_19/n85 ), .ZN(\unit_fetch/adder_out[4] ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U84  ( .A(
        \unit_fetch/unit_adder/add_19/n73 ), .B(
        \unit_fetch/unit_programCounter/ffi_7/n4 ), .ZN(
        \unit_fetch/adder_out[7] ) );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U90  ( .A1(
        \unit_fetch/unit_adder/add_19/n77 ), .A2(
        \unit_fetch/unit_programCounter/ffi_6/n4 ), .ZN(
        \unit_fetch/unit_adder/add_19/n73 ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U63  ( .A(
        \unit_fetch/unit_adder/add_19/n57 ), .B(
        \unit_fetch/unit_programCounter/ffi_11/n4 ), .Z(
        \unit_fetch/adder_out[11] ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U70  ( .A1(n1642), .A2(
        \unit_fetch/pc_regout[10] ), .ZN(\unit_fetch/unit_adder/add_19/n57 )
         );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U73  ( .A(
        \unit_fetch/unit_adder/add_19/n66 ), .B(
        \unit_fetch/unit_programCounter/ffi_9/n4 ), .Z(
        \unit_fetch/adder_out[9] ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U81  ( .A1(
        \unit_fetch/unit_adder/add_19/n69 ), .A2(\unit_fetch/pc_regout[8] ), 
        .ZN(\unit_fetch/unit_adder/add_19/n66 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U51  ( .A(
        \unit_fetch/unit_adder/add_19/n48 ), .B(
        \unit_fetch/unit_adder/add_19/n47 ), .ZN(\unit_fetch/adder_out[13] )
         );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U59  ( .A1(
        \unit_fetch/unit_adder/add_19/n52 ), .A2(
        \unit_fetch/unit_programCounter/ffi_12/n4 ), .ZN(
        \unit_fetch/unit_adder/add_19/n48 ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U22  ( .A(n1641), .B(
        \unit_fetch/unit_programCounter/ffi_18/n4 ), .Z(
        \unit_fetch/adder_out[18] ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U27  ( .A(
        \unit_fetch/unit_adder/add_19/n29 ), .B(
        \unit_fetch/unit_adder/add_19/n28 ), .ZN(\unit_fetch/adder_out[17] )
         );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U36  ( .A1(
        \unit_fetch/unit_adder/add_19/n33 ), .A2(
        \unit_fetch/unit_adder/add_19/n32 ), .ZN(
        \unit_fetch/unit_adder/add_19/n29 ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U35  ( .A(
        \unit_fetch/unit_adder/add_19/n33 ), .B(
        \unit_fetch/unit_adder/add_19/n32 ), .Z(\unit_fetch/adder_out[16] ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U41  ( .A1(
        \unit_fetch/unit_adder/add_19/n42 ), .A2(
        \unit_fetch/unit_adder/add_19/n34 ), .ZN(
        \unit_fetch/unit_adder/add_19/n33 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U40  ( .A(
        \unit_fetch/unit_adder/add_19/n38 ), .B(
        \unit_fetch/unit_adder/add_19/n37 ), .ZN(\unit_fetch/adder_out[15] )
         );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U47  ( .A1(
        \unit_fetch/unit_adder/add_19/n43 ), .A2(
        \unit_fetch/unit_adder/add_19/n41 ), .ZN(
        \unit_fetch/unit_adder/add_19/n38 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U46  ( .A(
        \unit_fetch/unit_adder/add_19/n42 ), .B(
        \unit_fetch/unit_adder/add_19/n41 ), .ZN(\unit_fetch/adder_out[14] )
         );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U53  ( .A1(n1642), .A2(
        \unit_fetch/unit_adder/add_19/n44 ), .ZN(
        \unit_fetch/unit_adder/add_19/n43 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U80  ( .A(
        \unit_fetch/unit_adder/add_19/n69 ), .B(
        \unit_fetch/unit_programCounter/ffi_8/n4 ), .ZN(
        \unit_fetch/adder_out[8] ) );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U85  ( .A1(
        \unit_fetch/unit_adder/add_19/n77 ), .A2(
        \unit_fetch/unit_adder/add_19/n70 ), .ZN(
        \unit_fetch/unit_adder/add_19/n69 ) );
  XOR2_X1 \unit_fetch/unit_adder/add_19/U58  ( .A(
        \unit_fetch/unit_adder/add_19/n52 ), .B(
        \unit_fetch/unit_programCounter/ffi_12/n4 ), .Z(
        \unit_fetch/adder_out[12] ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U64  ( .A1(n1642), .A2(
        \unit_fetch/unit_adder/add_19/n53 ), .ZN(
        \unit_fetch/unit_adder/add_19/n52 ) );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U15  ( .A1(
        \unit_fetch/unit_adder/add_19/n15 ), .A2(
        \unit_fetch/unit_programCounter/ffi_20/n4 ), .ZN(
        \unit_fetch/unit_adder/add_19/n12 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U19  ( .A1(\unit_fetch/pc_regout[18] ), .A2(\unit_fetch/pc_regout[19] ), .ZN(\unit_fetch/unit_adder/add_19/n15 ) );
  XNOR2_X1 \unit_fetch/unit_adder/add_19/U17  ( .A(
        \unit_fetch/unit_adder/add_19/n18 ), .B(
        \unit_fetch/unit_adder/add_19/n17 ), .ZN(\unit_fetch/adder_out[19] )
         );
  NOR2_X1 \unit_fetch/unit_adder/add_19/U23  ( .A1(n1641), .A2(
        \unit_fetch/unit_programCounter/ffi_18/n4 ), .ZN(
        \unit_fetch/unit_adder/add_19/n18 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U55  ( .A1(\unit_fetch/pc_regout[12] ), .A2(\unit_fetch/pc_regout[13] ), .ZN(\unit_fetch/unit_adder/add_19/n45 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U97  ( .A1(\unit_fetch/pc_regout[4] ), 
        .A2(\unit_fetch/pc_regout[5] ), .ZN(\unit_fetch/unit_adder/add_19/n79 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U43  ( .A1(\unit_fetch/pc_regout[14] ), .A2(\unit_fetch/pc_regout[15] ), .ZN(\unit_fetch/unit_adder/add_19/n35 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U86  ( .A1(\unit_fetch/pc_regout[6] ), 
        .A2(\unit_fetch/pc_regout[7] ), .ZN(\unit_fetch/unit_adder/add_19/n70 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U77  ( .A1(\unit_fetch/pc_regout[8] ), 
        .A2(\unit_fetch/pc_regout[9] ), .ZN(\unit_fetch/unit_adder/add_19/n63 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U106  ( .A1(\unit_fetch/pc_regout[3] ), .A2(\unit_fetch/pc_regout[2] ), .ZN(\unit_fetch/unit_adder/add_19/n86 ) );
  NAND2_X1 \unit_fetch/unit_adder/add_19/U66  ( .A1(\unit_fetch/pc_regout[10] ), .A2(\unit_fetch/pc_regout[11] ), .ZN(\unit_fetch/unit_adder/add_19/n54 ) );
  HA_X1 \unit_fetch/unit_adder/add_19/U9  ( .A(
        \unit_fetch/unit_adder/add_19/n9 ), .B(\unit_fetch/pc_regout[23] ), 
        .CO(\unit_fetch/unit_adder/add_19/n8 ), .S(\unit_fetch/adder_out[23] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U8  ( .A(
        \unit_fetch/unit_adder/add_19/n8 ), .B(\unit_fetch/pc_regout[24] ), 
        .CO(\unit_fetch/unit_adder/add_19/n7 ), .S(\unit_fetch/adder_out[24] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U7  ( .A(
        \unit_fetch/unit_adder/add_19/n7 ), .B(\unit_fetch/pc_regout[25] ), 
        .CO(\unit_fetch/unit_adder/add_19/n6 ), .S(\unit_fetch/adder_out[25] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U6  ( .A(
        \unit_fetch/unit_adder/add_19/n6 ), .B(\unit_fetch/pc_regout[26] ), 
        .CO(\unit_fetch/unit_adder/add_19/n5 ), .S(\unit_fetch/adder_out[26] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U5  ( .A(
        \unit_fetch/unit_adder/add_19/n5 ), .B(\unit_fetch/pc_regout[27] ), 
        .CO(\unit_fetch/unit_adder/add_19/n4 ), .S(\unit_fetch/adder_out[27] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U4  ( .A(
        \unit_fetch/unit_adder/add_19/n4 ), .B(\unit_fetch/pc_regout[28] ), 
        .CO(\unit_fetch/unit_adder/add_19/n3 ), .S(\unit_fetch/adder_out[28] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U3  ( .A(
        \unit_fetch/unit_adder/add_19/n3 ), .B(\unit_fetch/pc_regout[29] ), 
        .CO(\unit_fetch/unit_adder/add_19/n2 ), .S(\unit_fetch/adder_out[29] )
         );
  HA_X1 \unit_fetch/unit_adder/add_19/U2  ( .A(
        \unit_fetch/unit_adder/add_19/n2 ), .B(\unit_fetch/pc_regout[30] ), 
        .CO(\unit_fetch/unit_adder/add_19/n1 ), .S(\unit_fetch/adder_out[30] )
         );
  DFF_X1 \unit_decode/Areg/ffi_19/Q_reg  ( .D(n3042), .CK(n3087), .Q(n1645) );
  DFF_X1 \unit_decode/Areg/ffi_8/Q_reg  ( .D(n3031), .CK(n3087), .Q(n1647) );
  DFF_X1 \unit_decode/IMMreg/ffi_10/Q_reg  ( .D(n3018), .CK(n3087), .Q(n1667)
         );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_0/Q_reg  ( .D(n2935), .CK(n3004), 
        .Q(wr_address[0]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_2/Q_reg  ( .D(n2937), .CK(n3004), 
        .Q(wr_address[2]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_4/Q_reg  ( .D(n2939), .CK(n3004), 
        .Q(wr_address[4]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_4/n5 ), .CK(CLK), .Q(
        \unit_control/cw2delay[4] ) );
  DFF_X1 \unit_control/uut_fourth_stage/ffi_4/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_4/n5 ), .CK(CLK), .Q(\cw_mem[4] )
         );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_3/Q_reg  ( .D(n2938), .CK(n3004), 
        .Q(wr_address[3]) );
  DFF_X1 \unit_execution/COMP_REG5_RD2OUT/ffi_1/Q_reg  ( .D(n2936), .CK(n3004), 
        .Q(wr_address[1]) );
  DFF_X1 \unit_control/uut_third_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_3/n5 ), .CK(CLK), .Q(
        \unit_control/cw2delay[3] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_12/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[12] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_14/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_14/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[14] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_9/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_24/n3 ), .CK(CLK), .Q(
        \unit_control/cw1delay[9] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_13/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[13] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_3/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[3] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_10/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[10] ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_17/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_17/n5 ), .CK(CLK), .Q(
        \unit_control/cw1delay[17] ) );
  DFFRS_X1 \unit_control/uut_second_stage/ffi_4/Q_reg  ( .D(n4), .CK(CLK), 
        .RN(1'b1), .SN(1'b1), .Q(\unit_control/cw1delay[4] ) );
  DFFRS_X1 \unit_fetch/unit_npcregister/ffi_29/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_29/n5 ), .CK(n2933), .RN(1'b1), .SN(
        1'b1), .QN(\unit_fetch/unit_npcregister/ffi_29/n4 ) );
  DFFRS_X1 \unit_fetch/unit_npcregister/ffi_19/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_19/n5 ), .CK(n2933), .RN(1'b1), .SN(
        1'b1), .QN(\unit_fetch/unit_npcregister/ffi_19/n4 ) );
  SDFFS_X1 \unit_decode/IMMreg/ffi_2/Q_reg  ( .D(n3011), .SI(1'b0), .SE(1'b0), 
        .CK(n3087), .SN(1'b1), .Q(n1665), .QN(\unit_decode/IMMreg/ffi_2/n4 )
         );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_13/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_13/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[13] ), .QN(\unit_fetch/unit_adder/add_19/n47 )
         );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_31/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_31/n5 ), .CK(n2933), .QN(n1606) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_0/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_0/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[0] ), .QN(
        \unit_fetch/unit_programCounter/ffi_0/n4 ) );
  DFFRS_X1 \unit_fetch/unit_npcregister/ffi_31/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_31/n5 ), .CK(n2933), .RN(1'b1), .SN(
        1'b1), .QN(\unit_fetch/unit_npcregister/ffi_31/n4 ) );
  DFF_X1 \unit_control/uut_second_stage/ffi_15/Q_reg  ( .D(n6), .CK(CLK), .QN(
        n1340) );
  DFF_X1 \unit_control/uut_second_stage/ffi_21/Q_reg  ( .D(
        \unit_control/uut_second_stage/ffi_21/n5 ), .CK(CLK), .Q(n1687), .QN(
        n1330) );
  DFF_X1 \unit_decode/IMMreg/ffi_25/Q_reg  ( .D(\unit_decode/IMMreg/ffi_25/n5 ), .CK(CLK), .Q(n1689), .QN(\unit_decode/IMMreg/ffi_25/n4 ) );
  DFF_X1 \unit_control/uut_third_stage/ffi_14/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_14/n5 ), .CK(CLK), .Q(n1673), .QN(
        n1336) );
  DFF_X1 \unit_control/uut_third_stage/ffi_13/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_13/n5 ), .CK(CLK), .Q(n1671), .QN(
        n1341) );
  DFF_X1 \unit_control/uut_third_stage/ffi_12/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_12/n5 ), .CK(CLK), .Q(n1655), .QN(
        n1338) );
  DFF_X1 \unit_control/uut_third_stage/ffi_10/Q_reg  ( .D(
        \unit_control/uut_third_stage/ffi_10/n5 ), .CK(CLK), .Q(n1661), .QN(
        n1342) );
  DFF_X1 \unit_control/uut_second_stage/ffi_22/Q_reg  ( .D(n1942), .CK(CLK), 
        .Q(\cw_dec[2] ), .QN(n1337) );
  DFFRS_X1 \unit_fetch/unit_npcregister/ffi_28/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_28/n5 ), .CK(n2933), .RN(1'b1), .SN(
        1'b1), .QN(\unit_fetch/unit_npcregister/ffi_28/n4 ) );
  SDFF_X1 \unit_decode/IMMreg/ffi_1/Q_reg  ( .D(1'b1), .SI(
        \unit_fetch/unit_instructionRegister/n39 ), .SE(n1942), .CK(n3087), 
        .Q(n1612), .QN(n1664) );
  DFF_X2 \unit_control/uut_fourth_stage/ffi_3/Q_reg  ( .D(
        \unit_control/uut_fourth_stage/ffi_3/n6 ), .CK(CLK), .Q(n1685), .QN(
        n1650) );
  DFF_X1 \unit_fetch/unit_programCounter/ffi_2/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_2/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[2] ), .QN(
        \unit_fetch/unit_programCounter/ffi_2/n4 ) );
  DFF_X1 \unit_fetch/unit_instructionRegister/regOut_reg[9]  ( .D(
        \unit_fetch/unit_instructionRegister/n89 ), .CK(CLK), .QN(
        \unit_fetch/unit_instructionRegister/n47 ) );
  DFF_X2 \unit_fetch/unit_programCounter/ffi_6/Q_reg  ( .D(
        \unit_fetch/unit_programCounter/ffi_6/n5 ), .CK(n2933), .Q(
        \unit_fetch/pc_regout[6] ), .QN(
        \unit_fetch/unit_programCounter/ffi_6/n4 ) );
  DFFRS_X1 \unit_fetch/unit_npcregister/ffi_0/Q_reg  ( .D(
        \unit_fetch/unit_npcregister/ffi_0/n5 ), .CK(n2933), .RN(1'b1), .SN(
        1'b1), .QN(\unit_fetch/unit_npcregister/ffi_0/n4 ) );
  OAI33_X1 U1731 ( .A1(1'b0), .A2(\unit_decode/IMMreg/ffi_2/n4 ), .A3(n1493), 
        .B1(n1494), .B2(n2607), .B3(n2611), .ZN(n1496) );
  OAI33_X1 U1732 ( .A1(1'b0), .A2(n1472), .A3(n1473), .B1(n1628), .B2(n2779), 
        .B3(n1567), .ZN(n1475) );
  OAI33_X1 U1733 ( .A1(1'b0), .A2(n1449), .A3(n1450), .B1(n1633), .B2(n2779), 
        .B3(\unit_decode/IMMreg/ffi_5/n4 ), .ZN(n1452) );
  OAI33_X1 U1734 ( .A1(1'b0), .A2(n2510), .A3(n1416), .B1(n1417), .B2(
        \unit_decode/IMMreg/ffi_11/n4 ), .B3(n2779), .ZN(n1419) );
  BUF_X1 U1735 ( .A(n2417), .Z(n1344) );
  XNOR2_X1 U1736 ( .A(n2150), .B(n1345), .ZN(n1360) );
  XNOR2_X1 U1737 ( .A(n1530), .B(n1612), .ZN(n1345) );
  BUF_X2 U1738 ( .A(n1344), .Z(n1346) );
  NAND2_X1 U1739 ( .A1(n2010), .A2(n2564), .ZN(n1547) );
  NAND2_X1 U1740 ( .A1(n2574), .A2(n2562), .ZN(n2564) );
  INV_X1 U1741 ( .A(n2103), .ZN(n1347) );
  INV_X1 U1742 ( .A(n1387), .ZN(n1348) );
  BUF_X1 U1743 ( .A(\unit_fetch/unit_adder/add_19/n89 ), .Z(n1349) );
  INV_X1 U1744 ( .A(n2135), .ZN(n1350) );
  INV_X1 U1745 ( .A(n1358), .ZN(n1351) );
  BUF_X1 U1746 ( .A(n1547), .Z(n1352) );
  NAND2_X1 U1747 ( .A1(n2639), .A2(n1374), .ZN(n1816) );
  XNOR2_X1 U1748 ( .A(n1442), .B(n1907), .ZN(n1374) );
  NOR2_X1 U1749 ( .A1(n1547), .A2(n2051), .ZN(n2045) );
  AOI21_X1 U1750 ( .B1(n1714), .B2(n1715), .A(n1353), .ZN(n2625) );
  NAND2_X1 U1751 ( .A1(n1764), .A2(n1765), .ZN(n1353) );
  NAND2_X1 U1752 ( .A1(n2424), .A2(n1766), .ZN(n1764) );
  NAND2_X1 U1753 ( .A1(n1395), .A2(n2484), .ZN(n2424) );
  INV_X2 U1754 ( .A(n1987), .ZN(n1986) );
  NAND2_X1 U1755 ( .A1(n1356), .A2(n1354), .ZN(n1598) );
  AND3_X2 U1756 ( .A1(n2008), .A2(n1980), .A3(n1355), .ZN(n1354) );
  OR2_X2 U1757 ( .A1(n2154), .A2(n1538), .ZN(n1355) );
  NAND2_X1 U1758 ( .A1(n2154), .A2(n1538), .ZN(n1980) );
  NAND2_X1 U1759 ( .A1(n2147), .A2(n1988), .ZN(n2008) );
  NAND2_X1 U1760 ( .A1(n1359), .A2(n1987), .ZN(n1356) );
  NAND2_X1 U1761 ( .A1(n1358), .A2(n1357), .ZN(n1987) );
  INV_X1 U1762 ( .A(n1967), .ZN(n1357) );
  INV_X1 U1763 ( .A(n2150), .ZN(n1358) );
  NAND2_X1 U1764 ( .A1(n1360), .A2(n1969), .ZN(n1359) );
  AND2_X1 U1765 ( .A1(n1529), .A2(n1968), .ZN(n1969) );
  BUF_X1 U1766 ( .A(n2643), .Z(n1361) );
  BUF_X1 U1767 ( .A(n1632), .Z(n1362) );
  XOR2_X1 U1768 ( .A(n2451), .B(n2199), .Z(n1632) );
  INV_X1 U1769 ( .A(n2211), .ZN(n1363) );
  XNOR2_X1 U1770 ( .A(\unit_decode/IMMreg/ffi_31/n4 ), .B(n1937), .ZN(n2210)
         );
  NOR2_X1 U1771 ( .A1(n1816), .A2(n2640), .ZN(n1364) );
  BUF_X1 U1772 ( .A(n2880), .Z(n1365) );
  OAI211_X1 U1773 ( .C1(n1886), .C2(\unit_control/n152 ), .A(n1799), .B(n1798), 
        .ZN(n1366) );
  OAI211_X1 U1774 ( .C1(n1886), .C2(\unit_control/n152 ), .A(n1799), .B(n1798), 
        .ZN(n1367) );
  NOR2_X2 U1775 ( .A1(n1887), .A2(n2740), .ZN(n1886) );
  NAND3_X1 U1776 ( .A1(n2195), .A2(n1828), .A3(n2484), .ZN(n1368) );
  INV_X1 U1777 ( .A(n2473), .ZN(n1369) );
  INV_X1 U1778 ( .A(n2286), .ZN(n1370) );
  NOR2_X1 U1779 ( .A1(n2303), .A2(n2302), .ZN(n2352) );
  AND2_X1 U1780 ( .A1(n1367), .A2(n1942), .ZN(n1559) );
  BUF_X1 U1781 ( .A(n2644), .Z(n1371) );
  INV_X1 U1782 ( .A(n1480), .ZN(n1372) );
  BUF_X1 U1783 ( .A(n1608), .Z(n1373) );
  INV_X1 U1784 ( .A(n2371), .ZN(n1375) );
  NAND2_X2 U1785 ( .A1(n2174), .A2(n1652), .ZN(n2120) );
  NOR2_X2 U1786 ( .A1(n1945), .A2(n2587), .ZN(n2174) );
  OR2_X1 U1787 ( .A1(\unit_fetch/unit_programCounter/ffi_16/n4 ), .A2(n1923), 
        .ZN(n1376) );
  NAND2_X1 U1788 ( .A1(n2671), .A2(n1376), .ZN(
        \unit_fetch/unit_programCounter/ffi_16/n5 ) );
  INV_X2 U1789 ( .A(n1925), .ZN(n1923) );
  BUF_X1 U1790 ( .A(n1879), .Z(n1377) );
  INV_X1 U1791 ( .A(n1736), .ZN(n1378) );
  NOR2_X2 U1792 ( .A1(n2488), .A2(n2196), .ZN(n2423) );
  AND2_X1 U1793 ( .A1(n1840), .A2(n1839), .ZN(n1569) );
  XNOR2_X1 U1794 ( .A(n2210), .B(n1797), .ZN(n1379) );
  INV_X2 U1795 ( .A(n1925), .ZN(n1924) );
  NOR2_X1 U1796 ( .A1(n1380), .A2(n1599), .ZN(n1813) );
  NAND2_X1 U1797 ( .A1(n1814), .A2(n2437), .ZN(n1380) );
  INV_X1 U1798 ( .A(n1455), .ZN(n1381) );
  AND2_X2 U1799 ( .A1(n2389), .A2(n2367), .ZN(n1382) );
  INV_X2 U1800 ( .A(n1382), .ZN(n2415) );
  AND2_X1 U1801 ( .A1(n1609), .A2(n1762), .ZN(n2414) );
  INV_X1 U1802 ( .A(n1385), .ZN(n1383) );
  AND2_X1 U1803 ( .A1(n1902), .A2(n2054), .ZN(n1384) );
  BUF_X1 U1804 ( .A(n1757), .Z(n1385) );
  INV_X1 U1805 ( .A(n2057), .ZN(n1386) );
  INV_X1 U1806 ( .A(n2158), .ZN(n1387) );
  INV_X1 U1807 ( .A(n2767), .ZN(n1388) );
  AOI221_X1 U1808 ( .B1(n1580), .B2(n2779), .C1(n2767), .C2(n2778), .A(
        \unit_decode/IMMreg/ffi_16/n4 ), .ZN(n2768) );
  BUF_X1 U1809 ( .A(n2624), .Z(n1389) );
  INV_X1 U1810 ( .A(n1664), .ZN(n1390) );
  BUF_X1 U1811 ( .A(n2623), .Z(n1391) );
  AOI21_X1 U1812 ( .B1(n1501), .B2(n2052), .A(n1500), .ZN(n1392) );
  AND2_X1 U1813 ( .A1(n1387), .A2(n2053), .ZN(n1393) );
  BUF_X1 U1814 ( .A(n1834), .Z(n1394) );
  XNOR2_X1 U1815 ( .A(n1938), .B(n1668), .ZN(n2197) );
  OAI21_X1 U1816 ( .B1(n1531), .B2(n2190), .A(n1830), .ZN(n1395) );
  OAI21_X1 U1817 ( .B1(n1531), .B2(n2190), .A(n1830), .ZN(n2195) );
  BUF_X1 U1818 ( .A(n2520), .Z(n1396) );
  CLKBUF_X3 U1819 ( .A(\unit_control/uut_third_stage/ffi_19/n5 ), .Z(n1934) );
  OAI21_X1 U1820 ( .B1(n1624), .B2(n1653), .A(n1528), .ZN(n2626) );
  BUF_X1 U1821 ( .A(n1529), .Z(n1528) );
  CLKBUF_X3 U1822 ( .A(n1915), .Z(n1941) );
  NOR2_X1 U1823 ( .A1(n2208), .A2(n2209), .ZN(n1881) );
  BUF_X1 U1824 ( .A(n2290), .Z(n1582) );
  OAI21_X1 U1825 ( .B1(n2079), .B2(n2502), .A(n2188), .ZN(n2111) );
  BUF_X1 U1826 ( .A(n1348), .Z(n1544) );
  OAI21_X1 U1827 ( .B1(n2608), .B2(n2609), .A(n1516), .ZN(n2616) );
  INV_X1 U1828 ( .A(n1537), .ZN(n2349) );
  INV_X1 U1829 ( .A(n1535), .ZN(n2404) );
  BUF_X1 U1830 ( .A(n2711), .Z(n1580) );
  BUF_X1 U1831 ( .A(n2542), .Z(n1589) );
  BUF_X1 U1832 ( .A(n2229), .Z(n1618) );
  AOI211_X1 U1833 ( .C1(n2845), .C2(n2889), .A(n2898), .B(n2871), .ZN(n2850)
         );
  NAND2_X1 U1834 ( .A1(n1383), .A2(\unit_decode/Areg/ffi_14/n4 ), .ZN(n1397)
         );
  OAI21_X1 U1835 ( .B1(n1514), .B2(n1935), .A(n1397), .ZN(n2228) );
  NOR4_X1 U1836 ( .A1(n2629), .A2(n2628), .A3(n2627), .A4(n2626), .ZN(n1398)
         );
  NAND4_X1 U1837 ( .A1(n1398), .A2(n2631), .A3(n2632), .A4(n2630), .ZN(n2634)
         );
  OAI22_X1 U1838 ( .A1(n2488), .A2(n2248), .B1(n2374), .B2(n1918), .ZN(n1399)
         );
  AOI21_X1 U1839 ( .B1(n1544), .B2(n2252), .A(n1399), .ZN(n1400) );
  NAND2_X1 U1840 ( .A1(n2288), .A2(n1575), .ZN(n1401) );
  NAND3_X1 U1841 ( .A1(n1401), .A2(n1400), .A3(n2294), .ZN(n2320) );
  AOI21_X1 U1842 ( .B1(n2756), .B2(n1845), .A(n2780), .ZN(n1402) );
  OAI211_X1 U1843 ( .C1(n2514), .C2(n2608), .A(n1844), .B(n2101), .ZN(n1403)
         );
  OAI21_X1 U1844 ( .B1(n2529), .B2(n2449), .A(n1843), .ZN(n1404) );
  NOR3_X1 U1845 ( .A1(n1402), .A2(n1403), .A3(n1404), .ZN(n1405) );
  OAI21_X1 U1846 ( .B1(n1651), .B2(n2544), .A(n1405), .ZN(n2913) );
  OAI221_X1 U1847 ( .B1(n1881), .B2(n2303), .C1(n1881), .C2(n2304), .A(n1379), 
        .ZN(n1406) );
  INV_X1 U1848 ( .A(n1696), .ZN(n1407) );
  NAND2_X1 U1849 ( .A1(n1406), .A2(n1407), .ZN(n1581) );
  NAND2_X1 U1850 ( .A1(n2750), .A2(n2612), .ZN(n1408) );
  INV_X1 U1851 ( .A(n1986), .ZN(n1409) );
  OAI221_X1 U1852 ( .B1(n1978), .B2(n1979), .C1(n1978), .C2(n1408), .A(n1409), 
        .ZN(n1981) );
  OAI22_X1 U1853 ( .A1(n2388), .A2(n1918), .B1(n1554), .B2(n2248), .ZN(n1410)
         );
  AOI21_X1 U1854 ( .B1(n1618), .B2(n2252), .A(n1410), .ZN(n1411) );
  NAND2_X1 U1855 ( .A1(n2288), .A2(n2230), .ZN(n1412) );
  NAND3_X1 U1856 ( .A1(n1412), .A2(n1411), .A3(n2294), .ZN(n2334) );
  NAND2_X1 U1857 ( .A1(n2593), .A2(n2504), .ZN(n1413) );
  NAND4_X1 U1858 ( .A1(n1725), .A2(n1726), .A3(n2509), .A4(n1413), .ZN(n1414)
         );
  INV_X1 U1859 ( .A(\unit_decode/IMMreg/ffi_11/n4 ), .ZN(n1415) );
  AOI22_X1 U1860 ( .A1(\unit_decode/IMMreg/ffi_11/n4 ), .A2(n2541), .B1(n2573), 
        .B2(n1415), .ZN(n1416) );
  INV_X1 U1861 ( .A(n2510), .ZN(n1417) );
  AOI21_X1 U1863 ( .B1(n2622), .B2(n1414), .A(n1419), .ZN(n1420) );
  OAI21_X1 U1864 ( .B1(n2544), .B2(n2638), .A(n1420), .ZN(n2703) );
  INV_X1 U1865 ( .A(n2288), .ZN(n1421) );
  OAI22_X1 U1866 ( .A1(n2773), .A2(n1589), .B1(n2291), .B2(n1624), .ZN(n1422)
         );
  AOI21_X1 U1867 ( .B1(n2711), .B2(n2175), .A(n1422), .ZN(n1423) );
  OAI211_X1 U1868 ( .C1(n2353), .C2(n1421), .A(n2294), .B(n1423), .ZN(n2442)
         );
  NOR4_X1 U1869 ( .A1(n2519), .A2(n2518), .A3(n2516), .A4(n2517), .ZN(n1424)
         );
  INV_X1 U1870 ( .A(n2522), .ZN(n1425) );
  INV_X1 U1871 ( .A(n1667), .ZN(n1426) );
  AOI22_X1 U1872 ( .A1(n1667), .A2(n2778), .B1(n2611), .B2(n1426), .ZN(n1427)
         );
  OAI222_X1 U1873 ( .A1(n1425), .A2(n1667), .B1(n1425), .B2(n2570), .C1(n2522), 
        .C2(n1427), .ZN(n1428) );
  NAND2_X1 U1874 ( .A1(n2633), .A2(n2617), .ZN(n1429) );
  OAI211_X1 U1875 ( .C1(n1424), .C2(n2780), .A(n1428), .B(n1429), .ZN(n2704)
         );
  OAI22_X1 U1876 ( .A1(n1918), .A2(n2267), .B1(n2248), .B2(n1629), .ZN(n1430)
         );
  OAI22_X1 U1877 ( .A1(n2291), .A2(n1626), .B1(n2171), .B2(n1633), .ZN(n1431)
         );
  NOR3_X1 U1878 ( .A1(n2174), .A2(n1430), .A3(n1431), .ZN(n2257) );
  OAI22_X1 U1879 ( .A1(n2611), .A2(n1670), .B1(\unit_decode/IMMreg/ffi_24/n4 ), 
        .B2(n2778), .ZN(n1432) );
  NOR3_X1 U1880 ( .A1(n2353), .A2(\unit_decode/IMMreg/ffi_24/n4 ), .A3(n2779), 
        .ZN(n1433) );
  AOI21_X1 U1881 ( .B1(n2353), .B2(n1432), .A(n1433), .ZN(n2354) );
  AOI21_X1 U1882 ( .B1(n1540), .B2(n1713), .A(n2446), .ZN(n1434) );
  MUX2_X1 U1883 ( .A(n1434), .B(n2447), .S(n1362), .Z(n2640) );
  INV_X1 U1884 ( .A(n2777), .ZN(n1435) );
  INV_X1 U1885 ( .A(n2757), .ZN(n1436) );
  AOI222_X1 U1886 ( .A1(n1435), .A2(n1436), .B1(n2465), .B2(n2593), .C1(n2406), 
        .C2(n2772), .ZN(n1845) );
  NOR3_X1 U1887 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_8/n4 ), .A3(n1589), 
        .ZN(n1437) );
  AOI21_X1 U1888 ( .B1(n1589), .B2(n2543), .A(n1437), .ZN(n1438) );
  NAND3_X1 U1889 ( .A1(n2538), .A2(n2539), .A3(n2540), .ZN(n1439) );
  NAND2_X1 U1890 ( .A1(n1439), .A2(n2622), .ZN(n1440) );
  OAI211_X1 U1891 ( .C1(n2630), .C2(n2544), .A(n1438), .B(n1440), .ZN(n2705)
         );
  AOI21_X1 U1892 ( .B1(n2209), .B2(n2208), .A(n1881), .ZN(n2304) );
  AND3_X1 U1893 ( .A1(n1609), .A2(n1879), .A3(n1784), .ZN(n1441) );
  NOR2_X1 U1894 ( .A1(n1441), .A2(n1551), .ZN(n1442) );
  NAND2_X1 U1895 ( .A1(n2571), .A2(n1643), .ZN(n1443) );
  AOI22_X1 U1896 ( .A1(n2175), .A2(n2510), .B1(n1619), .B2(n2775), .ZN(n1444)
         );
  NAND3_X1 U1897 ( .A1(n1443), .A2(n1444), .A3(n2120), .ZN(n2465) );
  AOI22_X1 U1898 ( .A1(n2537), .A2(n2596), .B1(n2027), .B2(n2535), .ZN(n1445)
         );
  AOI21_X1 U1899 ( .B1(n2772), .B2(n2508), .A(n1998), .ZN(n1446) );
  NAND3_X1 U1900 ( .A1(n1445), .A2(n1999), .A3(n1446), .ZN(n1447) );
  INV_X1 U1901 ( .A(n1680), .ZN(n1448) );
  AOI22_X1 U1902 ( .A1(n1680), .A2(n2573), .B1(n2541), .B2(n1448), .ZN(n1449)
         );
  INV_X1 U1903 ( .A(n1633), .ZN(n1450) );
  AOI21_X1 U1905 ( .B1(n2622), .B2(n1447), .A(n1452), .ZN(n1453) );
  OAI21_X1 U1906 ( .B1(n2632), .B2(n2544), .A(n1453), .ZN(n2917) );
  NAND4_X1 U1907 ( .A1(n1840), .A2(n1382), .A3(n1701), .A4(n1839), .ZN(n1454)
         );
  INV_X1 U1908 ( .A(n2368), .ZN(n1455) );
  AOI21_X1 U1909 ( .B1(n1454), .B2(n1455), .A(n1907), .ZN(n1906) );
  OAI21_X1 U1910 ( .B1(n1776), .B2(n1775), .A(n1777), .ZN(n1456) );
  NAND3_X1 U1911 ( .A1(n2198), .A2(n1779), .A3(n1778), .ZN(n1457) );
  NAND2_X1 U1912 ( .A1(n1457), .A2(n1456), .ZN(n2473) );
  NOR3_X1 U1913 ( .A1(\unit_fetch/unit_adder/add_19/n79 ), .A2(
        \unit_fetch/unit_adder/add_19/n45 ), .A3(
        \unit_fetch/unit_adder/add_19/n35 ), .ZN(n1458) );
  NAND3_X1 U1914 ( .A1(\unit_fetch/pc_regout[17] ), .A2(
        \unit_fetch/pc_regout[16] ), .A3(n1458), .ZN(n1640) );
  INV_X1 U1915 ( .A(n2302), .ZN(n1459) );
  AOI21_X1 U1916 ( .B1(n2301), .B2(n1459), .A(n2303), .ZN(n1460) );
  NOR2_X1 U1917 ( .A1(n2333), .A2(n1460), .ZN(n1461) );
  NOR2_X1 U1918 ( .A1(n1881), .A2(n1461), .ZN(n1866) );
  NAND2_X1 U1919 ( .A1(n2188), .A2(n2079), .ZN(n1462) );
  NAND3_X1 U1920 ( .A1(n1462), .A2(n1853), .A3(n1553), .ZN(n1601) );
  AOI21_X1 U1921 ( .B1(n1978), .B2(n1463), .A(n1464), .ZN(n2628) );
  INV_X1 U1922 ( .A(n1969), .ZN(n1463) );
  INV_X1 U1923 ( .A(n1613), .ZN(n1464) );
  OAI22_X1 U1924 ( .A1(n1370), .A2(n1919), .B1(n1549), .B2(n2773), .ZN(n1465)
         );
  OAI21_X1 U1925 ( .B1(n1582), .B2(n1543), .A(n2120), .ZN(n1466) );
  NOR2_X1 U1926 ( .A1(n1465), .A2(n1466), .ZN(n2460) );
  XOR2_X1 U1927 ( .A(n2521), .B(n1396), .Z(n2633) );
  OAI211_X1 U1928 ( .C1(n1984), .C2(n2552), .A(n1983), .B(n1982), .ZN(n1467)
         );
  AOI21_X1 U1929 ( .B1(n2534), .B2(n2596), .A(n1467), .ZN(n1468) );
  AOI22_X1 U1930 ( .A1(n2027), .A2(n2593), .B1(n2533), .B2(n2772), .ZN(n1469)
         );
  OAI211_X1 U1931 ( .C1(n2551), .C2(n2545), .A(n1468), .B(n1469), .ZN(n1470)
         );
  INV_X1 U1932 ( .A(n1567), .ZN(n1471) );
  AOI22_X1 U1933 ( .A1(n1567), .A2(n2541), .B1(n2573), .B2(n1471), .ZN(n1472)
         );
  INV_X1 U1934 ( .A(n1628), .ZN(n1473) );
  AOI21_X1 U1936 ( .B1(n2622), .B2(n1470), .A(n1475), .ZN(n1476) );
  OAI21_X1 U1937 ( .B1(n2631), .B2(n2544), .A(n1476), .ZN(n2916) );
  INV_X1 U1938 ( .A(n1839), .ZN(n1477) );
  AOI21_X1 U1939 ( .B1(n1557), .B2(n1840), .A(n1477), .ZN(n2368) );
  INV_X1 U1940 ( .A(n2302), .ZN(n1478) );
  AND3_X1 U1941 ( .A1(n2300), .A2(n2304), .A3(n1478), .ZN(n1658) );
  AND3_X1 U1942 ( .A1(\unit_fetch/pc_regout[22] ), .A2(
        \unit_fetch/pc_regout[21] ), .A3(\unit_fetch/unit_adder/add_19/n89 ), 
        .ZN(\unit_fetch/unit_adder/add_19/n9 ) );
  NAND2_X1 U1943 ( .A1(\unit_fetch/pc_regout[21] ), .A2(
        \unit_fetch/unit_adder/add_19/n89 ), .ZN(n1479) );
  XNOR2_X1 U1944 ( .A(\unit_fetch/pc_regout[22] ), .B(n1479), .ZN(
        \unit_fetch/adder_out[22] ) );
  INV_X1 U1945 ( .A(n1553), .ZN(n1480) );
  OAI21_X1 U1946 ( .B1(n2194), .B2(n2111), .A(n2110), .ZN(n1481) );
  NAND2_X1 U1947 ( .A1(n1851), .A2(n1601), .ZN(n1482) );
  AOI21_X1 U1948 ( .B1(n1480), .B2(n1481), .A(n1482), .ZN(n1852) );
  AOI22_X1 U1949 ( .A1(n2775), .A2(n2605), .B1(n2474), .B2(n2571), .ZN(n1483)
         );
  NAND2_X1 U1950 ( .A1(n2175), .A2(n2135), .ZN(n1484) );
  NAND3_X1 U1951 ( .A1(n1484), .A2(n1483), .A3(n2120), .ZN(n2504) );
  NAND2_X1 U1952 ( .A1(n1912), .A2(n1622), .ZN(n1485) );
  XOR2_X1 U1953 ( .A(n1634), .B(n1485), .Z(n2632) );
  AOI22_X1 U1954 ( .A1(n2534), .A2(n2593), .B1(n2598), .B2(n2027), .ZN(n1486)
         );
  AOI22_X1 U1955 ( .A1(n2607), .A2(n2592), .B1(n2535), .B2(n2594), .ZN(n1487)
         );
  NAND3_X1 U1956 ( .A1(n1940), .A2(n1619), .A3(n2554), .ZN(n1488) );
  OAI211_X1 U1957 ( .C1(n2609), .C2(n2552), .A(n1487), .B(n1488), .ZN(n1489)
         );
  OAI22_X1 U1958 ( .A1(n2548), .A2(n2024), .B1(n2515), .B2(n1984), .ZN(n1490)
         );
  AOI211_X1 U1959 ( .C1(n2537), .C2(n2772), .A(n1489), .B(n1490), .ZN(n1491)
         );
  INV_X1 U1960 ( .A(n1565), .ZN(n1492) );
  AOI22_X1 U1961 ( .A1(n1565), .A2(n2573), .B1(n2570), .B2(n1492), .ZN(n1493)
         );
  INV_X1 U1962 ( .A(\unit_decode/IMMreg/ffi_2/n4 ), .ZN(n1494) );
  AOI21_X1 U1964 ( .B1(n2627), .B2(n2617), .A(n1496), .ZN(n1497) );
  OAI221_X1 U1965 ( .B1(n2780), .B2(n1486), .C1(n2780), .C2(n1491), .A(n1497), 
        .ZN(n2915) );
  INV_X1 U1966 ( .A(n1903), .ZN(n1498) );
  NOR2_X1 U1967 ( .A1(n2303), .A2(n1498), .ZN(n1659) );
  AND3_X1 U1968 ( .A1(n2367), .A2(n1569), .A3(n1877), .ZN(n1784) );
  INV_X1 U1969 ( .A(n2425), .ZN(n1499) );
  AOI21_X1 U1970 ( .B1(n2426), .B2(n2427), .A(n1499), .ZN(n2446) );
  OR2_X1 U1971 ( .A1(n2523), .A2(n1393), .ZN(n1500) );
  NAND2_X1 U1972 ( .A1(n1562), .A2(n1912), .ZN(n1501) );
  AOI21_X1 U1973 ( .B1(n2052), .B2(n1501), .A(n1500), .ZN(n2525) );
  NOR3_X1 U1974 ( .A1(\unit_fetch/unit_adder/add_19/n86 ), .A2(n1640), .A3(
        \unit_fetch/unit_adder/add_19/n54 ), .ZN(n1502) );
  NAND2_X1 U1975 ( .A1(n1637), .A2(n1502), .ZN(n1641) );
  OAI211_X1 U1976 ( .C1(n1865), .C2(n1833), .A(n1863), .B(n1832), .ZN(n1503)
         );
  XOR2_X1 U1977 ( .A(n2307), .B(n2213), .Z(n1504) );
  XNOR2_X1 U1978 ( .A(n1503), .B(n1504), .ZN(n2648) );
  OAI22_X1 U1979 ( .A1(n1920), .A2(n1617), .B1(n1554), .B2(n2030), .ZN(n1505)
         );
  INV_X1 U1980 ( .A(n2029), .ZN(n1506) );
  NOR2_X1 U1981 ( .A1(n1505), .A2(n1506), .ZN(n2760) );
  INV_X1 U1982 ( .A(n1981), .ZN(n1507) );
  OAI21_X1 U1983 ( .B1(n2007), .B2(n1507), .A(n1991), .ZN(n1508) );
  XOR2_X1 U1984 ( .A(n1988), .B(n1628), .Z(n1509) );
  XNOR2_X1 U1985 ( .A(n1508), .B(n1509), .ZN(n2631) );
  AND3_X1 U1986 ( .A1(n1342), .A2(n1690), .A3(n1338), .ZN(n1897) );
  AOI22_X1 U1987 ( .A1(\unit_fetch/adder_out[31] ), .A2(n1927), .B1(n1929), 
        .B2(n2686), .ZN(n1510) );
  OAI21_X1 U1988 ( .B1(\unit_fetch/unit_npcregister/ffi_31/n4 ), .B2(n1922), 
        .A(n1510), .ZN(\unit_fetch/unit_npcregister/ffi_31/n5 ) );
  AND4_X1 U1989 ( .A1(n2828), .A2(n2846), .A3(n2836), .A4(n2831), .ZN(n1511)
         );
  NOR2_X1 U1990 ( .A1(n1933), .A2(n1511), .ZN(
        \unit_fetch/unit_instructionRegister/n80 ) );
  BUF_X2 U1991 ( .A(\unit_fetch/pc_regout[2] ), .Z(n1603) );
  XOR2_X1 U1992 ( .A(n1941), .B(\unit_decode/IMMreg/ffi_14/n4 ), .Z(n1512) );
  INV_X2 U1993 ( .A(n1542), .ZN(n1921) );
  INV_X1 U1994 ( .A(n1542), .ZN(n1922) );
  OR2_X1 U1995 ( .A1(n1528), .A2(n2778), .ZN(n1516) );
  INV_X4 U1996 ( .A(RST), .ZN(n1942) );
  NAND2_X1 U2006 ( .A1(n2472), .A2(n2426), .ZN(n2480) );
  NAND2_X1 U2007 ( .A1(n1526), .A2(n2767), .ZN(n2426) );
  INV_X1 U2008 ( .A(n2197), .ZN(n1526) );
  XNOR2_X1 U2009 ( .A(n2488), .B(n1527), .ZN(n2486) );
  INV_X1 U2010 ( .A(n2196), .ZN(n1527) );
  XNOR2_X1 U2011 ( .A(n1908), .B(\unit_decode/IMMreg/ffi_15/n4 ), .ZN(n2196)
         );
  NAND2_X1 U2012 ( .A1(n2610), .A2(n1653), .ZN(n1529) );
  INV_X1 U2013 ( .A(\unit_control/uut_third_stage/ffi_9/n5 ), .ZN(n1530) );
  INV_X1 U2014 ( .A(n2767), .ZN(n2711) );
  AOI21_X1 U2015 ( .B1(n2075), .B2(n2074), .A(n2073), .ZN(n1531) );
  BUF_X1 U2016 ( .A(n1351), .Z(n1532) );
  BUF_X1 U2017 ( .A(n2493), .Z(n1533) );
  INV_X1 U2018 ( .A(n1575), .ZN(n1534) );
  MUX2_X1 U2019 ( .A(\unit_decode/NPC1reg/ffi_31/n4 ), .B(
        \unit_decode/Areg/ffi_31/n4 ), .S(n1935), .Z(n2587) );
  AND4_X1 U2020 ( .A1(n2133), .A2(n2294), .A3(n2132), .A4(n2131), .ZN(n1535)
         );
  NAND2_X1 U2021 ( .A1(n1760), .A2(n2095), .ZN(n1608) );
  BUF_X1 U2022 ( .A(n2445), .Z(n1536) );
  OAI21_X1 U2023 ( .B1(n2472), .B2(n2473), .A(n2425), .ZN(n2445) );
  OR3_X1 U2024 ( .A1(n2160), .A2(n2159), .A3(n2174), .ZN(n1537) );
  XNOR2_X1 U2025 ( .A(n1915), .B(n1665), .ZN(n1538) );
  OAI211_X1 U2026 ( .C1(n2051), .C2(n2050), .A(n2049), .B(n2048), .ZN(n1539)
         );
  OR2_X1 U2027 ( .A1(n1769), .A2(n2414), .ZN(n1649) );
  BUF_X1 U2028 ( .A(n1715), .Z(n1540) );
  XOR2_X1 U2029 ( .A(n1722), .B(n2431), .Z(n2437) );
  AND2_X1 U2030 ( .A1(n1366), .A2(n1942), .ZN(n1541) );
  CLKBUF_X3 U2031 ( .A(n2927), .Z(n1932) );
  INV_X1 U2032 ( .A(n2708), .ZN(n1542) );
  BUF_X1 U2033 ( .A(n2125), .Z(n1543) );
  MUX2_X1 U2034 ( .A(\unit_decode/Areg/ffi_5/n4 ), .B(
        \unit_decode/NPC1reg/ffi_5/n4 ), .S(n1757), .Z(n2161) );
  BUF_X1 U2035 ( .A(n2497), .Z(n1545) );
  INV_X1 U2036 ( .A(n1589), .ZN(n1546) );
  AND2_X1 U2037 ( .A1(n1386), .A2(n1545), .ZN(n1548) );
  XOR2_X1 U2038 ( .A(n1643), .B(n2202), .Z(n2431) );
  BUF_X2 U2039 ( .A(n2574), .Z(n1549) );
  BUF_X1 U2040 ( .A(n2625), .Z(n1550) );
  BUF_X1 U2041 ( .A(n1381), .Z(n1551) );
  AND2_X1 U2042 ( .A1(n1770), .A2(n1578), .ZN(n1552) );
  XOR2_X1 U2043 ( .A(n2192), .B(n2228), .Z(n1553) );
  BUF_X2 U2044 ( .A(n2228), .Z(n1554) );
  BUF_X1 U2045 ( .A(n2008), .Z(n1555) );
  XNOR2_X1 U2046 ( .A(n1556), .B(n1616), .ZN(n2053) );
  XNOR2_X1 U2047 ( .A(n1623), .B(\unit_decode/IMMreg/ffi_9/n4 ), .ZN(n2067) );
  NAND2_X1 U2048 ( .A1(n2417), .A2(n2200), .ZN(n1557) );
  MUX2_X1 U2049 ( .A(\unit_decode/NPC1reg/ffi_5/n4 ), .B(
        \unit_decode/Areg/ffi_5/n4 ), .S(n1911), .Z(n1558) );
  BUF_X1 U2050 ( .A(n1934), .Z(n1560) );
  BUF_X1 U2051 ( .A(\unit_control/uut_third_stage/ffi_9/n5 ), .Z(n1561) );
  BUF_X1 U2052 ( .A(n1350), .Z(n1590) );
  BUF_X1 U2053 ( .A(n2045), .Z(n1562) );
  OR2_X2 U2054 ( .A1(n2162), .A2(n1512), .ZN(n2109) );
  OR2_X1 U2055 ( .A1(n1606), .A2(n1924), .ZN(n1563) );
  NAND2_X1 U2056 ( .A1(n1563), .A2(n1564), .ZN(
        \unit_fetch/unit_programCounter/ffi_31/n5 ) );
  AOI22_X1 U2057 ( .A1(n2686), .A2(n1929), .B1(\unit_fetch/adder_out[31] ), 
        .B2(n1926), .ZN(n1564) );
  INV_X1 U2058 ( .A(n2607), .ZN(n1565) );
  BUF_X1 U2059 ( .A(n2645), .Z(n1566) );
  INV_X1 U2060 ( .A(n1662), .ZN(n1567) );
  XNOR2_X1 U2061 ( .A(n2150), .B(n1756), .ZN(n1568) );
  OR2_X1 U2062 ( .A1(n2423), .A2(n1701), .ZN(n1570) );
  AND4_X1 U2063 ( .A1(n2770), .A2(n1585), .A3(n2769), .A4(n1584), .ZN(n1571)
         );
  OR2_X1 U2064 ( .A1(n1676), .A2(n1602), .ZN(n1572) );
  AND2_X1 U2065 ( .A1(n1581), .A2(n1860), .ZN(n1573) );
  XNOR2_X1 U2066 ( .A(n2318), .B(n1574), .ZN(n2647) );
  INV_X1 U2067 ( .A(n2708), .ZN(n1925) );
  INV_X1 U2068 ( .A(n1732), .ZN(n2507) );
  BUF_X1 U2069 ( .A(n2289), .Z(n1918) );
  CLKBUF_X3 U2070 ( .A(n1932), .Z(n1933) );
  AND2_X1 U2071 ( .A1(n2029), .A2(n1995), .ZN(n2757) );
  AND2_X1 U2072 ( .A1(n2029), .A2(n1948), .ZN(n2549) );
  INV_X1 U2073 ( .A(n2741), .ZN(n2816) );
  AND3_X1 U2074 ( .A1(n1889), .A2(n1804), .A3(n1803), .ZN(n1700) );
  AND2_X1 U2075 ( .A1(n2029), .A2(n1953), .ZN(n2601) );
  NAND2_X1 U2076 ( .A1(n1811), .A2(n1810), .ZN(n2786) );
  INV_X1 U2077 ( .A(n2875), .ZN(n2889) );
  BUF_X1 U2078 ( .A(n2875), .Z(n1587) );
  INV_X1 U2079 ( .A(n2598), .ZN(n2545) );
  INV_X1 U2080 ( .A(n2782), .ZN(n1810) );
  INV_X1 U2081 ( .A(n2596), .ZN(n2548) );
  OAI21_X1 U2082 ( .B1(n2737), .B2(\unit_fetch/unit_instructionRegister/n55 ), 
        .A(n2715), .ZN(n2782) );
  INV_X1 U2083 ( .A(n2193), .ZN(n1592) );
  NAND2_X1 U2084 ( .A1(n2732), .A2(n1891), .ZN(n2875) );
  OAI21_X1 U2085 ( .B1(n2824), .B2(n2733), .A(n2813), .ZN(n2929) );
  INV_X1 U2086 ( .A(n2777), .ZN(n2592) );
  INV_X1 U2087 ( .A(n2319), .ZN(n1574) );
  INV_X1 U2088 ( .A(n2774), .ZN(n2772) );
  INV_X1 U2089 ( .A(n2729), .ZN(n2732) );
  INV_X1 U2090 ( .A(n2611), .ZN(n2541) );
  XNOR2_X1 U2091 ( .A(n2210), .B(n1797), .ZN(n1883) );
  INV_X1 U2092 ( .A(n2736), .ZN(n2737) );
  INV_X1 U2093 ( .A(n1643), .ZN(n2432) );
  INV_X1 U2094 ( .A(n2587), .ZN(n1575) );
  NAND3_X1 U2095 ( .A1(n2712), .A2(\unit_fetch/unit_instructionRegister/n64 ), 
        .A3(n1333), .ZN(n2736) );
  OR2_X1 U2096 ( .A1(n2143), .A2(n2123), .ZN(n2291) );
  INV_X1 U2097 ( .A(n2778), .ZN(n2573) );
  INV_X1 U2098 ( .A(n2779), .ZN(n2570) );
  NAND2_X1 U2099 ( .A1(n1896), .A2(\unit_fetch/unit_programCounter/ffi_3/n4 ), 
        .ZN(n2729) );
  AND4_X1 U2100 ( .A1(\unit_fetch/unit_programCounter/ffi_18/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_20/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_28/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_10/n4 ), .ZN(n1677) );
  INV_X1 U2101 ( .A(n2713), .ZN(n2712) );
  OR3_X1 U2102 ( .A1(\unit_fetch/unit_instructionRegister/n64 ), .A2(n1333), 
        .A3(n2713), .ZN(n2735) );
  INV_X1 U2103 ( .A(n2776), .ZN(n1576) );
  INV_X1 U2104 ( .A(n2617), .ZN(n2544) );
  INV_X1 U2105 ( .A(\unit_fetch/unit_programCounter/ffi_4/n4 ), .ZN(n1896) );
  INV_X1 U2106 ( .A(n2780), .ZN(n2622) );
  NOR2_X1 U2107 ( .A1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .ZN(n2869) );
  NAND3_X1 U2108 ( .A1(n1331), .A2(\unit_fetch/unit_instructionRegister/n65 ), 
        .A3(\unit_fetch/unit_instructionRegister/n66 ), .ZN(n2713) );
  OR2_X1 U2109 ( .A1(n1538), .A2(n1966), .ZN(n2552) );
  INV_X1 U2110 ( .A(n2552), .ZN(n1577) );
  NAND2_X1 U2111 ( .A1(n1770), .A2(n1578), .ZN(n2262) );
  NOR2_X1 U2112 ( .A1(n1579), .A2(n1573), .ZN(n1578) );
  OAI21_X1 U2113 ( .B1(n1903), .B2(n1572), .A(n1859), .ZN(n1579) );
  NAND4_X1 U2114 ( .A1(n1812), .A2(n1364), .A3(n1898), .A4(n1813), .ZN(n2650)
         );
  AND4_X2 U2115 ( .A1(n1884), .A2(n1835), .A3(n1836), .A4(n2649), .ZN(n1812)
         );
  NOR2_X1 U2116 ( .A1(n2624), .A2(n2623), .ZN(n1875) );
  XNOR2_X1 U2117 ( .A(n2058), .B(n2498), .ZN(n2623) );
  XNOR2_X1 U2118 ( .A(n1349), .B(\unit_fetch/unit_programCounter/ffi_21/n4 ), 
        .ZN(\unit_fetch/adder_out[21] ) );
  NAND2_X1 U2119 ( .A1(n1571), .A2(n1583), .ZN(n2771) );
  INV_X1 U2120 ( .A(n2139), .ZN(n1583) );
  NAND2_X1 U2121 ( .A1(n2465), .A2(n2592), .ZN(n1584) );
  INV_X1 U2122 ( .A(n2140), .ZN(n1585) );
  XNOR2_X1 U2123 ( .A(n2067), .B(n2151), .ZN(n2494) );
  OAI21_X1 U2124 ( .B1(n1911), .B2(n1515), .A(n1586), .ZN(n2151) );
  NAND2_X1 U2125 ( .A1(n1914), .A2(\unit_decode/Areg/ffi_9/n4 ), .ZN(n1586) );
  NAND2_X1 U2126 ( .A1(n2791), .A2(n2829), .ZN(n2728) );
  NOR2_X1 U2127 ( .A1(n2729), .A2(n1588), .ZN(n2791) );
  AND2_X1 U2128 ( .A1(n1603), .A2(\unit_fetch/pc_regout[1] ), .ZN(n1588) );
  NAND2_X1 U2129 ( .A1(n1593), .A2(n1591), .ZN(n1594) );
  NOR2_X1 U2130 ( .A1(n1570), .A2(n2193), .ZN(n1591) );
  NAND2_X1 U2131 ( .A1(n1553), .A2(n2194), .ZN(n1593) );
  AND2_X1 U2132 ( .A1(n1593), .A2(n1592), .ZN(n2484) );
  XNOR2_X1 U2133 ( .A(n2192), .B(n2228), .ZN(n2485) );
  NOR2_X1 U2134 ( .A1(n1829), .A2(n1594), .ZN(n1876) );
  OAI21_X1 U2135 ( .B1(n2109), .B2(n1595), .A(n1760), .ZN(n2194) );
  INV_X1 U2136 ( .A(n2095), .ZN(n1595) );
  NAND2_X1 U2137 ( .A1(n2046), .A2(n2045), .ZN(n2075) );
  XNOR2_X1 U2138 ( .A(n2172), .B(n2019), .ZN(n2051) );
  OAI21_X1 U2139 ( .B1(n1513), .B2(n1934), .A(n1596), .ZN(n2172) );
  NAND2_X1 U2140 ( .A1(n1911), .A2(\unit_decode/Areg/ffi_6/n4 ), .ZN(n1596) );
  NAND2_X1 U2141 ( .A1(n1597), .A2(n1598), .ZN(n2046) );
  AOI21_X1 U2142 ( .B1(n2005), .B2(n1555), .A(n2565), .ZN(n1597) );
  NOR2_X1 U2143 ( .A1(n2562), .A2(n2574), .ZN(n2565) );
  NAND2_X1 U2144 ( .A1(n1991), .A2(n1990), .ZN(n2005) );
  NAND4_X1 U2145 ( .A1(n1651), .A2(n1695), .A3(n1657), .A4(n1649), .ZN(n1599)
         );
  XNOR2_X1 U2146 ( .A(n1837), .B(n1373), .ZN(n1651) );
  XNOR2_X1 U2147 ( .A(n2487), .B(n1600), .ZN(n1657) );
  INV_X1 U2148 ( .A(n1719), .ZN(n1600) );
  OAI21_X1 U2149 ( .B1(n1882), .B2(n1838), .A(n1659), .ZN(n1739) );
  NAND2_X1 U2150 ( .A1(n1620), .A2(n1394), .ZN(n1882) );
  NAND3_X1 U2151 ( .A1(n1395), .A2(n1828), .A3(n2484), .ZN(n1620) );
  NAND2_X1 U2152 ( .A1(n1635), .A2(n1708), .ZN(n1834) );
  NAND3_X1 U2153 ( .A1(n1635), .A2(n1708), .A3(n1880), .ZN(n1879) );
  NAND2_X1 U2154 ( .A1(n1601), .A2(n2484), .ZN(n2487) );
  NOR2_X1 U2155 ( .A1(n2191), .A2(n2501), .ZN(n2079) );
  NAND2_X1 U2156 ( .A1(n2195), .A2(n1876), .ZN(n1609) );
  INV_X1 U2157 ( .A(n1860), .ZN(n1602) );
  OAI21_X1 U2158 ( .B1(n1906), .B2(n1694), .A(n1905), .ZN(n1903) );
  OR2_X1 U2159 ( .A1(RST), .A2(n2142), .ZN(n2708) );
  OAI211_X1 U2160 ( .C1(n1886), .C2(\unit_control/n152 ), .A(n1799), .B(n1798), 
        .ZN(n2142) );
  NAND2_X1 U2161 ( .A1(n1607), .A2(n1603), .ZN(n1604) );
  BUF_X1 U2162 ( .A(n2795), .Z(n1605) );
  INV_X1 U2163 ( .A(n1892), .ZN(n2878) );
  XNOR2_X1 U2164 ( .A(\unit_fetch/unit_adder/add_19/n1 ), .B(n1606), .ZN(
        \unit_fetch/adder_out[31] ) );
  BUF_X1 U2165 ( .A(\unit_fetch/pc_regout[3] ), .Z(n1607) );
  BUF_X1 U2166 ( .A(n2649), .Z(n1610) );
  AND2_X1 U2167 ( .A1(n2655), .A2(n2654), .ZN(n1611) );
  INV_X1 U2168 ( .A(n1646), .ZN(n2542) );
  NAND2_X1 U2169 ( .A1(n1568), .A2(n1969), .ZN(n1613) );
  OR3_X1 U2170 ( .A1(n2794), .A2(n2929), .A3(
        \unit_fetch/unit_instructionRegister/n70 ), .ZN(n1614) );
  INV_X1 U2171 ( .A(n2925), .ZN(n2794) );
  BUF_X1 U2172 ( .A(n2494), .Z(n1615) );
  BUF_X2 U2173 ( .A(n1915), .Z(n1616) );
  AND2_X1 U2174 ( .A1(n1951), .A2(n1538), .ZN(n2593) );
  INV_X1 U2175 ( .A(n1941), .ZN(n1937) );
  INV_X1 U2176 ( .A(n1618), .ZN(n1617) );
  INV_X1 U2177 ( .A(n1628), .ZN(n1619) );
  INV_X1 U2178 ( .A(n2147), .ZN(n2603) );
  BUF_X1 U2179 ( .A(n2738), .Z(n1621) );
  AOI211_X1 U2180 ( .C1(n2814), .C2(n2745), .A(n2783), .B(n2795), .ZN(n2738)
         );
  BUF_X1 U2181 ( .A(n2564), .Z(n1622) );
  BUF_X2 U2182 ( .A(n1911), .Z(n1935) );
  CLKBUF_X3 U2183 ( .A(\unit_control/uut_third_stage/ffi_19/n5 ), .Z(n1910) );
  BUF_X1 U2184 ( .A(\unit_control/uut_third_stage/ffi_9/n5 ), .Z(n1623) );
  INV_X1 U2185 ( .A(n2612), .ZN(n1624) );
  NAND2_X1 U2186 ( .A1(n1755), .A2(n1758), .ZN(n2610) );
  INV_X1 U2187 ( .A(n1941), .ZN(n1938) );
  CLKBUF_X3 U2188 ( .A(n1941), .Z(n1940) );
  INV_X1 U2189 ( .A(n1941), .ZN(n1909) );
  AND4_X1 U2190 ( .A1(n1812), .A2(n1898), .A3(n1813), .A4(n1815), .ZN(n1625)
         );
  INV_X1 U2191 ( .A(n2098), .ZN(n1626) );
  BUF_X1 U2192 ( .A(n2051), .Z(n1627) );
  NAND2_X1 U2193 ( .A1(n1367), .A2(n1942), .ZN(n2927) );
  INV_X1 U2194 ( .A(n2603), .ZN(n1628) );
  OAI21_X1 U2195 ( .B1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .B2(n2822), 
        .A(n2889), .ZN(n2818) );
  NAND2_X1 U2196 ( .A1(n2818), .A2(n2828), .ZN(n2741) );
  INV_X1 U2197 ( .A(n2090), .ZN(n1629) );
  INV_X1 U2198 ( .A(n1544), .ZN(n1630) );
  OR2_X1 U2199 ( .A1(n2738), .A2(\unit_control/n152 ), .ZN(n1798) );
  INV_X1 U2200 ( .A(n2082), .ZN(n1631) );
  INV_X1 U2201 ( .A(n2251), .ZN(n1633) );
  BUF_X1 U2202 ( .A(n2010), .Z(n1634) );
  AOI21_X1 U2203 ( .B1(n1632), .B2(n2445), .A(n2428), .ZN(n1635) );
  BUF_X1 U2204 ( .A(n2565), .Z(n1636) );
  INV_X1 U2205 ( .A(\unit_fetch/pc_regout[19] ), .ZN(
        \unit_fetch/unit_adder/add_19/n17 ) );
  INV_X1 U2206 ( .A(\unit_fetch/pc_regout[17] ), .ZN(
        \unit_fetch/unit_adder/add_19/n28 ) );
  INV_X1 U2207 ( .A(\unit_fetch/pc_regout[16] ), .ZN(
        \unit_fetch/unit_adder/add_19/n32 ) );
  INV_X1 U2208 ( .A(\unit_fetch/unit_adder/add_19/n35 ), .ZN(
        \unit_fetch/unit_adder/add_19/n34 ) );
  INV_X1 U2209 ( .A(\unit_fetch/pc_regout[15] ), .ZN(
        \unit_fetch/unit_adder/add_19/n37 ) );
  INV_X1 U2210 ( .A(\unit_fetch/pc_regout[14] ), .ZN(
        \unit_fetch/unit_adder/add_19/n41 ) );
  INV_X1 U2211 ( .A(\unit_fetch/unit_adder/add_19/n43 ), .ZN(
        \unit_fetch/unit_adder/add_19/n42 ) );
  INV_X1 U2212 ( .A(\unit_fetch/unit_adder/add_19/n54 ), .ZN(
        \unit_fetch/unit_adder/add_19/n53 ) );
  INV_X1 U2213 ( .A(\unit_fetch/unit_adder/add_19/n78 ), .ZN(
        \unit_fetch/unit_adder/add_19/n77 ) );
  INV_X1 U2214 ( .A(\unit_fetch/pc_regout[5] ), .ZN(
        \unit_fetch/unit_adder/add_19/n81 ) );
  INV_X1 U2215 ( .A(\unit_fetch/pc_regout[4] ), .ZN(
        \unit_fetch/unit_adder/add_19/n84 ) );
  INV_X1 U2216 ( .A(n1604), .ZN(\unit_fetch/unit_adder/add_19/n85 ) );
  NAND3_X1 U2217 ( .A1(n1638), .A2(\unit_fetch/unit_adder/add_19/n12 ), .A3(
        n1637), .ZN(n1639) );
  AND2_X1 U2218 ( .A1(n1637), .A2(\unit_fetch/unit_adder/add_19/n78 ), .ZN(
        n1642) );
  NOR2_X1 U2219 ( .A1(\unit_fetch/unit_adder/add_19/n54 ), .A2(
        \unit_fetch/unit_adder/add_19/n86 ), .ZN(n1638) );
  NOR2_X1 U2220 ( .A1(\unit_fetch/unit_adder/add_19/n63 ), .A2(
        \unit_fetch/unit_adder/add_19/n70 ), .ZN(n1637) );
  NOR2_X1 U2221 ( .A1(n1639), .A2(n1640), .ZN(
        \unit_fetch/unit_adder/add_19/n89 ) );
  NOR2_X1 U2222 ( .A1(\unit_fetch/unit_adder/add_19/n79 ), .A2(n1604), .ZN(
        \unit_fetch/unit_adder/add_19/n78 ) );
  NOR2_X1 U2223 ( .A1(\unit_fetch/unit_adder/add_19/n54 ), .A2(
        \unit_fetch/unit_adder/add_19/n45 ), .ZN(
        \unit_fetch/unit_adder/add_19/n44 ) );
  INV_X1 U2224 ( .A(n1649), .ZN(n2641) );
  MUX2_X1 U2225 ( .A(n1644), .B(n1645), .S(n1934), .Z(n1643) );
  BUF_X2 U2226 ( .A(\unit_control/uut_third_stage/ffi_19/n5 ), .Z(n1911) );
  NOR2_X1 U2227 ( .A1(n2908), .A2(n1603), .ZN(n2845) );
  AOI211_X4 U2228 ( .C1(n2789), .C2(\unit_fetch/pc_regout[3] ), .A(n2790), .B(
        n2730), .ZN(n2924) );
  MUX2_X1 U2229 ( .A(\unit_decode/Areg/ffi_2/n4 ), .B(
        \unit_decode/NPC1reg/ffi_2/n4 ), .S(n1913), .Z(n2154) );
  MUX2_X1 U2230 ( .A(n1647), .B(n1648), .S(n1757), .Z(n1646) );
  INV_X1 U2231 ( .A(n1616), .ZN(n1936) );
  OAI21_X1 U2232 ( .B1(n2494), .B2(n2069), .A(n2495), .ZN(n2493) );
  INV_X1 U2233 ( .A(n1913), .ZN(n1914) );
  AND2_X2 U2234 ( .A1(n1873), .A2(n1872), .ZN(n2588) );
  NAND3_X1 U2235 ( .A1(n1848), .A2(n1611), .A3(n1849), .ZN(n2707) );
  NOR2_X1 U2236 ( .A1(n2927), .A2(n1383), .ZN(n2710) );
  AND2_X1 U2237 ( .A1(n1383), .A2(n1541), .ZN(n2709) );
  OR3_X1 U2238 ( .A1(n2081), .A2(n2080), .A3(n1733), .ZN(n1732) );
  BUF_X2 U2239 ( .A(n2709), .Z(n1927) );
  INV_X1 U2240 ( .A(n2775), .ZN(n2248) );
  BUF_X2 U2241 ( .A(n2710), .Z(n1930) );
  BUF_X2 U2242 ( .A(n2709), .Z(n1926) );
  BUF_X2 U2243 ( .A(n2710), .Z(n1929) );
  XNOR2_X1 U2244 ( .A(n2734), .B(n2929), .ZN(n2795) );
  NOR2_X1 U2245 ( .A1(n2794), .A2(n2924), .ZN(n2734) );
  NOR2_X1 U2246 ( .A1(\unit_fetch/unit_programCounter/ffi_5/n4 ), .A2(n2876), 
        .ZN(n2790) );
  AOI221_X1 U2247 ( .B1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n2845), 
        .C1(\unit_fetch/pc_regout[1] ), .C2(n2845), .A(n2729), .ZN(n2730) );
  OAI211_X1 U2248 ( .C1(n1896), .C2(\unit_fetch/unit_programCounter/ffi_3/n4 ), 
        .A(n2728), .B(n2727), .ZN(n2925) );
  NOR3_X1 U2249 ( .A1(n2816), .A2(n2723), .A3(n2782), .ZN(n2740) );
  NOR2_X1 U2250 ( .A1(\unit_decode/RD1reg/ffi_1/n4 ), .A2(n2786), .ZN(n2723)
         );
  NOR2_X1 U2251 ( .A1(n2724), .A2(n2745), .ZN(n1811) );
  OAI221_X1 U2252 ( .B1(n2737), .B2(\unit_fetch/unit_instructionRegister/n60 ), 
        .C1(n2736), .C2(\unit_fetch/unit_instructionRegister/n53 ), .A(n2735), 
        .ZN(n2745) );
  INV_X1 U2253 ( .A(\unit_fetch/unit_programCounter/ffi_11/n4 ), .ZN(n2861) );
  NAND2_X1 U2254 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(n2869), 
        .ZN(n2876) );
  NOR2_X1 U2255 ( .A1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .A2(
        \unit_fetch/pc_regout[0] ), .ZN(n2908) );
  INV_X1 U2256 ( .A(n2901), .ZN(n2867) );
  NOR2_X1 U2257 ( .A1(n2819), .A2(n2825), .ZN(n2901) );
  INV_X1 U2258 ( .A(n2593), .ZN(n2550) );
  INV_X1 U2259 ( .A(n2289), .ZN(n2175) );
  AND2_X1 U2260 ( .A1(n1671), .A2(n1336), .ZN(n2617) );
  AND2_X1 U2261 ( .A1(n1577), .A2(n2622), .ZN(n2606) );
  INV_X1 U2262 ( .A(RST), .ZN(n1943) );
  NAND2_X1 U2263 ( .A1(n2572), .A2(n1655), .ZN(n2779) );
  NAND2_X1 U2264 ( .A1(n1341), .A2(n1336), .ZN(n2780) );
  INV_X1 U2265 ( .A(n2932), .ZN(n2808) );
  BUF_X2 U2266 ( .A(n2710), .Z(n1931) );
  BUF_X2 U2267 ( .A(n2709), .Z(n1928) );
  AND2_X1 U2268 ( .A1(n2706), .A2(n1942), .ZN(n2944) );
  AND2_X1 U2269 ( .A1(n2700), .A2(n1942), .ZN(n2957) );
  AND2_X1 U2270 ( .A1(n2699), .A2(n1943), .ZN(n2958) );
  AND2_X1 U2271 ( .A1(n2694), .A2(n1942), .ZN(n2963) );
  AND2_X1 U2272 ( .A1(n2696), .A2(n1942), .ZN(n2961) );
  AND2_X1 U2273 ( .A1(n2689), .A2(n1943), .ZN(n2968) );
  AND2_X1 U2274 ( .A1(n2695), .A2(n1942), .ZN(n2962) );
  AND2_X1 U2275 ( .A1(n2697), .A2(n1942), .ZN(n2960) );
  AND2_X1 U2276 ( .A1(n2690), .A2(n1943), .ZN(n2967) );
  AND2_X1 U2277 ( .A1(n2693), .A2(n1942), .ZN(n2964) );
  AND2_X1 U2278 ( .A1(n2692), .A2(n1943), .ZN(n2965) );
  AND2_X1 U2279 ( .A1(n2691), .A2(n1942), .ZN(n2966) );
  AND2_X1 U2280 ( .A1(n2703), .A2(n1942), .ZN(n2951) );
  AND2_X1 U2281 ( .A1(n2704), .A2(n1942), .ZN(n2950) );
  AND2_X1 U2282 ( .A1(n2701), .A2(n1942), .ZN(n2956) );
  AND2_X1 U2283 ( .A1(n2702), .A2(n1942), .ZN(n2955) );
  AND2_X1 U2284 ( .A1(n2688), .A2(n1942), .ZN(n2969) );
  AND2_X1 U2285 ( .A1(n2705), .A2(n1942), .ZN(n2948) );
  AND2_X1 U2286 ( .A1(n2687), .A2(n1943), .ZN(n2970) );
  AND2_X1 U2287 ( .A1(n2686), .A2(n1943), .ZN(n2971) );
  AND2_X1 U2288 ( .A1(n2698), .A2(n1942), .ZN(n2959) );
  NAND4_X1 U2289 ( .A1(n1976), .A2(n1975), .A3(n1974), .A4(n1973), .ZN(n2910)
         );
  NAND2_X1 U2290 ( .A1(n2570), .A2(n1664), .ZN(n1971) );
  AOI22_X1 U2291 ( .A1(n2602), .A2(n2553), .B1(n2595), .B2(n1740), .ZN(n1975)
         );
  NAND2_X1 U2292 ( .A1(n1960), .A2(n2622), .ZN(n1976) );
  OAI21_X1 U2293 ( .B1(n2774), .B2(n2549), .A(n1959), .ZN(n1960) );
  AOI211_X1 U2294 ( .C1(n2596), .C2(n2594), .A(n1958), .B(n1957), .ZN(n1959)
         );
  NOR2_X1 U2295 ( .A1(n2601), .A2(n2545), .ZN(n1957) );
  OAI22_X1 U2296 ( .A1(n2760), .A2(n2558), .B1(n2757), .B2(n2515), .ZN(n2516)
         );
  OAI22_X1 U2297 ( .A1(n2551), .A2(n2777), .B1(n2529), .B2(n2548), .ZN(n2517)
         );
  OAI22_X1 U2298 ( .A1(n2546), .A2(n2528), .B1(n2514), .B2(n2545), .ZN(n2518)
         );
  OAI21_X1 U2299 ( .B1(n2547), .B2(n2552), .A(n2513), .ZN(n2519) );
  AOI22_X1 U2300 ( .A1(n2512), .A2(n2772), .B1(n2593), .B2(n2511), .ZN(n2513)
         );
  OAI211_X1 U2301 ( .C1(\unit_fetch/unit_programCounter/ffi_30/n4 ), .C2(n1924), .A(n2657), .B(n2656), .ZN(\unit_fetch/unit_programCounter/ffi_30/n5 ) );
  OAI211_X1 U2302 ( .C1(\unit_fetch/unit_npcregister/ffi_30/n4 ), .C2(n1924), 
        .A(n2657), .B(n2656), .ZN(\unit_fetch/unit_npcregister/ffi_30/n5 ) );
  NAND2_X1 U2303 ( .A1(n1927), .A2(\unit_fetch/adder_out[30] ), .ZN(n2656) );
  OAI211_X1 U2304 ( .C1(n2247), .C2(n2780), .A(n2246), .B(n2245), .ZN(n2687)
         );
  AOI21_X1 U2305 ( .B1(n2326), .B2(n2244), .A(n2243), .ZN(n2245) );
  NOR3_X1 U2306 ( .A1(n2779), .A2(n2244), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2243) );
  NAND2_X1 U2307 ( .A1(n2653), .A2(n2617), .ZN(n2246) );
  NOR3_X1 U2308 ( .A1(n2238), .A2(n2237), .A3(n2236), .ZN(n2247) );
  OAI22_X1 U2309 ( .A1(n2323), .A2(n2558), .B1(n2313), .B2(n2548), .ZN(n2236)
         );
  OAI22_X1 U2310 ( .A1(n2349), .A2(n2552), .B1(n2282), .B2(n2515), .ZN(n2237)
         );
  OAI211_X1 U2311 ( .C1(n2381), .C2(n2777), .A(n2235), .B(n2234), .ZN(n2238)
         );
  AOI22_X1 U2312 ( .A1(n2233), .A2(n2598), .B1(n2772), .B2(n2232), .ZN(n2234)
         );
  INV_X1 U2313 ( .A(n2257), .ZN(n2233) );
  AOI22_X1 U2314 ( .A1(n2231), .A2(n2593), .B1(n2554), .B2(n2320), .ZN(n2235)
         );
  INV_X1 U2315 ( .A(n2285), .ZN(n2231) );
  OAI21_X1 U2316 ( .B1(\unit_fetch/unit_programCounter/ffi_22/n4 ), .B2(n1924), 
        .A(n2665), .ZN(\unit_fetch/unit_programCounter/ffi_22/n5 ) );
  OAI21_X1 U2317 ( .B1(\unit_fetch/unit_programCounter/ffi_24/n4 ), .B2(n1924), 
        .A(n2663), .ZN(\unit_fetch/unit_programCounter/ffi_24/n5 ) );
  OAI21_X1 U2318 ( .B1(\unit_fetch/unit_programCounter/ffi_25/n4 ), .B2(n1924), 
        .A(n2662), .ZN(\unit_fetch/unit_programCounter/ffi_25/n5 ) );
  OAI21_X1 U2319 ( .B1(\unit_fetch/unit_programCounter/ffi_20/n4 ), .B2(n1923), 
        .A(n2667), .ZN(\unit_fetch/unit_programCounter/ffi_20/n5 ) );
  OAI21_X1 U2320 ( .B1(\unit_fetch/unit_programCounter/ffi_23/n4 ), .B2(n1923), 
        .A(n2664), .ZN(\unit_fetch/unit_programCounter/ffi_23/n5 ) );
  OAI21_X1 U2321 ( .B1(\unit_fetch/unit_programCounter/ffi_21/n4 ), .B2(n1923), 
        .A(n2666), .ZN(\unit_fetch/unit_programCounter/ffi_21/n5 ) );
  OAI21_X1 U2322 ( .B1(\unit_fetch/unit_npcregister/ffi_22/n4 ), .B2(n1921), 
        .A(n2665), .ZN(\unit_fetch/unit_npcregister/ffi_22/n5 ) );
  AOI22_X1 U2323 ( .A1(n1930), .A2(n2695), .B1(n1927), .B2(
        \unit_fetch/adder_out[22] ), .ZN(n2665) );
  OAI21_X1 U2324 ( .B1(n2385), .B2(n2780), .A(n1792), .ZN(n2695) );
  INV_X1 U2325 ( .A(n1793), .ZN(n1792) );
  OAI21_X1 U2326 ( .B1(n1374), .B2(n2544), .A(n1794), .ZN(n1793) );
  AOI21_X1 U2327 ( .B1(n2387), .B2(n1347), .A(n2386), .ZN(n1794) );
  NOR3_X1 U2328 ( .A1(n2779), .A2(n2388), .A3(\unit_decode/IMMreg/ffi_22/n4 ), 
        .ZN(n2386) );
  NOR3_X1 U2329 ( .A1(n2384), .A2(n2383), .A3(n2382), .ZN(n2385) );
  OAI22_X1 U2330 ( .A1(n2438), .A2(n2515), .B1(n2381), .B2(n2505), .ZN(n2382)
         );
  OAI22_X1 U2331 ( .A1(n2410), .A2(n2548), .B1(n1535), .B2(n2558), .ZN(n2383)
         );
  OAI211_X1 U2332 ( .C1(n2468), .C2(n2552), .A(n2380), .B(n2379), .ZN(n2384)
         );
  AOI22_X1 U2333 ( .A1(n2592), .A2(n2394), .B1(n2463), .B2(n2554), .ZN(n2379)
         );
  AOI22_X1 U2334 ( .A1(n2405), .A2(n2593), .B1(n2598), .B2(n2393), .ZN(n2380)
         );
  OAI21_X1 U2335 ( .B1(\unit_fetch/unit_npcregister/ffi_20/n4 ), .B2(n1921), 
        .A(n2667), .ZN(\unit_fetch/unit_npcregister/ffi_20/n5 ) );
  AOI22_X1 U2336 ( .A1(n1930), .A2(n2697), .B1(n1928), .B2(
        \unit_fetch/adder_out[20] ), .ZN(n2667) );
  OAI211_X1 U2337 ( .C1(n2422), .C2(n2780), .A(n2421), .B(n2420), .ZN(n2697)
         );
  NAND2_X1 U2338 ( .A1(n2570), .A2(n1678), .ZN(n2418) );
  NAND2_X1 U2339 ( .A1(n2641), .A2(n2617), .ZN(n2421) );
  NOR3_X1 U2340 ( .A1(n2413), .A2(n2412), .A3(n2411), .ZN(n2422) );
  OAI22_X1 U2341 ( .A1(n2410), .A2(n2545), .B1(n2438), .B2(n2548), .ZN(n2411)
         );
  OAI22_X1 U2342 ( .A1(n2439), .A2(n2515), .B1(n2462), .B2(n2552), .ZN(n2412)
         );
  OAI211_X1 U2343 ( .C1(n2468), .C2(n2558), .A(n2409), .B(n2408), .ZN(n2413)
         );
  AOI22_X1 U2344 ( .A1(n2407), .A2(n2592), .B1(n2554), .B2(n2406), .ZN(n2408)
         );
  AOI22_X1 U2345 ( .A1(n2405), .A2(n2772), .B1(n2593), .B2(n2404), .ZN(n2409)
         );
  OAI21_X1 U2346 ( .B1(\unit_fetch/unit_npcregister/ffi_23/n4 ), .B2(n1921), 
        .A(n2664), .ZN(\unit_fetch/unit_npcregister/ffi_23/n5 ) );
  AOI22_X1 U2347 ( .A1(n1931), .A2(n2694), .B1(n1928), .B2(
        \unit_fetch/adder_out[23] ), .ZN(n2664) );
  OAI211_X1 U2348 ( .C1(n2378), .C2(n2780), .A(n2377), .B(n2376), .ZN(n2694)
         );
  AOI21_X1 U2349 ( .B1(n2375), .B2(n2374), .A(n2373), .ZN(n2376) );
  NOR3_X1 U2350 ( .A1(n2779), .A2(n2374), .A3(\unit_decode/IMMreg/ffi_23/n4 ), 
        .ZN(n2373) );
  NAND2_X1 U2351 ( .A1(n2646), .A2(n2617), .ZN(n2377) );
  NOR3_X1 U2352 ( .A1(n2366), .A2(n2365), .A3(n2364), .ZN(n2378) );
  OAI22_X1 U2353 ( .A1(n1535), .A2(n2515), .B1(n2381), .B2(n2545), .ZN(n2364)
         );
  OAI22_X1 U2354 ( .A1(n2410), .A2(n2558), .B1(n2363), .B2(n2774), .ZN(n2365)
         );
  OAI211_X1 U2355 ( .C1(n2468), .C2(n2528), .A(n2362), .B(n2361), .ZN(n2366)
         );
  AOI22_X1 U2356 ( .A1(n1577), .A2(n2464), .B1(n2463), .B2(n2592), .ZN(n2361)
         );
  AOI22_X1 U2357 ( .A1(n2405), .A2(n2596), .B1(n2593), .B2(n2393), .ZN(n2362)
         );
  OAI21_X1 U2358 ( .B1(\unit_fetch/unit_npcregister/ffi_24/n4 ), .B2(n1921), 
        .A(n2663), .ZN(\unit_fetch/unit_npcregister/ffi_24/n5 ) );
  AOI22_X1 U2359 ( .A1(n1930), .A2(n2693), .B1(n1926), .B2(
        \unit_fetch/adder_out[24] ), .ZN(n2663) );
  OAI211_X1 U2360 ( .C1(n2360), .C2(n2780), .A(n2359), .B(n2358), .ZN(n2693)
         );
  AOI211_X1 U2361 ( .C1(n2606), .C2(n2404), .A(n2357), .B(n2356), .ZN(n2358)
         );
  OAI22_X1 U2362 ( .A1(n2410), .A2(n2450), .B1(n2448), .B2(n2438), .ZN(n2356)
         );
  OAI21_X1 U2363 ( .B1(n2355), .B2(n2608), .A(n2354), .ZN(n2357) );
  NAND2_X1 U2364 ( .A1(n1371), .A2(n2617), .ZN(n2359) );
  AOI211_X1 U2365 ( .C1(n2592), .C2(n2442), .A(n2351), .B(n2350), .ZN(n2360)
         );
  OAI22_X1 U2366 ( .A1(n2349), .A2(n2505), .B1(n2363), .B2(n2545), .ZN(n2350)
         );
  OAI22_X1 U2367 ( .A1(n2348), .A2(n2548), .B1(n2381), .B2(n2550), .ZN(n2351)
         );
  OAI21_X1 U2368 ( .B1(\unit_fetch/unit_npcregister/ffi_21/n4 ), .B2(n1921), 
        .A(n2666), .ZN(\unit_fetch/unit_npcregister/ffi_21/n5 ) );
  AOI22_X1 U2369 ( .A1(n1930), .A2(n2696), .B1(n1928), .B2(
        \unit_fetch/adder_out[21] ), .ZN(n2666) );
  OAI211_X1 U2370 ( .C1(n1361), .C2(n2544), .A(n2403), .B(n2402), .ZN(n2696)
         );
  OAI21_X1 U2371 ( .B1(n2401), .B2(n2400), .A(n2622), .ZN(n2402) );
  NAND2_X1 U2372 ( .A1(n2399), .A2(n2398), .ZN(n2400) );
  AOI22_X1 U2373 ( .A1(n2535), .A2(n2464), .B1(n2463), .B2(n1577), .ZN(n2398)
         );
  AOI22_X1 U2374 ( .A1(n2593), .A2(n2397), .B1(n2404), .B2(n2596), .ZN(n2399)
         );
  OAI211_X1 U2375 ( .C1(n2468), .C2(n2515), .A(n2396), .B(n2395), .ZN(n2401)
         );
  AOI22_X1 U2376 ( .A1(n2592), .A2(n2406), .B1(n2394), .B2(n2554), .ZN(n2395)
         );
  AOI22_X1 U2377 ( .A1(n2405), .A2(n2598), .B1(n2772), .B2(n2393), .ZN(n2396)
         );
  NAND2_X1 U2378 ( .A1(n2570), .A2(n1682), .ZN(n2392) );
  OAI21_X1 U2379 ( .B1(\unit_fetch/unit_npcregister/ffi_5/n4 ), .B2(n1921), 
        .A(n2682), .ZN(\unit_fetch/unit_npcregister/ffi_5/n5 ) );
  OAI21_X1 U2380 ( .B1(\unit_fetch/unit_npcregister/ffi_6/n4 ), .B2(n1921), 
        .A(n2681), .ZN(\unit_fetch/unit_npcregister/ffi_6/n5 ) );
  OAI21_X1 U2381 ( .B1(\unit_fetch/unit_npcregister/ffi_3/n4 ), .B2(n1921), 
        .A(n2684), .ZN(\unit_fetch/unit_npcregister/ffi_3/n5 ) );
  OAI21_X1 U2382 ( .B1(\unit_fetch/unit_npcregister/ffi_4/n4 ), .B2(n1921), 
        .A(n2683), .ZN(\unit_fetch/unit_npcregister/ffi_4/n5 ) );
  OAI21_X1 U2383 ( .B1(\unit_fetch/unit_programCounter/ffi_6/n4 ), .B2(n1922), 
        .A(n2681), .ZN(\unit_fetch/unit_programCounter/ffi_6/n5 ) );
  OAI211_X1 U2384 ( .C1(n2018), .C2(n2780), .A(n2017), .B(n2016), .ZN(n2918)
         );
  NAND2_X1 U2385 ( .A1(n2636), .A2(n2617), .ZN(n2017) );
  NOR3_X1 U2386 ( .A1(n2004), .A2(n2003), .A3(n2002), .ZN(n2018) );
  OAI22_X1 U2387 ( .A1(n2774), .A2(n2760), .B1(n2757), .B2(n2545), .ZN(n2002)
         );
  OAI22_X1 U2388 ( .A1(n2547), .A2(n2550), .B1(n2546), .B2(n2548), .ZN(n2003)
         );
  OAI211_X1 U2389 ( .C1(n2549), .C2(n2515), .A(n2001), .B(n2000), .ZN(n2004)
         );
  AOI22_X1 U2390 ( .A1(n2554), .A2(n2597), .B1(n2594), .B2(n2592), .ZN(n2000)
         );
  AOI22_X1 U2391 ( .A1(n2537), .A2(n2535), .B1(n1577), .B2(n2534), .ZN(n2001)
         );
  OAI21_X1 U2392 ( .B1(\unit_fetch/unit_programCounter/ffi_3/n4 ), .B2(n1922), 
        .A(n2684), .ZN(\unit_fetch/unit_programCounter/ffi_3/n5 ) );
  AOI22_X1 U2393 ( .A1(n2594), .A2(n2555), .B1(n2554), .B2(n2553), .ZN(n1983)
         );
  INV_X1 U2394 ( .A(n2595), .ZN(n1984) );
  OAI21_X1 U2395 ( .B1(\unit_fetch/unit_programCounter/ffi_27/n4 ), .B2(n1924), 
        .A(n2660), .ZN(\unit_fetch/unit_programCounter/ffi_27/n5 ) );
  OAI21_X1 U2396 ( .B1(\unit_fetch/unit_programCounter/ffi_5/n4 ), .B2(n1922), 
        .A(n2682), .ZN(\unit_fetch/unit_programCounter/ffi_5/n5 ) );
  OAI211_X1 U2397 ( .C1(n2601), .C2(n2515), .A(n1997), .B(n1996), .ZN(n1998)
         );
  NAND2_X1 U2398 ( .A1(n2554), .A2(n2594), .ZN(n1996) );
  AOI22_X1 U2399 ( .A1(n2592), .A2(n2595), .B1(n2597), .B2(n1577), .ZN(n1997)
         );
  AOI22_X1 U2400 ( .A1(n2536), .A2(n2598), .B1(n2593), .B2(n2533), .ZN(n1999)
         );
  OAI21_X1 U2401 ( .B1(\unit_fetch/unit_programCounter/ffi_4/n4 ), .B2(n1922), 
        .A(n2683), .ZN(\unit_fetch/unit_programCounter/ffi_4/n5 ) );
  OAI211_X1 U2402 ( .C1(n2579), .C2(n2780), .A(n2578), .B(n2577), .ZN(n2706)
         );
  AOI22_X1 U2403 ( .A1(n2573), .A2(n1652), .B1(n2572), .B2(n2571), .ZN(n2575)
         );
  NAND2_X1 U2404 ( .A1(n2570), .A2(n1652), .ZN(n2576) );
  NAND2_X1 U2405 ( .A1(n2629), .A2(n2617), .ZN(n2578) );
  NOR3_X1 U2406 ( .A1(n2561), .A2(n2560), .A3(n2559), .ZN(n2579) );
  OAI211_X1 U2407 ( .C1(n2601), .C2(n2558), .A(n2557), .B(n2556), .ZN(n2559)
         );
  AOI22_X1 U2408 ( .A1(n2597), .A2(n2555), .B1(n2554), .B2(n2595), .ZN(n2556)
         );
  AOI22_X1 U2409 ( .A1(n2553), .A2(n2592), .B1(n2594), .B2(n1577), .ZN(n2557)
         );
  INV_X1 U2410 ( .A(n2609), .ZN(n2553) );
  OAI22_X1 U2411 ( .A1(n2551), .A2(n2550), .B1(n2549), .B2(n2548), .ZN(n2560)
         );
  OAI22_X1 U2412 ( .A1(n2547), .A2(n2774), .B1(n2546), .B2(n2545), .ZN(n2561)
         );
  OAI21_X1 U2413 ( .B1(\unit_fetch/unit_programCounter/ffi_28/n4 ), .B2(n1924), 
        .A(n2659), .ZN(\unit_fetch/unit_programCounter/ffi_28/n5 ) );
  OAI21_X1 U2414 ( .B1(\unit_fetch/unit_programCounter/ffi_26/n4 ), .B2(n1924), 
        .A(n2661), .ZN(\unit_fetch/unit_programCounter/ffi_26/n5 ) );
  OAI21_X1 U2415 ( .B1(\unit_fetch/unit_npcregister/ffi_25/n4 ), .B2(n1921), 
        .A(n2662), .ZN(\unit_fetch/unit_npcregister/ffi_25/n5 ) );
  OAI21_X1 U2416 ( .B1(n2347), .B2(n2544), .A(n2346), .ZN(n2692) );
  AOI21_X1 U2417 ( .B1(n2622), .B2(n2345), .A(n2344), .ZN(n2346) );
  OAI211_X1 U2418 ( .C1(n2410), .C2(n2449), .A(n2343), .B(n2342), .ZN(n2344)
         );
  AOI21_X1 U2419 ( .B1(n2393), .B2(n1740), .A(n2341), .ZN(n2342) );
  OAI21_X1 U2420 ( .B1(n2340), .B2(n2339), .A(n2338), .ZN(n2341) );
  AOI22_X1 U2421 ( .A1(n2405), .A2(n2602), .B1(n2604), .B2(n2404), .ZN(n2343)
         );
  INV_X1 U2422 ( .A(n2355), .ZN(n2405) );
  INV_X1 U2423 ( .A(n2397), .ZN(n2410) );
  OAI211_X1 U2424 ( .C1(n2363), .C2(n2550), .A(n2337), .B(n2336), .ZN(n2345)
         );
  AOI22_X1 U2425 ( .A1(n2335), .A2(n2772), .B1(n2592), .B2(n2464), .ZN(n2336)
         );
  AOI22_X1 U2426 ( .A1(n1537), .A2(n2598), .B1(n2596), .B2(n2334), .ZN(n2337)
         );
  INV_X1 U2427 ( .A(n1566), .ZN(n2347) );
  OAI21_X1 U2428 ( .B1(\unit_fetch/unit_programCounter/ffi_7/n4 ), .B2(n1922), 
        .A(n2680), .ZN(\unit_fetch/unit_programCounter/ffi_7/n5 ) );
  AOI22_X1 U2429 ( .A1(n1931), .A2(n2919), .B1(n1927), .B2(
        \unit_fetch/adder_out[7] ), .ZN(n2680) );
  OAI21_X1 U2430 ( .B1(n2039), .B2(n2544), .A(n2038), .ZN(n2919) );
  AOI21_X1 U2431 ( .B1(n2037), .B2(n2622), .A(n2036), .ZN(n2038) );
  NOR2_X1 U2432 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_7/n4 ), .ZN(n2035)
         );
  AOI22_X1 U2433 ( .A1(n2535), .A2(n2533), .B1(n2122), .B2(n2772), .ZN(n2031)
         );
  AOI22_X1 U2434 ( .A1(n2537), .A2(n2555), .B1(n1577), .B2(n2027), .ZN(n2032)
         );
  INV_X1 U2435 ( .A(n2549), .ZN(n2027) );
  AOI211_X1 U2436 ( .C1(n2598), .C2(n2532), .A(n2026), .B(n2025), .ZN(n2033)
         );
  OAI22_X1 U2437 ( .A1(n2547), .A2(n2548), .B1(n2757), .B2(n2550), .ZN(n2025)
         );
  OAI22_X1 U2438 ( .A1(n2601), .A2(n2528), .B1(n2024), .B2(n2777), .ZN(n2026)
         );
  INV_X1 U2439 ( .A(n2597), .ZN(n2024) );
  INV_X1 U2440 ( .A(n1389), .ZN(n2039) );
  OAI21_X1 U2441 ( .B1(\unit_fetch/unit_programCounter/ffi_17/n4 ), .B2(n1923), 
        .A(n2670), .ZN(\unit_fetch/unit_programCounter/ffi_17/n5 ) );
  OAI21_X1 U2442 ( .B1(\unit_fetch/unit_programCounter/ffi_18/n4 ), .B2(n1923), 
        .A(n2669), .ZN(\unit_fetch/unit_programCounter/ffi_18/n5 ) );
  OAI21_X1 U2443 ( .B1(\unit_fetch/unit_programCounter/ffi_11/n4 ), .B2(n1923), 
        .A(n2676), .ZN(\unit_fetch/unit_programCounter/ffi_11/n5 ) );
  OAI21_X1 U2444 ( .B1(\unit_fetch/unit_adder/add_19/n47 ), .B2(n1923), .A(
        n2674), .ZN(\unit_fetch/unit_programCounter/ffi_13/n5 ) );
  OAI21_X1 U2445 ( .B1(\unit_fetch/unit_npcregister/ffi_28/n4 ), .B2(n1922), 
        .A(n2659), .ZN(\unit_fetch/unit_npcregister/ffi_28/n5 ) );
  OAI21_X1 U2446 ( .B1(n2297), .B2(n2296), .A(n2622), .ZN(n2298) );
  OAI22_X1 U2447 ( .A1(n2313), .A2(n2545), .B1(n2355), .B2(n2777), .ZN(n2296)
         );
  OAI21_X1 U2448 ( .B1(n2774), .B2(n2285), .A(n2284), .ZN(n2297) );
  AOI22_X1 U2449 ( .A1(n2593), .A2(n2283), .B1(n2335), .B2(n2596), .ZN(n2284)
         );
  INV_X1 U2450 ( .A(n2323), .ZN(n2283) );
  AOI211_X1 U2451 ( .C1(n2606), .C2(n2334), .A(n2281), .B(n2280), .ZN(n2299)
         );
  OAI22_X1 U2452 ( .A1(n2348), .A2(n2448), .B1(n2450), .B2(n2363), .ZN(n2280)
         );
  INV_X1 U2453 ( .A(n2393), .ZN(n2348) );
  OAI21_X1 U2454 ( .B1(n2349), .B2(n2608), .A(n2279), .ZN(n2281) );
  AOI21_X1 U2455 ( .B1(n2326), .B2(n2278), .A(n2277), .ZN(n2279) );
  NOR3_X1 U2456 ( .A1(n2779), .A2(n2278), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2277) );
  OAI21_X1 U2457 ( .B1(\unit_fetch/unit_npcregister/ffi_27/n4 ), .B2(n1921), 
        .A(n2660), .ZN(\unit_fetch/unit_npcregister/ffi_27/n5 ) );
  OAI211_X1 U2458 ( .C1(n2648), .C2(n2544), .A(n2317), .B(n2316), .ZN(n2690)
         );
  OAI21_X1 U2459 ( .B1(n2315), .B2(n2314), .A(n2622), .ZN(n2316) );
  OAI22_X1 U2460 ( .A1(n2774), .A2(n2313), .B1(n2349), .B2(n2548), .ZN(n2314)
         );
  OAI21_X1 U2461 ( .B1(n2323), .B2(n2545), .A(n2312), .ZN(n2315) );
  AOI22_X1 U2462 ( .A1(n2335), .A2(n2593), .B1(n2592), .B2(n2397), .ZN(n2312)
         );
  AOI211_X1 U2463 ( .C1(n2606), .C2(n2393), .A(n2311), .B(n2310), .ZN(n2317)
         );
  OAI22_X1 U2464 ( .A1(n2355), .A2(n2448), .B1(n2450), .B2(n2381), .ZN(n2310)
         );
  OAI21_X1 U2465 ( .B1(n2363), .B2(n2608), .A(n2309), .ZN(n2311) );
  AOI21_X1 U2466 ( .B1(n2308), .B2(n2307), .A(n2306), .ZN(n2309) );
  NOR3_X1 U2467 ( .A1(n2779), .A2(n2307), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2306) );
  OAI21_X1 U2468 ( .B1(\unit_fetch/unit_npcregister/ffi_26/n4 ), .B2(n1921), 
        .A(n2661), .ZN(\unit_fetch/unit_npcregister/ffi_26/n5 ) );
  OAI21_X1 U2469 ( .B1(n2647), .B2(n2544), .A(n2332), .ZN(n2691) );
  AOI21_X1 U2470 ( .B1(n2622), .B2(n2331), .A(n2330), .ZN(n2332) );
  OAI211_X1 U2471 ( .C1(n2355), .C2(n2449), .A(n2329), .B(n2328), .ZN(n2330)
         );
  AOI22_X1 U2472 ( .A1(n2604), .A2(n2397), .B1(n2602), .B2(n2393), .ZN(n2328)
         );
  AOI211_X1 U2473 ( .C1(n2327), .C2(n2326), .A(n2325), .B(n2324), .ZN(n2329)
         );
  AND2_X1 U2474 ( .A1(n2334), .A2(n1740), .ZN(n2324) );
  NOR3_X1 U2475 ( .A1(n2779), .A2(n2327), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2325) );
  AND3_X1 U2476 ( .A1(n2295), .A2(n2294), .A3(n2293), .ZN(n2355) );
  INV_X1 U2477 ( .A(n2292), .ZN(n2293) );
  OAI22_X1 U2478 ( .A1(n2291), .A2(n1549), .B1(n1582), .B2(n1918), .ZN(n2292)
         );
  AOI22_X1 U2479 ( .A1(n2288), .A2(n2287), .B1(n2286), .B2(n2775), .ZN(n2295)
         );
  OAI211_X1 U2480 ( .C1(n2774), .C2(n2323), .A(n2322), .B(n2321), .ZN(n2331)
         );
  AOI22_X1 U2481 ( .A1(n2335), .A2(n2598), .B1(n2592), .B2(n2404), .ZN(n2321)
         );
  INV_X1 U2482 ( .A(n2282), .ZN(n2335) );
  AOI22_X1 U2483 ( .A1(n1537), .A2(n2593), .B1(n2596), .B2(n2320), .ZN(n2322)
         );
  OAI21_X1 U2484 ( .B1(\unit_fetch/unit_npcregister/ffi_9/n4 ), .B2(n1921), 
        .A(n2678), .ZN(\unit_fetch/unit_npcregister/ffi_9/n5 ) );
  OAI21_X1 U2485 ( .B1(\unit_fetch/unit_npcregister/ffi_11/n4 ), .B2(n1921), 
        .A(n2676), .ZN(\unit_fetch/unit_npcregister/ffi_11/n5 ) );
  AOI22_X1 U2486 ( .A1(n1931), .A2(n2703), .B1(n1928), .B2(
        \unit_fetch/adder_out[11] ), .ZN(n2676) );
  AOI22_X1 U2487 ( .A1(n2596), .A2(n2511), .B1(n2508), .B2(n1577), .ZN(n1725)
         );
  NOR2_X1 U2488 ( .A1(n1728), .A2(n1727), .ZN(n1726) );
  NOR2_X1 U2489 ( .A1(n2505), .A2(n2506), .ZN(n1727) );
  OAI21_X1 U2490 ( .B1(n2529), .B2(n2558), .A(n1729), .ZN(n1728) );
  AOI21_X1 U2491 ( .B1(n1732), .B2(n1731), .A(n1730), .ZN(n1729) );
  NOR2_X1 U2492 ( .A1(n2760), .A2(n2515), .ZN(n1730) );
  INV_X1 U2493 ( .A(n2545), .ZN(n1731) );
  AOI22_X1 U2494 ( .A1(n2536), .A2(n2554), .B1(n2592), .B2(n2533), .ZN(n2509)
         );
  OAI21_X1 U2495 ( .B1(\unit_fetch/unit_programCounter/ffi_15/n4 ), .B2(n1923), 
        .A(n2672), .ZN(\unit_fetch/unit_programCounter/ffi_15/n5 ) );
  OAI21_X1 U2496 ( .B1(\unit_fetch/unit_programCounter/ffi_9/n4 ), .B2(n1922), 
        .A(n2678), .ZN(\unit_fetch/unit_programCounter/ffi_9/n5 ) );
  AOI22_X1 U2497 ( .A1(n1930), .A2(n2920), .B1(n1926), .B2(
        \unit_fetch/adder_out[9] ), .ZN(n2678) );
  OAI211_X1 U2498 ( .C1(n2066), .C2(n2780), .A(n2065), .B(n2064), .ZN(n2920)
         );
  AOI211_X1 U2499 ( .C1(n1740), .C2(n2508), .A(n2063), .B(n2062), .ZN(n2064)
         );
  OAI22_X1 U2500 ( .A1(n2547), .A2(n2450), .B1(n2546), .B2(n2449), .ZN(n2062)
         );
  INV_X1 U2501 ( .A(n2533), .ZN(n2546) );
  OAI21_X1 U2502 ( .B1(n2551), .B2(n2448), .A(n2061), .ZN(n2063) );
  NAND2_X1 U2503 ( .A1(n2570), .A2(n1684), .ZN(n2059) );
  INV_X1 U2504 ( .A(n2757), .ZN(n2508) );
  NAND2_X1 U2505 ( .A1(n1391), .A2(n2617), .ZN(n2065) );
  AOI211_X1 U2506 ( .C1(n2596), .C2(n2532), .A(n2044), .B(n2043), .ZN(n2066)
         );
  OAI22_X1 U2507 ( .A1(n2529), .A2(n2550), .B1(n2549), .B2(n2777), .ZN(n2043)
         );
  OAI22_X1 U2508 ( .A1(n2774), .A2(n2514), .B1(n2527), .B2(n2545), .ZN(n2044)
         );
  OAI21_X1 U2509 ( .B1(\unit_fetch/unit_npcregister/ffi_13/n4 ), .B2(n1922), 
        .A(n2674), .ZN(\unit_fetch/unit_npcregister/ffi_13/n5 ) );
  AOI22_X1 U2510 ( .A1(n1931), .A2(n2913), .B1(n1926), .B2(
        \unit_fetch/adder_out[13] ), .ZN(n2674) );
  NAND2_X1 U2511 ( .A1(n2511), .A2(n2602), .ZN(n1843) );
  NAND2_X1 U2512 ( .A1(n2532), .A2(n2604), .ZN(n1844) );
  NAND2_X1 U2513 ( .A1(n2570), .A2(n1672), .ZN(n2099) );
  AOI22_X1 U2514 ( .A1(n2598), .A2(n2407), .B1(n2596), .B2(n2512), .ZN(n2756)
         );
  OAI21_X1 U2515 ( .B1(\unit_fetch/unit_npcregister/ffi_18/n4 ), .B2(n1921), 
        .A(n2669), .ZN(\unit_fetch/unit_npcregister/ffi_18/n5 ) );
  AOI22_X1 U2516 ( .A1(n1930), .A2(n2699), .B1(n1928), .B2(
        \unit_fetch/adder_out[18] ), .ZN(n2669) );
  OAI211_X1 U2517 ( .C1(n2459), .C2(n2780), .A(n2458), .B(n2457), .ZN(n2699)
         );
  NOR3_X1 U2518 ( .A1(n2456), .A2(n2455), .A3(n2454), .ZN(n2457) );
  NOR2_X1 U2519 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_18/n4 ), .ZN(n2453)
         );
  OAI22_X1 U2520 ( .A1(n2450), .A2(n2461), .B1(n2460), .B2(n2449), .ZN(n2455)
         );
  INV_X1 U2521 ( .A(n2606), .ZN(n2449) );
  OAI22_X1 U2522 ( .A1(n2506), .A2(n2448), .B1(n2462), .B2(n2608), .ZN(n2456)
         );
  NAND2_X1 U2523 ( .A1(n2640), .A2(n2617), .ZN(n2458) );
  AOI211_X1 U2524 ( .C1(n2593), .C2(n2442), .A(n2441), .B(n2440), .ZN(n2459)
         );
  OAI22_X1 U2525 ( .A1(n2507), .A2(n2777), .B1(n2439), .B2(n2548), .ZN(n2440)
         );
  OAI22_X1 U2526 ( .A1(n1535), .A2(n2505), .B1(n2438), .B2(n2545), .ZN(n2441)
         );
  OAI21_X1 U2527 ( .B1(\unit_fetch/unit_npcregister/ffi_17/n4 ), .B2(n1921), 
        .A(n2670), .ZN(\unit_fetch/unit_npcregister/ffi_17/n5 ) );
  AOI22_X1 U2528 ( .A1(n1930), .A2(n2700), .B1(n1928), .B2(
        \unit_fetch/adder_out[17] ), .ZN(n2670) );
  OAI211_X1 U2529 ( .C1(n2479), .C2(n2780), .A(n2478), .B(n2477), .ZN(n2700)
         );
  NAND2_X1 U2530 ( .A1(n2570), .A2(n1666), .ZN(n2475) );
  NAND2_X1 U2531 ( .A1(n2642), .A2(n2617), .ZN(n2478) );
  NOR3_X1 U2532 ( .A1(n2471), .A2(n2470), .A3(n2469), .ZN(n2479) );
  OAI211_X1 U2533 ( .C1(n2468), .C2(n2545), .A(n2467), .B(n2466), .ZN(n2469)
         );
  AOI22_X1 U2534 ( .A1(n2592), .A2(n2504), .B1(n2465), .B2(n1577), .ZN(n2466)
         );
  AOI22_X1 U2535 ( .A1(n2772), .A2(n2464), .B1(n2463), .B2(n2593), .ZN(n2467)
         );
  INV_X1 U2536 ( .A(n2442), .ZN(n2468) );
  OAI22_X1 U2537 ( .A1(n2462), .A2(n2548), .B1(n2461), .B2(n2558), .ZN(n2470)
         );
  INV_X1 U2538 ( .A(n2406), .ZN(n2461) );
  OAI22_X1 U2539 ( .A1(n2507), .A2(n2528), .B1(n2460), .B2(n2515), .ZN(n2471)
         );
  OAI21_X1 U2540 ( .B1(\unit_fetch/unit_npcregister/ffi_16/n4 ), .B2(n1921), 
        .A(n2671), .ZN(\unit_fetch/unit_npcregister/ffi_16/n5 ) );
  AOI22_X1 U2541 ( .A1(n1930), .A2(n2701), .B1(n1928), .B2(
        \unit_fetch/adder_out[16] ), .ZN(n2671) );
  OAI21_X1 U2542 ( .B1(n2483), .B2(n2544), .A(n2482), .ZN(n2701) );
  AOI21_X1 U2543 ( .B1(n1749), .B2(n2622), .A(n1748), .ZN(n2482) );
  OR2_X1 U2544 ( .A1(n2481), .A2(n2768), .ZN(n1748) );
  NOR3_X1 U2545 ( .A1(n1580), .A2(n2611), .A3(n1668), .ZN(n2481) );
  NOR3_X1 U2546 ( .A1(n1754), .A2(n1753), .A3(n1751), .ZN(n1750) );
  OAI21_X1 U2547 ( .B1(n2514), .B2(n2528), .A(n1752), .ZN(n1751) );
  NAND2_X1 U2548 ( .A1(n2442), .A2(n2772), .ZN(n1752) );
  NOR2_X1 U2549 ( .A1(n2527), .A2(n2777), .ZN(n1753) );
  OAI22_X1 U2550 ( .A1(n2462), .A2(n2550), .B1(n2439), .B2(n2545), .ZN(n1754)
         );
  AOI22_X1 U2551 ( .A1(n2596), .A2(n2406), .B1(n2535), .B2(n2407), .ZN(n2766)
         );
  AOI22_X1 U2552 ( .A1(n2555), .A2(n2465), .B1(n1577), .B2(n2512), .ZN(n2765)
         );
  INV_X1 U2553 ( .A(n1550), .ZN(n2483) );
  OAI21_X1 U2554 ( .B1(\unit_fetch/unit_programCounter/ffi_14/n4 ), .B2(n1923), 
        .A(n2673), .ZN(\unit_fetch/unit_programCounter/ffi_14/n5 ) );
  OAI21_X1 U2555 ( .B1(\unit_fetch/unit_programCounter/ffi_29/n4 ), .B2(n1924), 
        .A(n2658), .ZN(\unit_fetch/unit_programCounter/ffi_29/n5 ) );
  OAI21_X1 U2556 ( .B1(\unit_fetch/unit_npcregister/ffi_15/n4 ), .B2(n1921), 
        .A(n2672), .ZN(\unit_fetch/unit_npcregister/ffi_15/n5 ) );
  AOI22_X1 U2557 ( .A1(n1930), .A2(n2702), .B1(n1928), .B2(
        \unit_fetch/adder_out[15] ), .ZN(n2672) );
  OAI21_X1 U2558 ( .B1(n1657), .B2(n2544), .A(n2492), .ZN(n2702) );
  AOI21_X1 U2559 ( .B1(n2622), .B2(n2764), .A(n2491), .ZN(n2492) );
  NOR2_X1 U2560 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_15/n4 ), .ZN(n2490)
         );
  NOR2_X1 U2561 ( .A1(n2121), .A2(n1741), .ZN(n2761) );
  NAND2_X1 U2562 ( .A1(n1747), .A2(n1742), .ZN(n1741) );
  AOI22_X1 U2563 ( .A1(n2406), .A2(n2593), .B1(n2463), .B2(n2772), .ZN(n1742)
         );
  NAND2_X1 U2564 ( .A1(n2122), .A2(n2592), .ZN(n1747) );
  OAI22_X1 U2565 ( .A1(n2514), .A2(n2552), .B1(n2527), .B2(n2528), .ZN(n2121)
         );
  AOI22_X1 U2566 ( .A1(n2555), .A2(n2512), .B1(n2535), .B2(n2465), .ZN(n2762)
         );
  INV_X1 U2567 ( .A(n2507), .ZN(n2512) );
  AOI22_X1 U2568 ( .A1(n2598), .A2(n2394), .B1(n2596), .B2(n2407), .ZN(n2763)
         );
  OAI21_X1 U2569 ( .B1(\unit_fetch/unit_npcregister/ffi_14/n4 ), .B2(n1921), 
        .A(n2673), .ZN(\unit_fetch/unit_npcregister/ffi_14/n5 ) );
  AOI22_X1 U2570 ( .A1(n1931), .A2(n2914), .B1(n1928), .B2(
        \unit_fetch/adder_out[14] ), .ZN(n2673) );
  OAI21_X1 U2571 ( .B1(n2637), .B2(n2544), .A(n2116), .ZN(n2914) );
  AOI21_X1 U2572 ( .B1(n1822), .B2(n2622), .A(n1817), .ZN(n2116) );
  NAND2_X1 U2573 ( .A1(n2114), .A2(n1686), .ZN(n1817) );
  NAND2_X1 U2574 ( .A1(n2122), .A2(n2604), .ZN(n1818) );
  NOR2_X1 U2575 ( .A1(n2115), .A2(n1820), .ZN(n1819) );
  NOR2_X1 U2576 ( .A1(n2507), .A2(n2608), .ZN(n1820) );
  NOR2_X1 U2577 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_14/n4 ), .ZN(n2113)
         );
  NAND2_X1 U2578 ( .A1(n2504), .A2(n2602), .ZN(n1821) );
  NAND2_X1 U2579 ( .A1(n2511), .A2(n2606), .ZN(n2114) );
  NAND2_X1 U2580 ( .A1(n2758), .A2(n1823), .ZN(n1822) );
  NOR2_X1 U2581 ( .A1(n1825), .A2(n1824), .ZN(n1823) );
  NOR2_X1 U2582 ( .A1(n2760), .A2(n2777), .ZN(n1824) );
  INV_X1 U2583 ( .A(n2759), .ZN(n1825) );
  AOI22_X1 U2584 ( .A1(n2598), .A2(n2406), .B1(n2596), .B2(n2465), .ZN(n2759)
         );
  AOI22_X1 U2585 ( .A1(n2593), .A2(n2407), .B1(n2772), .B2(n2394), .ZN(n2758)
         );
  OAI21_X1 U2586 ( .B1(\unit_fetch/unit_npcregister/ffi_29/n4 ), .B2(n1922), 
        .A(n2658), .ZN(\unit_fetch/unit_npcregister/ffi_29/n5 ) );
  OAI211_X1 U2587 ( .C1(n2274), .C2(n2780), .A(n2273), .B(n2272), .ZN(n2688)
         );
  AOI211_X1 U2588 ( .C1(n2606), .C2(n2320), .A(n2271), .B(n2270), .ZN(n2272)
         );
  OAI22_X1 U2589 ( .A1(n2349), .A2(n2450), .B1(n2448), .B2(n2381), .ZN(n2270)
         );
  INV_X1 U2590 ( .A(n2334), .ZN(n2381) );
  INV_X1 U2591 ( .A(n2604), .ZN(n2448) );
  INV_X1 U2592 ( .A(n2602), .ZN(n2450) );
  OAI21_X1 U2593 ( .B1(n2282), .B2(n2608), .A(n2269), .ZN(n2271) );
  AOI21_X1 U2594 ( .B1(n2268), .B2(n2267), .A(n2266), .ZN(n2269) );
  NOR3_X1 U2595 ( .A1(n2779), .A2(n2267), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2266) );
  OAI21_X1 U2596 ( .B1(n2611), .B2(n1660), .A(n2265), .ZN(n2268) );
  NAND2_X1 U2597 ( .A1(n2573), .A2(n1660), .ZN(n2265) );
  NAND2_X1 U2598 ( .A1(n2652), .A2(n2617), .ZN(n2273) );
  AOI211_X1 U2599 ( .C1(n2592), .C2(n2393), .A(n2259), .B(n2258), .ZN(n2274)
         );
  OAI22_X1 U2600 ( .A1(n2323), .A2(n2548), .B1(n2285), .B2(n2545), .ZN(n2258)
         );
  OAI22_X1 U2601 ( .A1(n2313), .A2(n2550), .B1(n2257), .B2(n2774), .ZN(n2259)
         );
  NAND4_X1 U2602 ( .A1(n2294), .A2(n2256), .A3(n2255), .A4(n2254), .ZN(n2393)
         );
  NAND2_X1 U2603 ( .A1(n2253), .A2(n2288), .ZN(n2254) );
  NAND2_X1 U2604 ( .A1(n2252), .A2(n2251), .ZN(n2255) );
  INV_X1 U2605 ( .A(n2250), .ZN(n2256) );
  OAI21_X1 U2606 ( .B1(\unit_fetch/unit_npcregister/ffi_8/n4 ), .B2(n1922), 
        .A(n2679), .ZN(\unit_fetch/unit_npcregister/ffi_8/n5 ) );
  OAI21_X1 U2607 ( .B1(\unit_fetch/unit_programCounter/ffi_8/n4 ), .B2(n1922), 
        .A(n2679), .ZN(\unit_fetch/unit_programCounter/ffi_8/n5 ) );
  AOI22_X1 U2608 ( .A1(n1931), .A2(n2705), .B1(n1926), .B2(
        \unit_fetch/adder_out[8] ), .ZN(n2679) );
  AOI22_X1 U2609 ( .A1(n1577), .A2(n2537), .B1(n2536), .B2(n2535), .ZN(n2538)
         );
  INV_X1 U2610 ( .A(n2547), .ZN(n2536) );
  INV_X1 U2611 ( .A(n2551), .ZN(n2537) );
  NOR2_X1 U2612 ( .A1(n1993), .A2(n1977), .ZN(n2551) );
  AOI22_X1 U2613 ( .A1(n2534), .A2(n2592), .B1(n2555), .B2(n2533), .ZN(n2539)
         );
  OAI211_X1 U2614 ( .C1(n2146), .C2(n2030), .A(n2029), .B(n1985), .ZN(n2533)
         );
  INV_X1 U2615 ( .A(n2515), .ZN(n2555) );
  INV_X1 U2616 ( .A(n2601), .ZN(n2534) );
  AOI211_X1 U2617 ( .C1(n2593), .C2(n2532), .A(n2531), .B(n2530), .ZN(n2540)
         );
  OAI22_X1 U2618 ( .A1(n2529), .A2(n2545), .B1(n2757), .B2(n2548), .ZN(n2530)
         );
  OAI22_X1 U2619 ( .A1(n2549), .A2(n2528), .B1(n2774), .B2(n2527), .ZN(n2531)
         );
  INV_X1 U2620 ( .A(n1947), .ZN(n1948) );
  INV_X1 U2621 ( .A(n2760), .ZN(n2532) );
  OAI21_X1 U2622 ( .B1(\unit_fetch/unit_programCounter/ffi_12/n4 ), .B2(n1923), 
        .A(n2675), .ZN(\unit_fetch/unit_programCounter/ffi_12/n5 ) );
  OAI21_X1 U2623 ( .B1(\unit_fetch/unit_npcregister/ffi_12/n4 ), .B2(n1924), 
        .A(n2675), .ZN(\unit_fetch/unit_npcregister/ffi_12/n5 ) );
  AOI22_X1 U2624 ( .A1(n1931), .A2(n2912), .B1(n1928), .B2(
        \unit_fetch/adder_out[12] ), .ZN(n2675) );
  OAI211_X1 U2625 ( .C1(n2089), .C2(n2544), .A(n2088), .B(n2087), .ZN(n2912)
         );
  NAND2_X1 U2626 ( .A1(n2570), .A2(n1663), .ZN(n2085) );
  OAI21_X1 U2627 ( .B1(n2084), .B2(n2083), .A(n2622), .ZN(n2088) );
  OAI21_X1 U2628 ( .B1(n2460), .B2(n2505), .A(n2755), .ZN(n2083) );
  OAI22_X1 U2629 ( .A1(n2760), .A2(n2552), .B1(n2757), .B2(n2528), .ZN(n2752)
         );
  INV_X1 U2630 ( .A(n1994), .ZN(n1995) );
  OAI22_X1 U2631 ( .A1(n2529), .A2(n2515), .B1(n2527), .B2(n2558), .ZN(n2753)
         );
  INV_X1 U2632 ( .A(n2511), .ZN(n2527) );
  NAND4_X1 U2633 ( .A1(n2120), .A2(n2042), .A3(n2041), .A4(n2040), .ZN(n2511)
         );
  NAND2_X1 U2634 ( .A1(n1546), .A2(n2175), .ZN(n2040) );
  NAND2_X1 U2635 ( .A1(n2612), .A2(n2775), .ZN(n2041) );
  NAND2_X1 U2636 ( .A1(n2711), .A2(n2571), .ZN(n2042) );
  INV_X1 U2637 ( .A(n2122), .ZN(n2529) );
  NAND2_X1 U2638 ( .A1(n2028), .A2(n1734), .ZN(n2122) );
  AND2_X1 U2639 ( .A1(n2029), .A2(n1735), .ZN(n1734) );
  NAND2_X1 U2640 ( .A1(n1737), .A2(n1736), .ZN(n1735) );
  INV_X1 U2641 ( .A(n2030), .ZN(n1737) );
  NAND2_X1 U2642 ( .A1(n1544), .A2(n2175), .ZN(n2028) );
  OAI22_X1 U2643 ( .A1(n2506), .A2(n2545), .B1(n2514), .B2(n2548), .ZN(n2754)
         );
  INV_X1 U2644 ( .A(n2504), .ZN(n2514) );
  INV_X1 U2645 ( .A(n2465), .ZN(n2506) );
  INV_X1 U2646 ( .A(n2772), .ZN(n2505) );
  OAI22_X1 U2647 ( .A1(n2507), .A2(n2550), .B1(n2547), .B2(n2777), .ZN(n2084)
         );
  NOR2_X1 U2648 ( .A1(n1993), .A2(n1992), .ZN(n2547) );
  OAI22_X1 U2649 ( .A1(n2162), .A2(n2030), .B1(n1549), .B2(n1918), .ZN(n1992)
         );
  INV_X1 U2650 ( .A(n2029), .ZN(n1993) );
  AND2_X1 U2651 ( .A1(n2082), .A2(n2571), .ZN(n1733) );
  INV_X1 U2652 ( .A(n2451), .ZN(n2082) );
  INV_X1 U2653 ( .A(n2120), .ZN(n2080) );
  INV_X1 U2654 ( .A(n2635), .ZN(n2089) );
  OAI211_X1 U2655 ( .C1(n2227), .C2(n2780), .A(n2226), .B(n2225), .ZN(n2686)
         );
  AOI21_X1 U2656 ( .B1(n2326), .B2(n1534), .A(n2224), .ZN(n2225) );
  NOR3_X1 U2657 ( .A1(n2779), .A2(n1534), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2224) );
  NAND2_X1 U2658 ( .A1(n2651), .A2(n2617), .ZN(n2226) );
  NOR4_X1 U2659 ( .A1(n2185), .A2(n2184), .A3(n2183), .A4(n2182), .ZN(n2227)
         );
  OAI211_X1 U2660 ( .C1(n2285), .C2(n2548), .A(n2181), .B(n2180), .ZN(n2182)
         );
  NAND2_X1 U2661 ( .A1(n2232), .A2(n2598), .ZN(n2180) );
  NAND4_X1 U2662 ( .A1(n2179), .A2(n2178), .A3(n2177), .A4(n2176), .ZN(n2232)
         );
  NAND2_X1 U2663 ( .A1(n2230), .A2(n2175), .ZN(n2176) );
  INV_X1 U2664 ( .A(n2244), .ZN(n2230) );
  INV_X1 U2665 ( .A(n2174), .ZN(n2177) );
  INV_X1 U2666 ( .A(n2173), .ZN(n2178) );
  OAI22_X1 U2667 ( .A1(n2291), .A2(n1554), .B1(n2388), .B2(n2248), .ZN(n2173)
         );
  OAI211_X1 U2668 ( .C1(n2170), .C2(n2169), .A(\unit_decode/IMMreg/ffi_0/n4 ), 
        .B(n1576), .ZN(n2181) );
  OAI22_X1 U2669 ( .A1(n2374), .A2(n2248), .B1(n2587), .B2(n1918), .ZN(n2169)
         );
  OAI22_X1 U2670 ( .A1(n2171), .A2(n1630), .B1(n2291), .B2(n2488), .ZN(n2170)
         );
  AND2_X1 U2671 ( .A1(n2167), .A2(n2166), .ZN(n2285) );
  AOI22_X1 U2672 ( .A1(n2165), .A2(n2164), .B1(n2287), .B2(n2175), .ZN(n2166)
         );
  INV_X1 U2673 ( .A(n2278), .ZN(n2287) );
  INV_X1 U2674 ( .A(n2171), .ZN(n2165) );
  NOR2_X1 U2675 ( .A1(n2163), .A2(n2174), .ZN(n2167) );
  OAI22_X1 U2676 ( .A1(n2291), .A2(n1370), .B1(n1582), .B2(n2248), .ZN(n2163)
         );
  OAI22_X1 U2677 ( .A1(n2349), .A2(n2528), .B1(n2257), .B2(n2550), .ZN(n2183)
         );
  OAI22_X1 U2678 ( .A1(n2291), .A2(n1589), .B1(n2353), .B2(n1918), .ZN(n2159)
         );
  OAI22_X1 U2679 ( .A1(n2323), .A2(n2515), .B1(n2363), .B2(n2777), .ZN(n2184)
         );
  INV_X1 U2680 ( .A(n2320), .ZN(n2363) );
  NOR3_X1 U2681 ( .A1(n2157), .A2(n2156), .A3(n2174), .ZN(n2323) );
  OAI22_X1 U2682 ( .A1(n2291), .A2(n2155), .B1(n1631), .B2(n2248), .ZN(n2156)
         );
  OAI22_X1 U2683 ( .A1(n2313), .A2(n2558), .B1(n2282), .B2(n2552), .ZN(n2185)
         );
  NOR3_X1 U2684 ( .A1(n2153), .A2(n2152), .A3(n2174), .ZN(n2282) );
  OAI21_X1 U2685 ( .B1(n2248), .B2(n1759), .A(n1697), .ZN(n2152) );
  NOR3_X1 U2686 ( .A1(n2149), .A2(n2148), .A3(n2174), .ZN(n2313) );
  OAI22_X1 U2687 ( .A1(n2307), .A2(n1919), .B1(n2432), .B2(n2773), .ZN(n2148)
         );
  NAND2_X1 U2688 ( .A1(n2145), .A2(n2144), .ZN(n2171) );
  NOR2_X1 U2689 ( .A1(n1661), .A2(n1567), .ZN(n2144) );
  INV_X1 U2690 ( .A(n2143), .ZN(n2145) );
  OAI21_X1 U2691 ( .B1(\unit_fetch/unit_programCounter/ffi_19/n4 ), .B2(n1923), 
        .A(n2668), .ZN(\unit_fetch/unit_programCounter/ffi_19/n5 ) );
  OAI21_X1 U2692 ( .B1(\unit_fetch/unit_npcregister/ffi_19/n4 ), .B2(n1921), 
        .A(n2668), .ZN(\unit_fetch/unit_npcregister/ffi_19/n5 ) );
  AOI22_X1 U2693 ( .A1(n1930), .A2(n2698), .B1(n1928), .B2(
        \unit_fetch/adder_out[19] ), .ZN(n2668) );
  OAI21_X1 U2694 ( .B1(n2437), .B2(n2544), .A(n2436), .ZN(n2698) );
  AOI21_X1 U2695 ( .B1(n2622), .B2(n2771), .A(n2435), .ZN(n2436) );
  NOR2_X1 U2696 ( .A1(n2779), .A2(\unit_decode/IMMreg/ffi_19/n4 ), .ZN(n2434)
         );
  OAI22_X1 U2697 ( .A1(n2439), .A2(n2558), .B1(n2462), .B2(n2515), .ZN(n2139)
         );
  INV_X1 U2698 ( .A(n2394), .ZN(n2462) );
  NAND4_X1 U2699 ( .A1(n2120), .A2(n2106), .A3(n2105), .A4(n2104), .ZN(n2394)
         );
  NAND2_X1 U2700 ( .A1(n2103), .A2(n2571), .ZN(n2104) );
  INV_X1 U2701 ( .A(n2388), .ZN(n2103) );
  NAND2_X1 U2702 ( .A1(n1618), .A2(n2775), .ZN(n2105) );
  NAND2_X1 U2703 ( .A1(n2102), .A2(n2175), .ZN(n2106) );
  INV_X1 U2704 ( .A(n1554), .ZN(n2102) );
  INV_X1 U2705 ( .A(n2535), .ZN(n2558) );
  INV_X1 U2706 ( .A(n2463), .ZN(n2439) );
  NAND2_X1 U2707 ( .A1(n2119), .A2(n1743), .ZN(n2463) );
  NOR2_X1 U2708 ( .A1(n1691), .A2(n1744), .ZN(n1743) );
  NAND2_X1 U2709 ( .A1(n2120), .A2(n2118), .ZN(n1744) );
  NAND2_X1 U2710 ( .A1(n2117), .A2(n2571), .ZN(n2118) );
  INV_X1 U2711 ( .A(n2374), .ZN(n2117) );
  NAND2_X1 U2712 ( .A1(n1544), .A2(n2775), .ZN(n2119) );
  OAI22_X1 U2713 ( .A1(n1535), .A2(n2545), .B1(n2438), .B2(n2550), .ZN(n2140)
         );
  INV_X1 U2714 ( .A(n2464), .ZN(n2438) );
  NAND4_X1 U2715 ( .A1(n2138), .A2(n2294), .A3(n2137), .A4(n2136), .ZN(n2464)
         );
  NAND2_X1 U2716 ( .A1(n2339), .A2(n2288), .ZN(n2136) );
  INV_X1 U2717 ( .A(n2209), .ZN(n2339) );
  NAND2_X1 U2718 ( .A1(n2135), .A2(n2775), .ZN(n2137) );
  INV_X1 U2719 ( .A(n2134), .ZN(n2138) );
  NAND2_X1 U2720 ( .A1(n1797), .A2(n2288), .ZN(n2131) );
  NAND2_X1 U2721 ( .A1(n2522), .A2(n2775), .ZN(n2132) );
  INV_X1 U2722 ( .A(n2130), .ZN(n2133) );
  AOI22_X1 U2723 ( .A1(n2596), .A2(n2442), .B1(n2772), .B2(n2397), .ZN(n2769)
         );
  NAND4_X1 U2724 ( .A1(n2129), .A2(n2294), .A3(n2128), .A4(n2127), .ZN(n2397)
         );
  NAND2_X1 U2725 ( .A1(n2212), .A2(n2288), .ZN(n2127) );
  INV_X1 U2726 ( .A(n2126), .ZN(n2128) );
  OAI22_X1 U2727 ( .A1(n2432), .A2(n1920), .B1(n2146), .B2(n2248), .ZN(n2126)
         );
  INV_X1 U2728 ( .A(n2291), .ZN(n2252) );
  NOR2_X1 U2729 ( .A1(n1543), .A2(n1662), .ZN(n2288) );
  NAND2_X1 U2730 ( .A1(n2174), .A2(n2124), .ZN(n2294) );
  NAND2_X1 U2731 ( .A1(\unit_decode/IMMreg/ffi_6/n4 ), .A2(n1567), .ZN(n2124)
         );
  NAND2_X1 U2732 ( .A1(n1342), .A2(\unit_decode/IMMreg/ffi_3/n4 ), .ZN(n2123)
         );
  AOI22_X1 U2733 ( .A1(n2554), .A2(n2407), .B1(n1577), .B2(n2406), .ZN(n2770)
         );
  NAND2_X1 U2734 ( .A1(n2091), .A2(n1745), .ZN(n2406) );
  NOR2_X1 U2735 ( .A1(n1692), .A2(n1746), .ZN(n1745) );
  NAND2_X1 U2736 ( .A1(n2120), .A2(n2092), .ZN(n1746) );
  NAND2_X1 U2737 ( .A1(n2090), .A2(n2571), .ZN(n2092) );
  INV_X1 U2738 ( .A(n1543), .ZN(n2571) );
  INV_X1 U2739 ( .A(n2390), .ZN(n2090) );
  NAND2_X1 U2740 ( .A1(n1450), .A2(n2775), .ZN(n2091) );
  INV_X1 U2741 ( .A(n2460), .ZN(n2407) );
  INV_X1 U2742 ( .A(n2528), .ZN(n2554) );
  NOR2_X1 U2743 ( .A1(n1927), .A2(n1542), .ZN(n2922) );
  INV_X1 U2744 ( .A(n1800), .ZN(n1799) );
  OAI21_X1 U2745 ( .B1(n2786), .B2(n1801), .A(n2141), .ZN(n1800) );
  INV_X1 U2746 ( .A(\unit_control/n153 ), .ZN(n2141) );
  NAND2_X1 U2747 ( .A1(n1802), .A2(n1842), .ZN(n1801) );
  NAND2_X1 U2748 ( .A1(n2816), .A2(n2782), .ZN(n1888) );
  NAND2_X1 U2749 ( .A1(n1808), .A2(n1807), .ZN(n1803) );
  AND2_X1 U2750 ( .A1(n2815), .A2(n2784), .ZN(n1807) );
  NAND2_X1 U2751 ( .A1(n1809), .A2(n1805), .ZN(n1804) );
  AND2_X1 U2752 ( .A1(n1806), .A2(n2746), .ZN(n1805) );
  NAND4_X1 U2753 ( .A1(n1810), .A2(n1806), .A3(n1654), .A4(n2784), .ZN(n1809)
         );
  INV_X1 U2754 ( .A(n1890), .ZN(n1889) );
  OAI21_X1 U2755 ( .B1(n2815), .B2(n2784), .A(n2739), .ZN(n1890) );
  NOR2_X1 U2756 ( .A1(n1892), .A2(\unit_fetch/pc_regout[5] ), .ZN(n1891) );
  NAND4_X1 U2757 ( .A1(n1895), .A2(n1894), .A3(n1893), .A4(n1677), .ZN(n1892)
         );
  NOR2_X1 U2758 ( .A1(n2720), .A2(n2861), .ZN(n1893) );
  NOR2_X1 U2759 ( .A1(n2718), .A2(n2719), .ZN(n1894) );
  NOR2_X1 U2760 ( .A1(n2716), .A2(n2717), .ZN(n1895) );
  NAND2_X1 U2761 ( .A1(n1900), .A2(n1901), .ZN(n1899) );
  NOR2_X1 U2762 ( .A1(n2653), .A2(n2651), .ZN(n1900) );
  INV_X1 U2763 ( .A(n2652), .ZN(n1901) );
  INV_X1 U2764 ( .A(n1867), .ZN(n2590) );
  OAI21_X1 U2765 ( .B1(n2588), .B2(n1870), .A(n1868), .ZN(n1867) );
  NOR2_X1 U2766 ( .A1(n2586), .A2(n1869), .ZN(n1868) );
  NAND2_X1 U2767 ( .A1(n1690), .A2(n1655), .ZN(n1869) );
  NOR3_X1 U2768 ( .A1(n1534), .A2(n2585), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2586) );
  NAND2_X1 U2769 ( .A1(n2585), .A2(n1871), .ZN(n1870) );
  NOR2_X1 U2770 ( .A1(n1534), .A2(n1660), .ZN(n1871) );
  INV_X1 U2771 ( .A(n2583), .ZN(n1872) );
  OAI21_X1 U2772 ( .B1(n2582), .B2(n1874), .A(n2584), .ZN(n1873) );
  NAND2_X1 U2773 ( .A1(n2218), .A2(n2220), .ZN(n1874) );
  AOI21_X1 U2774 ( .B1(n2622), .B2(n2621), .A(n2620), .ZN(n2654) );
  AOI211_X1 U2775 ( .C1(n2617), .C2(n2626), .A(n2616), .B(n2615), .ZN(n2618)
         );
  NOR2_X1 U2776 ( .A1(n2612), .A2(n2611), .ZN(n2613) );
  NAND2_X1 U2777 ( .A1(n2572), .A2(n1661), .ZN(n2778) );
  NOR2_X1 U2778 ( .A1(n1336), .A2(n1341), .ZN(n2572) );
  NAND2_X1 U2779 ( .A1(n2535), .A2(n2622), .ZN(n2608) );
  NOR2_X1 U2780 ( .A1(n1963), .A2(\unit_decode/IMMreg/ffi_2/n4 ), .ZN(n2535)
         );
  NAND2_X1 U2781 ( .A1(n1390), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .ZN(n1963)
         );
  INV_X1 U2782 ( .A(n1549), .ZN(n2164) );
  NOR2_X1 U2783 ( .A1(n2515), .A2(n2780), .ZN(n2602) );
  MUX2_X1 U2784 ( .A(n1962), .B(n1961), .S(n1940), .Z(n2515) );
  NOR2_X1 U2785 ( .A1(n2528), .A2(n2780), .ZN(n2604) );
  MUX2_X1 U2786 ( .A(n1965), .B(n1964), .S(n1937), .Z(n2528) );
  OAI211_X1 U2787 ( .C1(n2601), .C2(n2774), .A(n2600), .B(n2599), .ZN(n2621)
         );
  AOI22_X1 U2788 ( .A1(n2598), .A2(n2597), .B1(n2596), .B2(n2595), .ZN(n2599)
         );
  MUX2_X1 U2789 ( .A(n1950), .B(n1949), .S(n1937), .Z(n2596) );
  INV_X1 U2790 ( .A(n1961), .ZN(n1949) );
  NAND2_X1 U2791 ( .A1(n1954), .A2(\unit_decode/IMMreg/ffi_2/n4 ), .ZN(n1961)
         );
  INV_X1 U2792 ( .A(n1962), .ZN(n1950) );
  INV_X1 U2793 ( .A(n1964), .ZN(n1955) );
  NAND2_X1 U2794 ( .A1(n1954), .A2(n1665), .ZN(n1964) );
  NOR2_X1 U2795 ( .A1(n1612), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .ZN(n1954)
         );
  INV_X1 U2796 ( .A(n1965), .ZN(n1956) );
  NAND2_X1 U2797 ( .A1(n1653), .A2(n1576), .ZN(n1965) );
  AOI22_X1 U2798 ( .A1(n2594), .A2(n2593), .B1(n2592), .B2(n2612), .ZN(n2600)
         );
  NAND2_X1 U2799 ( .A1(n1944), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .ZN(n2777)
         );
  INV_X1 U2800 ( .A(n1966), .ZN(n1951) );
  NAND2_X1 U2801 ( .A1(n1664), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .ZN(n1966)
         );
  NAND3_X1 U2802 ( .A1(n1909), .A2(\unit_decode/IMMreg/ffi_0/n4 ), .A3(n1576), 
        .ZN(n2774) );
  INV_X1 U2803 ( .A(n1952), .ZN(n1953) );
  INV_X1 U2804 ( .A(n2751), .ZN(n1946) );
  INV_X1 U2805 ( .A(n1945), .ZN(n1738) );
  NOR2_X1 U2806 ( .A1(n1781), .A2(n1780), .ZN(n1850) );
  OR2_X1 U2807 ( .A1(n2651), .A2(n1706), .ZN(n1780) );
  XNOR2_X1 U2808 ( .A(n2223), .B(n2583), .ZN(n2651) );
  XNOR2_X1 U2809 ( .A(n2587), .B(n2585), .ZN(n2583) );
  AOI21_X1 U2810 ( .B1(n2221), .B2(n2220), .A(n2219), .ZN(n2222) );
  INV_X1 U2811 ( .A(n2241), .ZN(n2221) );
  AOI21_X1 U2812 ( .B1(n2239), .B2(n2220), .A(n2219), .ZN(n2584) );
  NOR2_X1 U2813 ( .A1(n2244), .A2(n1363), .ZN(n2219) );
  OR2_X1 U2814 ( .A1(n2653), .A2(n2652), .ZN(n1781) );
  XNOR2_X1 U2815 ( .A(n2242), .B(n2581), .ZN(n2653) );
  INV_X1 U2816 ( .A(n2239), .ZN(n2240) );
  OAI21_X1 U2817 ( .B1(n2580), .B2(n2263), .A(n2215), .ZN(n2239) );
  AOI21_X1 U2818 ( .B1(n2218), .B2(n2217), .A(n2216), .ZN(n2241) );
  INV_X1 U2819 ( .A(n2215), .ZN(n2216) );
  INV_X1 U2820 ( .A(n2260), .ZN(n2217) );
  XNOR2_X1 U2821 ( .A(n2264), .B(n2580), .ZN(n2652) );
  NAND2_X1 U2822 ( .A1(n2215), .A2(n2214), .ZN(n2580) );
  NAND2_X1 U2823 ( .A1(n2267), .A2(n2213), .ZN(n2214) );
  NAND2_X1 U2824 ( .A1(n2253), .A2(n2305), .ZN(n2215) );
  INV_X1 U2825 ( .A(n2267), .ZN(n2253) );
  NAND2_X1 U2826 ( .A1(n2582), .A2(n2263), .ZN(n2264) );
  INV_X1 U2827 ( .A(n2261), .ZN(n2263) );
  INV_X1 U2828 ( .A(n2275), .ZN(n2276) );
  NOR2_X1 U2829 ( .A1(n2261), .A2(n2260), .ZN(n2275) );
  AND2_X1 U2830 ( .A1(n2278), .A2(n2210), .ZN(n2260) );
  NOR2_X1 U2831 ( .A1(n2278), .A2(n2210), .ZN(n2261) );
  AND2_X1 U2832 ( .A1(n1834), .A2(n1860), .ZN(n1771) );
  AND2_X1 U2833 ( .A1(n1862), .A2(n2643), .ZN(n1835) );
  NAND2_X1 U2834 ( .A1(n1569), .A2(n1827), .ZN(n1826) );
  INV_X1 U2835 ( .A(n1557), .ZN(n1827) );
  NOR2_X1 U2836 ( .A1(n1712), .A2(n1721), .ZN(n1714) );
  NOR2_X1 U2837 ( .A1(n2644), .A2(n2645), .ZN(n1884) );
  AOI21_X1 U2838 ( .B1(n1885), .B2(n1375), .A(n2301), .ZN(n1856) );
  AND2_X1 U2839 ( .A1(n1656), .A2(n1905), .ZN(n1904) );
  AND2_X1 U2840 ( .A1(n1795), .A2(n2352), .ZN(n1905) );
  OR2_X1 U2841 ( .A1(n2301), .A2(n2300), .ZN(n1795) );
  NAND2_X1 U2842 ( .A1(n1712), .A2(n2423), .ZN(n1765) );
  NOR2_X1 U2843 ( .A1(n2480), .A2(n1719), .ZN(n1766) );
  NOR2_X1 U2844 ( .A1(n1816), .A2(n2640), .ZN(n1815) );
  NOR2_X1 U2845 ( .A1(n1536), .A2(n1721), .ZN(n1713) );
  AOI21_X1 U2846 ( .B1(n2444), .B2(n2443), .A(n1536), .ZN(n2447) );
  NAND2_X1 U2847 ( .A1(n1715), .A2(n1724), .ZN(n2444) );
  NOR4_X1 U2848 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n2639)
         );
  OAI21_X1 U2849 ( .B1(n1548), .B2(n1384), .A(n2526), .ZN(n2630) );
  INV_X1 U2850 ( .A(n1392), .ZN(n2526) );
  INV_X1 U2851 ( .A(n1622), .ZN(n2566) );
  INV_X1 U2852 ( .A(n2562), .ZN(n2563) );
  XNOR2_X1 U2853 ( .A(n2111), .B(n2187), .ZN(n2635) );
  XNOR2_X1 U2854 ( .A(n2503), .B(n2502), .ZN(n2638) );
  AOI21_X1 U2855 ( .B1(n2521), .B2(n1396), .A(n2501), .ZN(n2503) );
  AOI21_X1 U2856 ( .B1(n2524), .B2(n2500), .A(n2499), .ZN(n2521) );
  AOI21_X1 U2857 ( .B1(n2498), .B2(n1545), .A(n2496), .ZN(n2499) );
  INV_X1 U2858 ( .A(n2495), .ZN(n2496) );
  NAND2_X1 U2859 ( .A1(n1902), .A2(n2054), .ZN(n2524) );
  NOR2_X1 U2860 ( .A1(n2525), .A2(n2057), .ZN(n2058) );
  INV_X1 U2861 ( .A(n2069), .ZN(n2057) );
  XNOR2_X1 U2862 ( .A(n2023), .B(n2022), .ZN(n2624) );
  XNOR2_X1 U2863 ( .A(n1630), .B(n2053), .ZN(n2022) );
  NOR2_X1 U2864 ( .A1(n2014), .A2(n2013), .ZN(n2021) );
  INV_X1 U2865 ( .A(n2050), .ZN(n2013) );
  AOI21_X1 U2866 ( .B1(n2567), .B2(n2011), .A(n1352), .ZN(n2014) );
  NAND2_X1 U2867 ( .A1(n2009), .A2(n1555), .ZN(n2567) );
  INV_X1 U2868 ( .A(n2005), .ZN(n2006) );
  INV_X1 U2869 ( .A(n2109), .ZN(n2096) );
  INV_X1 U2870 ( .A(n2187), .ZN(n2097) );
  AND2_X1 U2871 ( .A1(n2110), .A2(n1854), .ZN(n1853) );
  NAND2_X1 U2872 ( .A1(n2502), .A2(n2188), .ZN(n1854) );
  INV_X1 U2873 ( .A(n2107), .ZN(n2108) );
  INV_X1 U2874 ( .A(n2186), .ZN(n2501) );
  OAI21_X1 U2875 ( .B1(n1720), .B2(n2424), .A(n1716), .ZN(n1722) );
  NOR2_X1 U2876 ( .A1(n1717), .A2(n2429), .ZN(n1716) );
  INV_X1 U2877 ( .A(n2446), .ZN(n2443) );
  NOR2_X1 U2878 ( .A1(n1723), .A2(n1718), .ZN(n1717) );
  NAND2_X1 U2879 ( .A1(n1724), .A2(n1719), .ZN(n1718) );
  OR2_X1 U2880 ( .A1(n1723), .A2(n1721), .ZN(n1720) );
  INV_X1 U2881 ( .A(n1635), .ZN(n1723) );
  INV_X1 U2882 ( .A(n2646), .ZN(n1814) );
  NOR2_X1 U2883 ( .A1(n1699), .A2(n2370), .ZN(n1783) );
  INV_X1 U2884 ( .A(n1907), .ZN(n1785) );
  AND2_X1 U2885 ( .A1(n2648), .A2(n2647), .ZN(n1898) );
  OR2_X1 U2886 ( .A1(n1865), .A2(n1858), .ZN(n1832) );
  INV_X1 U2887 ( .A(n1885), .ZN(n1858) );
  OR2_X1 U2888 ( .A1(n1906), .A2(n2370), .ZN(n1885) );
  INV_X1 U2889 ( .A(n2204), .ZN(n2205) );
  AND2_X1 U2890 ( .A1(n1643), .A2(n2202), .ZN(n1701) );
  NOR2_X1 U2891 ( .A1(n1864), .A2(n1696), .ZN(n1863) );
  AND2_X1 U2892 ( .A1(n1797), .A2(n2211), .ZN(n1696) );
  INV_X1 U2893 ( .A(n2210), .ZN(n2211) );
  NOR2_X1 U2894 ( .A1(n1866), .A2(n2319), .ZN(n1864) );
  NOR2_X1 U2895 ( .A1(n2374), .A2(n2203), .ZN(n2301) );
  INV_X1 U2896 ( .A(n2206), .ZN(n2203) );
  NAND2_X1 U2897 ( .A1(n1658), .A2(n1574), .ZN(n1865) );
  AND2_X1 U2898 ( .A1(n2207), .A2(n2353), .ZN(n2302) );
  XNOR2_X1 U2899 ( .A(\unit_decode/IMMreg/ffi_24/n4 ), .B(n1909), .ZN(n2207)
         );
  XNOR2_X1 U2900 ( .A(n2374), .B(n2206), .ZN(n2300) );
  XNOR2_X1 U2901 ( .A(n1941), .B(\unit_decode/IMMreg/ffi_23/n4 ), .ZN(n2206)
         );
  XNOR2_X1 U2902 ( .A(n2146), .B(n2077), .ZN(n2502) );
  NAND2_X1 U2903 ( .A1(n2162), .A2(n1512), .ZN(n2107) );
  NAND2_X1 U2904 ( .A1(n2186), .A2(n2188), .ZN(n2190) );
  NAND2_X1 U2905 ( .A1(n2510), .A2(n2078), .ZN(n2188) );
  INV_X1 U2906 ( .A(n2077), .ZN(n2078) );
  INV_X1 U2907 ( .A(n2146), .ZN(n2510) );
  NAND2_X1 U2908 ( .A1(n2522), .A2(n2076), .ZN(n2186) );
  INV_X1 U2909 ( .A(n2155), .ZN(n2522) );
  XNOR2_X1 U2910 ( .A(n2155), .B(n2076), .ZN(n2520) );
  AND2_X1 U2911 ( .A1(n2168), .A2(n2053), .ZN(n2071) );
  NAND2_X1 U2912 ( .A1(n2135), .A2(n2068), .ZN(n2495) );
  INV_X1 U2913 ( .A(n2067), .ZN(n2068) );
  INV_X1 U2914 ( .A(n2151), .ZN(n2135) );
  NAND2_X1 U2915 ( .A1(n2229), .A2(n2020), .ZN(n2048) );
  INV_X1 U2916 ( .A(n2172), .ZN(n2229) );
  NAND2_X1 U2917 ( .A1(n2158), .A2(n2047), .ZN(n2049) );
  INV_X1 U2918 ( .A(n2053), .ZN(n2047) );
  INV_X1 U2919 ( .A(n2168), .ZN(n2158) );
  INV_X1 U2920 ( .A(n1558), .ZN(n2251) );
  AND2_X1 U2921 ( .A1(n2143), .A2(n2125), .ZN(n2562) );
  OR2_X1 U2922 ( .A1(n2154), .A2(n1538), .ZN(n1991) );
  INV_X1 U2923 ( .A(n1967), .ZN(n1756) );
  NOR2_X1 U2924 ( .A1(n1554), .A2(n2192), .ZN(n2193) );
  XNOR2_X1 U2925 ( .A(\unit_decode/IMMreg/ffi_14/n4 ), .B(n1938), .ZN(n2192)
         );
  AND2_X1 U2926 ( .A1(n1834), .A2(n1656), .ZN(n1831) );
  AOI21_X1 U2927 ( .B1(n2445), .B2(n1632), .A(n2428), .ZN(n2430) );
  NOR2_X1 U2928 ( .A1(n2451), .A2(n2199), .ZN(n2428) );
  NAND2_X1 U2929 ( .A1(n2474), .A2(n2198), .ZN(n2425) );
  XNOR2_X1 U2930 ( .A(n1616), .B(\unit_decode/IMMreg/ffi_17/n4 ), .ZN(n2198)
         );
  NAND2_X1 U2931 ( .A1(n1934), .A2(\unit_decode/Areg/ffi_17/n4 ), .ZN(n1779)
         );
  NAND2_X1 U2932 ( .A1(n1385), .A2(\unit_decode/NPC1reg/ffi_17/n4 ), .ZN(n1778) );
  AND3_X1 U2933 ( .A1(n1796), .A2(n1382), .A3(n1569), .ZN(n1656) );
  INV_X1 U2934 ( .A(n2200), .ZN(n2201) );
  XNOR2_X1 U2935 ( .A(n1941), .B(\unit_decode/IMMreg/ffi_20/n4 ), .ZN(n2200)
         );
  INV_X1 U2936 ( .A(n2290), .ZN(n2417) );
  AND2_X1 U2937 ( .A1(n2369), .A2(n2431), .ZN(n1796) );
  XNOR2_X1 U2938 ( .A(n1941), .B(\unit_decode/IMMreg/ffi_19/n4 ), .ZN(n2202)
         );
  XNOR2_X1 U2939 ( .A(n1941), .B(\unit_decode/IMMreg/ffi_22/n4 ), .ZN(n2204)
         );
  INV_X1 U2940 ( .A(n2745), .ZN(n1806) );
  NAND2_X1 U2941 ( .A1(\unit_decode/IMMreg/ffi_3/n4 ), .A2(n1946), .ZN(n2289)
         );
  XNOR2_X1 U2942 ( .A(n1660), .B(n1938), .ZN(n2305) );
  INV_X1 U2943 ( .A(n2305), .ZN(n2213) );
  INV_X1 U2944 ( .A(n1379), .ZN(n2319) );
  XNOR2_X1 U2945 ( .A(n2244), .B(n1363), .ZN(n2581) );
  INV_X1 U2946 ( .A(n2581), .ZN(n2220) );
  INV_X1 U2947 ( .A(n2304), .ZN(n2333) );
  NAND2_X1 U2948 ( .A1(n2417), .A2(n2200), .ZN(n2389) );
  INV_X1 U2949 ( .A(n2488), .ZN(n1736) );
  INV_X1 U2950 ( .A(n2327), .ZN(n1797) );
  INV_X1 U2951 ( .A(n2608), .ZN(n1740) );
  INV_X1 U2952 ( .A(n2289), .ZN(n1917) );
  INV_X1 U2953 ( .A(n2486), .ZN(n1719) );
  INV_X1 U2954 ( .A(n1393), .ZN(n2054) );
  NAND2_X1 U2955 ( .A1(n2304), .A2(n1883), .ZN(n1676) );
  XNOR2_X1 U2956 ( .A(n2388), .B(n2204), .ZN(n2369) );
  INV_X1 U2957 ( .A(n2369), .ZN(n1907) );
  INV_X1 U2958 ( .A(n2580), .ZN(n2218) );
  AND3_X1 U2959 ( .A1(n1821), .A2(n1819), .A3(n1818), .ZN(n1686) );
  INV_X1 U2960 ( .A(n2307), .ZN(n2212) );
  OR2_X1 U2961 ( .A1(n2291), .A2(n1532), .ZN(n1688) );
  AND2_X1 U2962 ( .A1(n1673), .A2(n1341), .ZN(n1690) );
  AND2_X1 U2963 ( .A1(n1736), .A2(n2175), .ZN(n1691) );
  AND2_X1 U2964 ( .A1(n2098), .A2(n2175), .ZN(n1692) );
  INV_X1 U2965 ( .A(n2300), .ZN(n2371) );
  AND2_X1 U2966 ( .A1(n1926), .A2(\unit_fetch/pc_regout[0] ), .ZN(n1693) );
  OR2_X1 U2967 ( .A1(n2301), .A2(n2370), .ZN(n1694) );
  AOI21_X1 U2968 ( .B1(n2443), .B2(n1362), .A(n2428), .ZN(n2429) );
  NOR2_X1 U2969 ( .A1(n2353), .A2(n2207), .ZN(n2303) );
  AND2_X1 U2970 ( .A1(n1875), .A2(n2638), .ZN(n1695) );
  OR2_X1 U2971 ( .A1(n2291), .A2(n1590), .ZN(n1697) );
  INV_X1 U2972 ( .A(n2423), .ZN(n1724) );
  INV_X1 U2973 ( .A(n1724), .ZN(n1721) );
  AND2_X1 U2974 ( .A1(n1904), .A2(n1861), .ZN(n1698) );
  AND2_X1 U2975 ( .A1(n1785), .A2(n1551), .ZN(n1699) );
  NAND2_X1 U2976 ( .A1(n1388), .A2(n2197), .ZN(n2472) );
  INV_X1 U2977 ( .A(\unit_control/n152 ), .ZN(n1842) );
  NAND2_X1 U2978 ( .A1(n2290), .A2(n2201), .ZN(n2367) );
  NOR2_X1 U2979 ( .A1(n2388), .A2(n2205), .ZN(n2370) );
  INV_X1 U2980 ( .A(n2198), .ZN(n1777) );
  AND2_X1 U2981 ( .A1(n1784), .A2(n1785), .ZN(n1702) );
  AND2_X1 U2982 ( .A1(n1662), .A2(n1652), .ZN(n1703) );
  AND2_X1 U2983 ( .A1(n1765), .A2(n2472), .ZN(n1704) );
  OR2_X1 U2984 ( .A1(n1569), .A2(n1827), .ZN(n1705) );
  NAND2_X1 U2985 ( .A1(n1690), .A2(n1661), .ZN(n1706) );
  NAND2_X1 U2986 ( .A1(n1709), .A2(n1712), .ZN(n1708) );
  NOR2_X1 U2987 ( .A1(n1711), .A2(n1710), .ZN(n1709) );
  NAND2_X1 U2988 ( .A1(n1369), .A2(n1632), .ZN(n1710) );
  NOR2_X1 U2989 ( .A1(n2486), .A2(n2423), .ZN(n1711) );
  INV_X1 U2990 ( .A(n2480), .ZN(n1712) );
  NAND2_X1 U2991 ( .A1(n2424), .A2(n1600), .ZN(n1715) );
  NAND3_X1 U2992 ( .A1(n1575), .A2(n1703), .A3(n1738), .ZN(n2029) );
  XNOR2_X1 U2993 ( .A(n1739), .B(n2333), .ZN(n2645) );
  NAND3_X1 U2994 ( .A1(n2765), .A2(n2766), .A3(n1750), .ZN(n1749) );
  NOR3_X1 U2995 ( .A1(n2187), .A2(n2485), .A3(n1608), .ZN(n2189) );
  NAND2_X1 U2996 ( .A1(n2107), .A2(n2109), .ZN(n2187) );
  INV_X1 U2997 ( .A(n2162), .ZN(n2286) );
  NAND2_X1 U2998 ( .A1(n1913), .A2(\unit_decode/NPC1reg/ffi_0/n4 ), .ZN(n1755)
         );
  INV_X1 U2999 ( .A(\unit_control/uut_third_stage/ffi_19/n5 ), .ZN(n1757) );
  NAND2_X1 U3000 ( .A1(\unit_control/uut_third_stage/ffi_19/n5 ), .A2(
        \unit_decode/Areg/ffi_0/n4 ), .ZN(n1758) );
  OAI21_X1 U3001 ( .B1(n1920), .B2(n1759), .A(n1688), .ZN(n2134) );
  INV_X1 U3002 ( .A(n2474), .ZN(n1759) );
  AND2_X1 U3003 ( .A1(n1778), .A2(n1779), .ZN(n2474) );
  NAND2_X1 U3004 ( .A1(n2098), .A2(n2093), .ZN(n1760) );
  OAI21_X1 U3005 ( .B1(n2108), .B2(n1373), .A(n1760), .ZN(n2110) );
  OAI211_X1 U3006 ( .C1(n1705), .C2(n2414), .A(n1761), .B(n1826), .ZN(n2643)
         );
  NAND2_X1 U3007 ( .A1(n2414), .A2(n1569), .ZN(n1761) );
  AND2_X1 U3008 ( .A1(n1879), .A2(n1763), .ZN(n1762) );
  AND2_X1 U3009 ( .A1(n1382), .A2(n1877), .ZN(n1763) );
  NAND2_X1 U3010 ( .A1(n1656), .A2(n1375), .ZN(n1857) );
  NAND2_X1 U3011 ( .A1(n1764), .A2(n1704), .ZN(n1768) );
  XNOR2_X1 U3012 ( .A(n1768), .B(n1767), .ZN(n2642) );
  INV_X1 U3013 ( .A(n2427), .ZN(n1767) );
  AND2_X1 U3014 ( .A1(n2416), .A2(n2415), .ZN(n1769) );
  NAND3_X1 U3015 ( .A1(n1368), .A2(n1698), .A3(n1771), .ZN(n1770) );
  NAND2_X1 U3016 ( .A1(n2685), .A2(n1772), .ZN(
        \unit_fetch/unit_programCounter/ffi_0/n5 ) );
  OR2_X1 U3017 ( .A1(n2922), .A2(\unit_fetch/unit_programCounter/ffi_0/n4 ), 
        .ZN(n1772) );
  NAND2_X1 U3018 ( .A1(n1773), .A2(n1866), .ZN(n2318) );
  NAND2_X1 U3019 ( .A1(n1774), .A2(n1658), .ZN(n1773) );
  NAND2_X1 U3020 ( .A1(n1833), .A2(n1858), .ZN(n1774) );
  NAND2_X1 U3021 ( .A1(n1368), .A2(n1831), .ZN(n1833) );
  INV_X1 U3022 ( .A(n1778), .ZN(n1775) );
  INV_X1 U3023 ( .A(n2473), .ZN(n2427) );
  INV_X1 U3024 ( .A(n1779), .ZN(n1776) );
  NAND2_X1 U3025 ( .A1(n1782), .A2(n1783), .ZN(n2372) );
  NAND3_X1 U3026 ( .A1(n1609), .A2(n1702), .A3(n1879), .ZN(n1782) );
  NAND3_X1 U3027 ( .A1(n1609), .A2(n1377), .A3(n1877), .ZN(n2416) );
  NAND2_X1 U3028 ( .A1(n1788), .A2(n1786), .ZN(n2644) );
  NAND2_X1 U3029 ( .A1(n1855), .A2(n1787), .ZN(n1786) );
  INV_X1 U3030 ( .A(n1882), .ZN(n1787) );
  OAI21_X1 U3031 ( .B1(n1790), .B2(n1882), .A(n1789), .ZN(n1788) );
  XNOR2_X1 U3032 ( .A(n1856), .B(n2352), .ZN(n1789) );
  NAND2_X1 U3033 ( .A1(n1856), .A2(n1791), .ZN(n1790) );
  INV_X1 U3034 ( .A(n1857), .ZN(n1791) );
  NAND3_X1 U3035 ( .A1(n1886), .A2(n1621), .A3(n2748), .ZN(n2785) );
  NAND3_X1 U3036 ( .A1(n1886), .A2(n1621), .A3(n2786), .ZN(n2787) );
  INV_X1 U3037 ( .A(n2748), .ZN(n1802) );
  INV_X1 U3038 ( .A(n2786), .ZN(n2742) );
  NAND3_X1 U3039 ( .A1(n1811), .A2(n1810), .A3(n1683), .ZN(n1808) );
  NOR2_X1 U3040 ( .A1(n1829), .A2(n2423), .ZN(n1828) );
  INV_X1 U3041 ( .A(n2430), .ZN(n1829) );
  AND2_X1 U3042 ( .A1(n2189), .A2(n1854), .ZN(n1830) );
  INV_X1 U3043 ( .A(n2642), .ZN(n1836) );
  AOI21_X1 U3044 ( .B1(n2111), .B2(n2097), .A(n2096), .ZN(n1837) );
  INV_X1 U3045 ( .A(n1904), .ZN(n1838) );
  NAND2_X1 U3046 ( .A1(n2390), .A2(n1841), .ZN(n1839) );
  XNOR2_X1 U3047 ( .A(n1908), .B(\unit_decode/IMMreg/ffi_21/n4 ), .ZN(n1841)
         );
  OR2_X1 U3048 ( .A1(n1841), .A2(n2390), .ZN(n1840) );
  XNOR2_X1 U3049 ( .A(n1941), .B(n1679), .ZN(n2199) );
  NAND2_X1 U3050 ( .A1(n2685), .A2(n1846), .ZN(
        \unit_fetch/unit_npcregister/ffi_0/n5 ) );
  NOR2_X1 U3051 ( .A1(n1693), .A2(n1847), .ZN(n1846) );
  NOR2_X1 U3052 ( .A1(n1924), .A2(\unit_fetch/unit_npcregister/ffi_0/n4 ), 
        .ZN(n1847) );
  NAND2_X1 U3053 ( .A1(n2707), .A2(n1930), .ZN(n2685) );
  OAI21_X1 U3054 ( .B1(n2650), .B2(n1899), .A(n1897), .ZN(n1848) );
  NAND2_X1 U3055 ( .A1(n1850), .A2(n1625), .ZN(n1849) );
  NAND2_X1 U3056 ( .A1(n2194), .A2(n1372), .ZN(n1851) );
  INV_X1 U3057 ( .A(n1852), .ZN(n2637) );
  NOR2_X1 U3058 ( .A1(n1857), .A2(n2352), .ZN(n1855) );
  NAND2_X1 U3059 ( .A1(n2305), .A2(n2212), .ZN(n1859) );
  NAND2_X1 U3060 ( .A1(n2307), .A2(n2213), .ZN(n1860) );
  NOR2_X1 U3061 ( .A1(n2319), .A2(n2333), .ZN(n1861) );
  NOR2_X1 U3062 ( .A1(n2625), .A2(n1852), .ZN(n1862) );
  NAND2_X1 U3063 ( .A1(n1880), .A2(n1878), .ZN(n1877) );
  INV_X1 U3064 ( .A(n2431), .ZN(n1878) );
  INV_X1 U3065 ( .A(n1701), .ZN(n1880) );
  NAND3_X1 U3066 ( .A1(n2747), .A2(n1700), .A3(n1888), .ZN(n1887) );
  NAND2_X1 U3067 ( .A1(n2075), .A2(n2052), .ZN(n1902) );
  OAI21_X1 U3068 ( .B1(\unit_fetch/unit_npcregister/ffi_7/n4 ), .B2(n1922), 
        .A(n2680), .ZN(\unit_fetch/unit_npcregister/ffi_7/n5 ) );
  OAI21_X1 U3069 ( .B1(\unit_fetch/unit_npcregister/ffi_10/n4 ), .B2(n1921), 
        .A(n2677), .ZN(\unit_fetch/unit_npcregister/ffi_10/n5 ) );
  OR2_X1 U3070 ( .A1(n1617), .A2(n2171), .ZN(n2179) );
  NAND2_X1 U3071 ( .A1(n2687), .A2(n1931), .ZN(n2657) );
  AOI22_X1 U3072 ( .A1(n1931), .A2(n2918), .B1(n1927), .B2(
        \unit_fetch/adder_out[6] ), .ZN(n2681) );
  AOI22_X1 U3073 ( .A1(n1929), .A2(n2706), .B1(n1927), .B2(
        \unit_fetch/adder_out[4] ), .ZN(n2683) );
  AOI22_X1 U3074 ( .A1(n1930), .A2(n2916), .B1(n1926), .B2(
        \unit_fetch/adder_out[3] ), .ZN(n2684) );
  AOI22_X1 U3075 ( .A1(n1931), .A2(n2917), .B1(n1927), .B2(
        \unit_fetch/adder_out[5] ), .ZN(n2682) );
  AOI22_X1 U3076 ( .A1(n1931), .A2(n2692), .B1(n1926), .B2(
        \unit_fetch/adder_out[25] ), .ZN(n2662) );
  AOI22_X1 U3077 ( .A1(n2688), .A2(n1929), .B1(n1927), .B2(
        \unit_fetch/adder_out[29] ), .ZN(n2658) );
  AOI22_X1 U3078 ( .A1(n2689), .A2(n1929), .B1(n1927), .B2(
        \unit_fetch/adder_out[28] ), .ZN(n2659) );
  AOI22_X1 U3079 ( .A1(n2691), .A2(n1929), .B1(n1926), .B2(
        \unit_fetch/adder_out[26] ), .ZN(n2661) );
  INV_X1 U3080 ( .A(n1616), .ZN(n1908) );
  NAND2_X1 U3081 ( .A1(n2251), .A2(n2012), .ZN(n2050) );
  XNOR2_X1 U3082 ( .A(n2161), .B(n2012), .ZN(n2010) );
  INV_X1 U3083 ( .A(n1539), .ZN(n2052) );
  OAI21_X1 U3084 ( .B1(n2619), .B2(n1909), .A(n2618), .ZN(n2620) );
  NOR2_X1 U3085 ( .A1(n1633), .A2(n1909), .ZN(n2595) );
  NOR2_X1 U3086 ( .A1(n1630), .A2(n1937), .ZN(n2597) );
  NOR2_X1 U3087 ( .A1(n1617), .A2(n1909), .ZN(n2594) );
  XNOR2_X1 U3088 ( .A(n1937), .B(\unit_decode/IMMreg/ffi_31/n4 ), .ZN(n2585)
         );
  NOR2_X1 U3089 ( .A1(n1937), .A2(n2776), .ZN(n1944) );
  INV_X1 U3090 ( .A(n1636), .ZN(n2011) );
  NOR2_X1 U3091 ( .A1(n2566), .A2(n1636), .ZN(n2568) );
  NAND2_X1 U3092 ( .A1(\unit_decode/IMMreg/ffi_0/n4 ), .A2(n1623), .ZN(n1968)
         );
  NAND2_X1 U3093 ( .A1(n1652), .A2(n1561), .ZN(n2143) );
  XNOR2_X1 U3094 ( .A(\unit_decode/IMMreg/ffi_11/n4 ), .B(n1939), .ZN(n2077)
         );
  XNOR2_X1 U3095 ( .A(n1667), .B(n1939), .ZN(n2076) );
  XNOR2_X1 U3096 ( .A(n1561), .B(n1680), .ZN(n2012) );
  XNOR2_X1 U3097 ( .A(n1623), .B(\unit_decode/IMMreg/ffi_6/n4 ), .ZN(n2019) );
  NAND2_X1 U3098 ( .A1(n1646), .A2(n2055), .ZN(n2069) );
  INV_X1 U3099 ( .A(n2055), .ZN(n2056) );
  XNOR2_X1 U3100 ( .A(n2372), .B(n2371), .ZN(n2646) );
  OAI22_X1 U3101 ( .A1(n1626), .A2(n2030), .B1(n1633), .B2(n1918), .ZN(n1994)
         );
  OAI22_X1 U3102 ( .A1(n2390), .A2(n1918), .B1(n2249), .B2(n2248), .ZN(n2250)
         );
  NAND2_X1 U3103 ( .A1(n2249), .A2(n2094), .ZN(n2095) );
  INV_X1 U3104 ( .A(n2249), .ZN(n2098) );
  AOI22_X1 U3105 ( .A1(n2690), .A2(n1929), .B1(n1927), .B2(
        \unit_fetch/adder_out[27] ), .ZN(n2660) );
  NAND2_X1 U3106 ( .A1(n1991), .A2(n1980), .ZN(n2007) );
  XNOR2_X1 U3107 ( .A(n2588), .B(n1534), .ZN(n2591) );
  NAND2_X1 U3108 ( .A1(n2164), .A2(n1940), .ZN(n2609) );
  OAI21_X1 U3109 ( .B1(n1567), .B2(\unit_decode/IMMreg/ffi_6/n4 ), .A(n1940), 
        .ZN(n2030) );
  NAND2_X1 U3110 ( .A1(n1661), .A2(n1940), .ZN(n1945) );
  INV_X1 U3111 ( .A(n2093), .ZN(n2094) );
  XNOR2_X1 U3112 ( .A(n1672), .B(n1936), .ZN(n2093) );
  BUF_X1 U3113 ( .A(n2046), .Z(n1912) );
  AOI22_X1 U3114 ( .A1(n1970), .A2(n1940), .B1(n2628), .B2(n2617), .ZN(n1974)
         );
  NAND2_X1 U3115 ( .A1(n2572), .A2(n1940), .ZN(n2611) );
  OAI21_X1 U3116 ( .B1(\unit_fetch/unit_programCounter/ffi_10/n4 ), .B2(n1922), 
        .A(n2677), .ZN(\unit_fetch/unit_programCounter/ffi_10/n5 ) );
  AOI22_X1 U3117 ( .A1(n1931), .A2(n2704), .B1(n1926), .B2(
        \unit_fetch/adder_out[10] ), .ZN(n2677) );
  NAND2_X1 U3118 ( .A1(n2542), .A2(n2056), .ZN(n2497) );
  XNOR2_X1 U3119 ( .A(\unit_control/uut_third_stage/ffi_9/n5 ), .B(n1681), 
        .ZN(n2055) );
  NAND2_X1 U3120 ( .A1(n2069), .A2(n2497), .ZN(n2523) );
  INV_X1 U3121 ( .A(n1533), .ZN(n2500) );
  INV_X1 U3122 ( .A(n1615), .ZN(n2498) );
  NOR2_X1 U3123 ( .A1(n2070), .A2(n2493), .ZN(n2074) );
  OAI21_X1 U3124 ( .B1(n2021), .B2(n1627), .A(n2048), .ZN(n2023) );
  OAI211_X1 U3125 ( .C1(n2051), .C2(n2050), .A(n2049), .B(n2048), .ZN(n2070)
         );
  INV_X1 U3126 ( .A(n2019), .ZN(n2020) );
  AOI222_X1 U3127 ( .A1(n2607), .A2(n2606), .B1(n2605), .B2(n2604), .C1(n1619), 
        .C2(n2602), .ZN(n2619) );
  AOI22_X1 U3128 ( .A1(n2597), .A2(n2535), .B1(n2592), .B2(n1619), .ZN(n1982)
         );
  OAI22_X1 U3129 ( .A1(n2171), .A2(n1628), .B1(n2291), .B2(n2146), .ZN(n2149)
         );
  NAND2_X1 U3130 ( .A1(n1619), .A2(n2175), .ZN(n1985) );
  NAND2_X1 U3131 ( .A1(n2252), .A2(n1619), .ZN(n2129) );
  NAND2_X1 U3132 ( .A1(n2603), .A2(n1989), .ZN(n1990) );
  OAI22_X1 U3133 ( .A1(n2024), .A2(n2550), .B1(n1532), .B2(n2777), .ZN(n1958)
         );
  OAI22_X1 U3134 ( .A1(n1590), .A2(n2030), .B1(n1532), .B2(n1918), .ZN(n1947)
         );
  OAI22_X1 U3135 ( .A1(n2171), .A2(n1532), .B1(n2209), .B2(n1920), .ZN(n2153)
         );
  INV_X1 U3136 ( .A(n1532), .ZN(n2605) );
  NOR2_X1 U3137 ( .A1(n1624), .A2(n2779), .ZN(n2614) );
  OAI22_X1 U3138 ( .A1(n1589), .A2(n2030), .B1(n1624), .B2(n1918), .ZN(n1952)
         );
  OAI22_X1 U3139 ( .A1(n2171), .A2(n1624), .B1(n2767), .B2(n2248), .ZN(n2160)
         );
  INV_X1 U3140 ( .A(n2610), .ZN(n2612) );
  AND2_X1 U3141 ( .A1(n1613), .A2(n1987), .ZN(n1916) );
  INV_X1 U3142 ( .A(n1988), .ZN(n1989) );
  XNOR2_X1 U3143 ( .A(n1981), .B(n2007), .ZN(n2627) );
  OAI21_X1 U3144 ( .B1(n1916), .B2(n2007), .A(n2006), .ZN(n2009) );
  OAI21_X1 U3145 ( .B1(n2493), .B2(n2072), .A(n2520), .ZN(n2073) );
  NOR3_X1 U3146 ( .A1(n2523), .A2(n2071), .A3(n2494), .ZN(n2072) );
  OAI21_X1 U3147 ( .B1(n2241), .B2(n1552), .A(n2240), .ZN(n2242) );
  AOI21_X1 U3148 ( .B1(n1552), .B2(n2584), .A(n2222), .ZN(n2223) );
  MUX2_X1 U3149 ( .A(n1956), .B(n1955), .S(n1940), .Z(n2598) );
  OAI21_X1 U3150 ( .B1(n2750), .B2(n2612), .A(n1940), .ZN(n1979) );
  NAND2_X1 U3151 ( .A1(n1616), .A2(\unit_decode/IMMreg/ffi_6/n4 ), .ZN(n2125)
         );
  OAI22_X1 U3152 ( .A1(n2448), .A2(n1565), .B1(n1628), .B2(n2449), .ZN(n1970)
         );
  OAI22_X1 U3153 ( .A1(n2155), .A2(n2030), .B1(n1565), .B2(n1918), .ZN(n1977)
         );
  OAI22_X1 U3154 ( .A1(n2171), .A2(n1565), .B1(n2327), .B2(n1918), .ZN(n2157)
         );
  OAI22_X1 U3155 ( .A1(n2291), .A2(n1565), .B1(n1631), .B2(n1919), .ZN(n2130)
         );
  OAI22_X1 U3156 ( .A1(n2155), .A2(n1919), .B1(n2154), .B2(n2773), .ZN(n2081)
         );
  INV_X1 U3157 ( .A(n2154), .ZN(n2607) );
  OAI211_X1 U3158 ( .C1(n2591), .C2(\unit_decode/IMMreg/ffi_31/n4 ), .A(n2590), 
        .B(n2589), .ZN(n2655) );
  INV_X1 U3159 ( .A(n1568), .ZN(n1978) );
  AND2_X1 U3160 ( .A1(n2707), .A2(n1942), .ZN(n2940) );
  NAND2_X1 U3161 ( .A1(n2262), .A2(n2275), .ZN(n2582) );
  XNOR2_X1 U3162 ( .A(n1552), .B(n2276), .ZN(n2649) );
  AOI21_X1 U3163 ( .B1(n2074), .B2(n2075), .A(n2073), .ZN(n2191) );
  OAI211_X1 U3164 ( .C1(n1610), .C2(n2544), .A(n2299), .B(n2298), .ZN(n2689)
         );
  XNOR2_X1 U3165 ( .A(\unit_decode/IMMreg/ffi_25/n4 ), .B(n1908), .ZN(n2208)
         );
  XNOR2_X1 U3166 ( .A(\unit_decode/IMMreg/ffi_3/n4 ), .B(
        \unit_control/uut_third_stage/ffi_9/n5 ), .ZN(n1988) );
  XNOR2_X1 U3167 ( .A(\unit_control/uut_third_stage/ffi_9/n5 ), .B(n1612), 
        .ZN(n1967) );
  INV_X1 U3168 ( .A(n1917), .ZN(n1919) );
  INV_X1 U3169 ( .A(n1917), .ZN(n1920) );
  INV_X1 U3170 ( .A(n1941), .ZN(n1939) );
  MUX2_X1 U3171 ( .A(\unit_decode/NPC1reg/ffi_1/n4 ), .B(
        \unit_decode/Areg/ffi_1/n4 ), .S(
        \unit_control/uut_third_stage/ffi_19/n5 ), .Z(n2150) );
  NAND3_X1 U3172 ( .A1(n1665), .A2(n1653), .A3(n1612), .ZN(n1962) );
  MUX2_X1 U3173 ( .A(\unit_decode/NPC1reg/ffi_7/n4 ), .B(
        \unit_decode/Areg/ffi_7/n4 ), .S(n1910), .Z(n2168) );
  MUX2_X1 U3174 ( .A(\unit_decode/NPC1reg/ffi_4/n4 ), .B(
        \unit_decode/Areg/ffi_4/n4 ), .S(n1911), .Z(n2574) );
  MUX2_X1 U3175 ( .A(\unit_decode/NPC1reg/ffi_3/n4 ), .B(
        \unit_decode/Areg/ffi_3/n4 ), .S(n1914), .Z(n2147) );
  MUX2_X1 U3176 ( .A(n2778), .B(n2611), .S(n1390), .Z(n1972) );
  MUX2_X1 U3177 ( .A(n1972), .B(n1971), .S(n2605), .Z(n1973) );
  MUX2_X1 U3178 ( .A(\unit_decode/NPC1reg/ffi_10/n4 ), .B(
        \unit_decode/Areg/ffi_10/n4 ), .S(n1910), .Z(n2155) );
  MUX2_X1 U3179 ( .A(\unit_decode/NPC1reg/ffi_11/n4 ), .B(
        \unit_decode/Areg/ffi_11/n4 ), .S(n1910), .Z(n2146) );
  MUX2_X1 U3180 ( .A(\unit_decode/NPC1reg/ffi_12/n4 ), .B(
        \unit_decode/Areg/ffi_12/n4 ), .S(n1910), .Z(n2162) );
  MUX2_X1 U3181 ( .A(\unit_decode/NPC1reg/ffi_13/n4 ), .B(
        \unit_decode/Areg/ffi_13/n4 ), .S(n1911), .Z(n2249) );
  XOR2_X1 U3182 ( .A(n1627), .B(n2021), .Z(n2636) );
  MUX2_X1 U3183 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_6/n4 ), .Z(
        n2015) );
  MUX2_X1 U3184 ( .A(n2015), .B(n2576), .S(n1618), .Z(n2016) );
  MUX2_X1 U3185 ( .A(\unit_decode/NPC1reg/ffi_15/n4 ), .B(
        \unit_decode/Areg/ffi_15/n4 ), .S(n1910), .Z(n2488) );
  NAND3_X1 U3186 ( .A1(n2033), .A2(n2032), .A3(n2031), .ZN(n2037) );
  MUX2_X1 U3187 ( .A(n2573), .B(n2541), .S(\unit_decode/IMMreg/ffi_7/n4 ), .Z(
        n2034) );
  MUX2_X1 U3188 ( .A(n2035), .B(n2034), .S(n1630), .Z(n2036) );
  MUX2_X1 U3189 ( .A(\unit_decode/NPC1reg/ffi_16/n4 ), .B(
        \unit_decode/Areg/ffi_16/n4 ), .S(n1934), .Z(n2767) );
  MUX2_X1 U3190 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_9/n4 ), .Z(
        n2060) );
  MUX2_X1 U3191 ( .A(n2060), .B(n2059), .S(n2135), .Z(n2061) );
  MUX2_X1 U3192 ( .A(\unit_decode/NPC1reg/ffi_18/n4 ), .B(
        \unit_decode/Areg/ffi_18/n4 ), .S(n1934), .Z(n2451) );
  MUX2_X1 U3193 ( .A(\unit_decode/NPC1reg/ffi_20/n4 ), .B(
        \unit_decode/Areg/ffi_20/n4 ), .S(n1910), .Z(n2290) );
  MUX2_X1 U3194 ( .A(n2611), .B(n2778), .S(n1663), .Z(n2086) );
  MUX2_X1 U3195 ( .A(n2086), .B(n2085), .S(n2286), .Z(n2087) );
  MUX2_X1 U3196 ( .A(\unit_decode/NPC1reg/ffi_21/n4 ), .B(
        \unit_decode/Areg/ffi_21/n4 ), .S(n1910), .Z(n2390) );
  MUX2_X1 U3197 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_13/n4 ), 
        .Z(n2100) );
  MUX2_X1 U3198 ( .A(n2100), .B(n2099), .S(n2098), .Z(n2101) );
  MUX2_X1 U3199 ( .A(\unit_decode/NPC1reg/ffi_22/n4 ), .B(
        \unit_decode/Areg/ffi_22/n4 ), .S(n1934), .Z(n2388) );
  MUX2_X1 U3200 ( .A(n2573), .B(n2541), .S(\unit_decode/IMMreg/ffi_14/n4 ), 
        .Z(n2112) );
  MUX2_X1 U3201 ( .A(n2113), .B(n2112), .S(n1554), .Z(n2115) );
  MUX2_X1 U3202 ( .A(\unit_decode/NPC1reg/ffi_23/n4 ), .B(
        \unit_decode/Areg/ffi_23/n4 ), .S(n1910), .Z(n2374) );
  MUX2_X1 U3203 ( .A(\unit_decode/NPC1reg/ffi_24/n4 ), .B(
        \unit_decode/Areg/ffi_24/n4 ), .S(n1910), .Z(n2353) );
  MUX2_X1 U3204 ( .A(\unit_decode/NPC1reg/ffi_27/n4 ), .B(
        \unit_decode/Areg/ffi_27/n4 ), .S(n1935), .Z(n2307) );
  MUX2_X1 U3205 ( .A(\unit_decode/NPC1reg/ffi_26/n4 ), .B(
        \unit_decode/Areg/ffi_26/n4 ), .S(n1560), .Z(n2327) );
  MUX2_X1 U3206 ( .A(\unit_decode/NPC1reg/ffi_25/n4 ), .B(
        \unit_decode/Areg/ffi_25/n4 ), .S(n1910), .Z(n2209) );
  MUX2_X1 U3207 ( .A(\unit_decode/NPC1reg/ffi_29/n4 ), .B(
        \unit_decode/Areg/ffi_29/n4 ), .S(n1935), .Z(n2267) );
  MUX2_X1 U3208 ( .A(\unit_decode/NPC1reg/ffi_28/n4 ), .B(
        \unit_decode/Areg/ffi_28/n4 ), .S(n1935), .Z(n2278) );
  MUX2_X1 U3209 ( .A(\unit_decode/NPC1reg/ffi_30/n4 ), .B(
        \unit_decode/Areg/ffi_30/n4 ), .S(n1560), .Z(n2244) );
  MUX2_X1 U3210 ( .A(n2541), .B(n2573), .S(n1660), .Z(n2308) );
  MUX2_X1 U3211 ( .A(n2573), .B(n2541), .S(\unit_decode/IMMreg/ffi_31/n4 ), 
        .Z(n2326) );
  MUX2_X1 U3212 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_25/n4 ), 
        .Z(n2340) );
  NAND3_X1 U3213 ( .A1(n2339), .A2(n2570), .A3(n1689), .ZN(n2338) );
  MUX2_X1 U3214 ( .A(n2541), .B(n2573), .S(n1674), .Z(n2375) );
  MUX2_X1 U3215 ( .A(n2573), .B(n2541), .S(\unit_decode/IMMreg/ffi_22/n4 ), 
        .Z(n2387) );
  MUX2_X1 U3216 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_21/n4 ), 
        .Z(n2391) );
  MUX2_X1 U3217 ( .A(n2392), .B(n2391), .S(n1629), .Z(n2403) );
  MUX2_X1 U3218 ( .A(n2778), .B(n2611), .S(\unit_decode/IMMreg/ffi_20/n4 ), 
        .Z(n2419) );
  MUX2_X1 U3219 ( .A(n2419), .B(n2418), .S(n1346), .Z(n2420) );
  MUX2_X1 U3220 ( .A(n2541), .B(n2573), .S(n1675), .Z(n2433) );
  MUX2_X1 U3221 ( .A(n2434), .B(n2433), .S(n2432), .Z(n2435) );
  MUX2_X1 U3222 ( .A(n2541), .B(n2573), .S(n1679), .Z(n2452) );
  MUX2_X1 U3223 ( .A(n2453), .B(n2452), .S(n1631), .Z(n2454) );
  MUX2_X1 U3224 ( .A(n2611), .B(n2778), .S(n1666), .Z(n2476) );
  MUX2_X1 U3225 ( .A(n2476), .B(n2475), .S(n2474), .Z(n2477) );
  MUX2_X1 U3226 ( .A(n2541), .B(n2573), .S(n1669), .Z(n2489) );
  MUX2_X1 U3227 ( .A(n2490), .B(n2489), .S(n1378), .Z(n2491) );
  MUX2_X1 U3228 ( .A(n2541), .B(n2573), .S(n1681), .Z(n2543) );
  XOR2_X1 U3229 ( .A(n1549), .B(n2563), .Z(n2569) );
  MUX2_X1 U3230 ( .A(n2569), .B(n2568), .S(n2567), .Z(n2629) );
  MUX2_X1 U3231 ( .A(n2576), .B(n2575), .S(n1549), .Z(n2577) );
  NAND3_X1 U3232 ( .A1(n2588), .A2(n1534), .A3(\unit_decode/IMMreg/ffi_31/n4 ), 
        .ZN(n2589) );
  MUX2_X1 U3233 ( .A(n2614), .B(n2613), .S(\unit_decode/IMMreg/ffi_0/n4 ), .Z(
        n2615) );
  NAND2_X1 U3235 ( .A1(n1337), .A2(n1942), .ZN(n2932) );
  OAI21_X1 U3236 ( .B1(n2736), .B2(\unit_fetch/unit_instructionRegister/n50 ), 
        .A(n2735), .ZN(n2714) );
  INV_X1 U3237 ( .A(n2714), .ZN(n2715) );
  OAI21_X1 U3238 ( .B1(\unit_fetch/unit_instructionRegister/n57 ), .B2(n2737), 
        .A(n2715), .ZN(n2724) );
  INV_X1 U3239 ( .A(n2876), .ZN(n2822) );
  NAND4_X1 U3240 ( .A1(\unit_fetch/unit_programCounter/ffi_27/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_16/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_23/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_24/n4 ), .ZN(n2720) );
  NAND4_X1 U3241 ( .A1(\unit_fetch/unit_programCounter/ffi_25/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_17/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_15/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_19/n4 ), .ZN(n2719) );
  NAND4_X1 U3242 ( .A1(\unit_fetch/unit_programCounter/ffi_7/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_22/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_30/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_26/n4 ), .ZN(n2718) );
  NAND4_X1 U3243 ( .A1(\unit_fetch/unit_programCounter/ffi_8/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_9/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_21/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_29/n4 ), .ZN(n2717) );
  NAND4_X1 U3244 ( .A1(\unit_fetch/unit_programCounter/ffi_12/n4 ), .A2(
        \unit_fetch/unit_adder/add_19/n47 ), .A3(
        \unit_fetch/unit_programCounter/ffi_6/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_14/n4 ), .ZN(n2716) );
  NAND3_X1 U3245 ( .A1(n2878), .A2(n2908), .A3(n1603), .ZN(n2817) );
  NAND2_X1 U3246 ( .A1(\unit_fetch/unit_programCounter/ffi_5/n4 ), .A2(n1896), 
        .ZN(n2839) );
  NOR2_X1 U3247 ( .A1(\unit_fetch/unit_programCounter/ffi_3/n4 ), .A2(n2839), 
        .ZN(n2882) );
  NOR3_X1 U3248 ( .A1(\unit_fetch/unit_programCounter/ffi_5/n4 ), .A2(n1896), 
        .A3(\unit_fetch/pc_regout[3] ), .ZN(n2721) );
  OAI21_X1 U3249 ( .B1(n2882), .B2(n2721), .A(n2878), .ZN(n2880) );
  NAND2_X1 U3250 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(n2908), 
        .ZN(n2847) );
  OAI22_X1 U3251 ( .A1(n2817), .A2(n2839), .B1(n2880), .B2(n2847), .ZN(n2722)
         );
  INV_X1 U3252 ( .A(n2722), .ZN(n2828) );
  INV_X1 U3253 ( .A(n2724), .ZN(n2784) );
  OAI221_X1 U3254 ( .B1(\unit_fetch/unit_programCounter/ffi_4/n4 ), .B2(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .C1(
        \unit_fetch/unit_programCounter/ffi_4/n4 ), .C2(
        \unit_fetch/unit_programCounter/ffi_3/n4 ), .A(
        \unit_fetch/unit_programCounter/ffi_5/n4 ), .ZN(n2725) );
  NAND2_X1 U3255 ( .A1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .ZN(n2829) );
  OAI21_X1 U3256 ( .B1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .B2(n2725), 
        .A(n2728), .ZN(n2815) );
  OAI221_X1 U3257 ( .B1(n2737), .B2(\unit_fetch/unit_instructionRegister/n54 ), 
        .C1(n2736), .C2(\unit_fetch/unit_instructionRegister/n49 ), .A(n2735), 
        .ZN(n2781) );
  NOR2_X1 U3258 ( .A1(RST), .A2(n2781), .ZN(n2739) );
  NAND2_X1 U3259 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .ZN(n2833) );
  INV_X1 U3260 ( .A(n2725), .ZN(n2726) );
  AOI22_X1 U3261 ( .A1(n2791), .A2(n2833), .B1(n2726), .B2(
        \unit_fetch/pc_regout[1] ), .ZN(n2814) );
  NAND3_X1 U3262 ( .A1(\unit_fetch/pc_regout[0] ), .A2(n2732), .A3(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .ZN(n2727) );
  INV_X1 U3263 ( .A(n2869), .ZN(n2731) );
  NOR2_X1 U3264 ( .A1(\unit_fetch/unit_programCounter/ffi_4/n4 ), .A2(n2731), 
        .ZN(n2789) );
  NAND2_X1 U3265 ( .A1(n2869), .A2(n1603), .ZN(n2824) );
  NAND2_X1 U3266 ( .A1(\unit_fetch/unit_programCounter/ffi_4/n4 ), .A2(
        \unit_fetch/pc_regout[3] ), .ZN(n2733) );
  NAND3_X1 U3267 ( .A1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .ZN(n2887) );
  NAND3_X1 U3268 ( .A1(n2732), .A2(n2731), .A3(n2887), .ZN(n2813) );
  OAI221_X1 U3269 ( .B1(n2737), .B2(\unit_fetch/unit_instructionRegister/n56 ), 
        .C1(n2736), .C2(\unit_fetch/unit_instructionRegister/n51 ), .A(n2735), 
        .ZN(n2783) );
  OAI211_X1 U3270 ( .C1(\unit_decode/RD1reg/ffi_1/n4 ), .C2(n2741), .A(
        \unit_decode/RD1reg/ffi_0/n4 ), .B(\unit_decode/RD1reg/ffi_2/n4 ), 
        .ZN(n2744) );
  INV_X1 U3271 ( .A(n2814), .ZN(n2746) );
  OAI22_X1 U3272 ( .A1(\unit_decode/RD1reg/ffi_4/n4 ), .A2(n2746), .B1(
        \unit_decode/RD1reg/ffi_3/n4 ), .B2(n2815), .ZN(n2743) );
  OAI21_X1 U3273 ( .B1(n2744), .B2(n2743), .A(n2742), .ZN(n2747) );
  NAND3_X1 U3274 ( .A1(\unit_decode/RD1reg/ffi_4/n4 ), .A2(
        \unit_decode/RD1reg/ffi_1/n4 ), .A3(\unit_decode/RD1reg/ffi_3/n4 ), 
        .ZN(n2748) );
  NOR2_X1 U3275 ( .A1(RST), .A2(\unit_decode/RD1reg/ffi_0/n4 ), .ZN(n2935) );
  NOR2_X1 U3276 ( .A1(RST), .A2(\unit_decode/RD1reg/ffi_1/n4 ), .ZN(n2936) );
  NOR2_X1 U3277 ( .A1(RST), .A2(\unit_decode/RD1reg/ffi_2/n4 ), .ZN(n2937) );
  NOR2_X1 U3278 ( .A1(RST), .A2(\unit_decode/RD1reg/ffi_3/n4 ), .ZN(n2938) );
  NOR2_X1 U3279 ( .A1(RST), .A2(\unit_decode/RD1reg/ffi_4/n4 ), .ZN(n2939) );
  NAND2_X1 U3280 ( .A1(n1938), .A2(n1653), .ZN(n2749) );
  OAI21_X1 U3281 ( .B1(n1936), .B2(n1653), .A(n2749), .ZN(n2750) );
  NAND2_X1 U3282 ( .A1(n1612), .A2(\unit_decode/IMMreg/ffi_2/n4 ), .ZN(n2776)
         );
  NAND3_X1 U3283 ( .A1(n1936), .A2(\unit_decode/IMMreg/ffi_6/n4 ), .A3(n1342), 
        .ZN(n2751) );
  AND2_X1 U3284 ( .A1(n1943), .A2(n2910), .ZN(n2941) );
  AND2_X1 U3285 ( .A1(n1943), .A2(n2915), .ZN(n2942) );
  AND2_X1 U3286 ( .A1(n1943), .A2(n2916), .ZN(n2943) );
  AND2_X1 U3287 ( .A1(n1943), .A2(n2917), .ZN(n2945) );
  AND2_X1 U3288 ( .A1(n1943), .A2(n2918), .ZN(n2946) );
  AND2_X1 U3289 ( .A1(n1943), .A2(n2919), .ZN(n2947) );
  NOR2_X1 U3290 ( .A1(\unit_decode/IMMreg/ffi_3/n4 ), .A2(n2751), .ZN(n2775)
         );
  INV_X1 U3291 ( .A(n2775), .ZN(n2773) );
  AND2_X1 U3292 ( .A1(n1943), .A2(n2920), .ZN(n2949) );
  NOR3_X1 U3293 ( .A1(n2754), .A2(n2753), .A3(n2752), .ZN(n2755) );
  AND2_X1 U3294 ( .A1(n1943), .A2(n2912), .ZN(n2952) );
  AND2_X1 U3295 ( .A1(n1943), .A2(n2913), .ZN(n2953) );
  AND2_X1 U3296 ( .A1(n1943), .A2(n2914), .ZN(n2954) );
  NAND3_X1 U3297 ( .A1(n2763), .A2(n2762), .A3(n2761), .ZN(n2764) );
  NOR2_X1 U3298 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_0/n4 ), .ZN(n2972) );
  NOR2_X1 U3299 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_1/n4 ), .ZN(n2973) );
  NOR2_X1 U3300 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_2/n4 ), .ZN(n2974) );
  NOR2_X1 U3301 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_3/n4 ), .ZN(n2975) );
  NOR2_X1 U3302 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_4/n4 ), .ZN(n2976) );
  NOR2_X1 U3303 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_5/n4 ), .ZN(n2977) );
  NOR2_X1 U3304 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_6/n4 ), .ZN(n2978) );
  NOR2_X1 U3305 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_7/n4 ), .ZN(n2979) );
  NOR2_X1 U3306 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_8/n4 ), .ZN(n2980) );
  NOR2_X1 U3307 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_9/n4 ), .ZN(n2981) );
  NOR2_X1 U3308 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_10/n4 ), .ZN(n2982)
         );
  NOR2_X1 U3309 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_11/n4 ), .ZN(n2983)
         );
  NOR2_X1 U3310 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_12/n4 ), .ZN(n2984)
         );
  NOR2_X1 U3311 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_13/n4 ), .ZN(n2985)
         );
  NOR2_X1 U3312 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_14/n4 ), .ZN(n2986)
         );
  NOR2_X1 U3313 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_15/n4 ), .ZN(n2987)
         );
  NOR2_X1 U3314 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_16/n4 ), .ZN(n2988)
         );
  NOR2_X1 U3315 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_17/n4 ), .ZN(n2989)
         );
  NOR2_X1 U3316 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_18/n4 ), .ZN(n2990)
         );
  NOR2_X1 U3317 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_19/n4 ), .ZN(n2991)
         );
  NOR2_X1 U3318 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_20/n4 ), .ZN(n2992)
         );
  NOR2_X1 U3319 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_21/n4 ), .ZN(n2993)
         );
  NOR2_X1 U3320 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_22/n4 ), .ZN(n2994)
         );
  NOR2_X1 U3321 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_23/n4 ), .ZN(n2995)
         );
  NOR2_X1 U3322 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_24/n4 ), .ZN(n2996)
         );
  NOR2_X1 U3323 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_25/n4 ), .ZN(n2997)
         );
  NOR2_X1 U3324 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_26/n4 ), .ZN(n2998)
         );
  NOR2_X1 U3325 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_27/n4 ), .ZN(n2999)
         );
  NOR2_X1 U3326 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_28/n4 ), .ZN(n3000)
         );
  NOR2_X1 U3327 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_29/n4 ), .ZN(n3001)
         );
  NOR2_X1 U3328 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_30/n4 ), .ZN(n3002)
         );
  NOR2_X1 U3329 ( .A1(RST), .A2(\unit_decode/NPC1reg/ffi_31/n4 ), .ZN(n3003)
         );
  AND2_X1 U3330 ( .A1(n1943), .A2(n2781), .ZN(n3005) );
  AND2_X1 U3331 ( .A1(n1943), .A2(n2782), .ZN(n3006) );
  AND2_X1 U3332 ( .A1(n1943), .A2(n2783), .ZN(n3007) );
  NOR2_X1 U3333 ( .A1(RST), .A2(n2784), .ZN(n3008) );
  NOR2_X1 U3334 ( .A1(RST), .A2(n1806), .ZN(n3009) );
  NOR2_X1 U3335 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n38 ), 
        .ZN(n3010) );
  NOR2_X1 U3336 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n40 ), 
        .ZN(n3011) );
  NOR2_X1 U3337 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n41 ), 
        .ZN(n3012) );
  NOR2_X1 U3338 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n42 ), 
        .ZN(n3013) );
  NOR2_X1 U3339 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n43 ), 
        .ZN(n3014) );
  NOR2_X1 U3340 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n45 ), 
        .ZN(n3015) );
  NOR2_X1 U3341 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n46 ), 
        .ZN(n3016) );
  NOR2_X1 U3342 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n47 ), 
        .ZN(n3017) );
  NOR2_X1 U3343 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n48 ), 
        .ZN(n3018) );
  NOR2_X1 U3344 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n49 ), 
        .ZN(n3019) );
  NOR2_X1 U3345 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n50 ), 
        .ZN(n3020) );
  NOR2_X1 U3346 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n51 ), 
        .ZN(n3021) );
  NOR2_X1 U3347 ( .A1(RST), .A2(\unit_fetch/unit_instructionRegister/n53 ), 
        .ZN(n3022) );
  AND2_X1 U3348 ( .A1(\unit_decode/registerA[0] ), .A2(n1942), .ZN(n3023) );
  AND2_X1 U3349 ( .A1(\unit_decode/registerA[1] ), .A2(n1942), .ZN(n3024) );
  AND2_X1 U3350 ( .A1(\unit_decode/registerA[2] ), .A2(n1942), .ZN(n3025) );
  AND2_X1 U3351 ( .A1(\unit_decode/registerA[3] ), .A2(n1942), .ZN(n3026) );
  AND2_X1 U3352 ( .A1(\unit_decode/registerA[4] ), .A2(n1942), .ZN(n3027) );
  AND2_X1 U3353 ( .A1(\unit_decode/registerA[5] ), .A2(n1942), .ZN(n3028) );
  AND2_X1 U3354 ( .A1(\unit_decode/registerA[6] ), .A2(n1942), .ZN(n3029) );
  AND2_X1 U3355 ( .A1(\unit_decode/registerA[7] ), .A2(n1942), .ZN(n3030) );
  AND2_X1 U3356 ( .A1(\unit_decode/registerA[8] ), .A2(n1942), .ZN(n3031) );
  AND2_X1 U3357 ( .A1(\unit_decode/registerA[9] ), .A2(n1942), .ZN(n3032) );
  AND2_X1 U3358 ( .A1(\unit_decode/registerA[10] ), .A2(n1942), .ZN(n3033) );
  AND2_X1 U3359 ( .A1(\unit_decode/registerA[11] ), .A2(n1942), .ZN(n3034) );
  AND2_X1 U3360 ( .A1(\unit_decode/registerA[12] ), .A2(n1942), .ZN(n3035) );
  AND2_X1 U3361 ( .A1(\unit_decode/registerA[13] ), .A2(n1942), .ZN(n3036) );
  AND2_X1 U3362 ( .A1(\unit_decode/registerA[14] ), .A2(n1942), .ZN(n3037) );
  AND2_X1 U3363 ( .A1(\unit_decode/registerA[15] ), .A2(n1942), .ZN(n3038) );
  AND2_X1 U3364 ( .A1(\unit_decode/registerA[16] ), .A2(n1942), .ZN(n3039) );
  AND2_X1 U3365 ( .A1(\unit_decode/registerA[17] ), .A2(n1942), .ZN(n3040) );
  AND2_X1 U3366 ( .A1(\unit_decode/registerA[18] ), .A2(n1942), .ZN(n3041) );
  AND2_X1 U3367 ( .A1(\unit_decode/registerA[19] ), .A2(n1943), .ZN(n3042) );
  AND2_X1 U3368 ( .A1(\unit_decode/registerA[20] ), .A2(n1942), .ZN(n3043) );
  AND2_X1 U3369 ( .A1(\unit_decode/registerA[21] ), .A2(n1942), .ZN(n3044) );
  AND2_X1 U3370 ( .A1(\unit_decode/registerA[22] ), .A2(n1942), .ZN(n3045) );
  AND2_X1 U3371 ( .A1(\unit_decode/registerA[23] ), .A2(n1942), .ZN(n3046) );
  AND2_X1 U3372 ( .A1(\unit_decode/registerA[24] ), .A2(n1942), .ZN(n3047) );
  AND2_X1 U3373 ( .A1(\unit_decode/registerA[25] ), .A2(n1942), .ZN(n3048) );
  AND2_X1 U3374 ( .A1(\unit_decode/registerA[26] ), .A2(n1943), .ZN(n3049) );
  AND2_X1 U3375 ( .A1(\unit_decode/registerA[27] ), .A2(n1943), .ZN(n3050) );
  AND2_X1 U3376 ( .A1(\unit_decode/registerA[28] ), .A2(n1943), .ZN(n3051) );
  AND2_X1 U3377 ( .A1(\unit_decode/registerA[29] ), .A2(n1943), .ZN(n3052) );
  AND2_X1 U3378 ( .A1(\unit_decode/registerA[30] ), .A2(n1943), .ZN(n3053) );
  AND2_X1 U3379 ( .A1(\unit_decode/registerA[31] ), .A2(n1943), .ZN(n3054) );
  NOR2_X1 U3380 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_0/n4 ), .ZN(
        n3055) );
  NOR2_X1 U3381 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_1/n4 ), .ZN(
        n3056) );
  NOR2_X1 U3382 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_2/n4 ), .ZN(
        n3057) );
  NOR2_X1 U3383 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_3/n4 ), .ZN(
        n3058) );
  NOR2_X1 U3384 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_4/n4 ), .ZN(
        n3059) );
  NOR2_X1 U3385 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_5/n4 ), .ZN(
        n3060) );
  NOR2_X1 U3386 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_6/n4 ), .ZN(
        n3061) );
  NOR2_X1 U3387 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_7/n4 ), .ZN(
        n3062) );
  NOR2_X1 U3388 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_8/n4 ), .ZN(
        n3063) );
  NOR2_X1 U3389 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_9/n4 ), .ZN(
        n3064) );
  NOR2_X1 U3390 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_10/n4 ), .ZN(
        n3065) );
  NOR2_X1 U3391 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_11/n4 ), .ZN(
        n3066) );
  NOR2_X1 U3392 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_12/n4 ), .ZN(
        n3067) );
  NOR2_X1 U3393 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_13/n4 ), .ZN(
        n3068) );
  NOR2_X1 U3394 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_14/n4 ), .ZN(
        n3069) );
  NOR2_X1 U3395 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_15/n4 ), .ZN(
        n3070) );
  NOR2_X1 U3396 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_16/n4 ), .ZN(
        n3071) );
  NOR2_X1 U3397 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_17/n4 ), .ZN(
        n3072) );
  NOR2_X1 U3398 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_18/n4 ), .ZN(
        n3073) );
  NOR2_X1 U3399 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_19/n4 ), .ZN(
        n3074) );
  NOR2_X1 U3400 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_20/n4 ), .ZN(
        n3075) );
  NOR2_X1 U3401 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_21/n4 ), .ZN(
        n3076) );
  NOR2_X1 U3402 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_22/n4 ), .ZN(
        n3077) );
  NOR2_X1 U3403 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_23/n4 ), .ZN(
        n3078) );
  NOR2_X1 U3404 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_24/n4 ), .ZN(
        n3079) );
  NOR2_X1 U3405 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_25/n4 ), .ZN(
        n3080) );
  NOR2_X1 U3406 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_26/n4 ), .ZN(
        n3081) );
  NOR2_X1 U3407 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_27/n4 ), .ZN(
        n3082) );
  NOR2_X1 U3408 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_28/n4 ), .ZN(
        n3083) );
  NOR2_X1 U3409 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_29/n4 ), .ZN(
        n3084) );
  NOR2_X1 U3410 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_30/n4 ), .ZN(
        n3085) );
  NOR2_X1 U3411 ( .A1(RST), .A2(\unit_fetch/unit_npcregister/ffi_31/n4 ), .ZN(
        n3086) );
  NOR2_X1 U3412 ( .A1(RST), .A2(n1340), .ZN(
        \unit_control/uut_third_stage/ffi_15/n5 ) );
  NAND2_X1 U3413 ( .A1(\unit_control/uut_third_stage/ffi_15/n5 ), .A2(
        \cw_dec[2] ), .ZN(n2810) );
  OR2_X1 U3414 ( .A1(\unit_fetch/unit_instructionRegister/n63 ), .A2(n2810), 
        .ZN(n2812) );
  NAND4_X1 U3415 ( .A1(n1340), .A2(n3022), .A3(n1330), .A4(\cw_dec[2] ), .ZN(
        n2811) );
  OAI21_X1 U3416 ( .B1(n1687), .B2(n2812), .A(n2811), .ZN(n2934) );
  NOR4_X1 U3417 ( .A1(\unit_control/n153 ), .A2(\unit_control/n152 ), .A3(
        n2786), .A4(n2785), .ZN(\unit_control/next_state[0] ) );
  NOR3_X1 U3418 ( .A1(\unit_control/n153 ), .A2(\unit_control/n152 ), .A3(
        n2787), .ZN(\unit_control/next_state[1] ) );
  AND2_X1 U3419 ( .A1(\unit_control/cw2delay[3] ), .A2(n1943), .ZN(
        \unit_control/uut_fourth_stage/ffi_3/n6 ) );
  AND2_X1 U3420 ( .A1(\unit_control/cw2delay[4] ), .A2(n1943), .ZN(
        \unit_control/uut_fourth_stage/ffi_4/n5 ) );
  NOR2_X1 U3421 ( .A1(n2794), .A2(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n73 ) );
  INV_X1 U3422 ( .A(n2929), .ZN(n2793) );
  NAND2_X1 U3423 ( .A1(\unit_fetch/unit_instructionRegister/n73 ), .A2(n2793), 
        .ZN(n2792) );
  NAND2_X1 U3424 ( .A1(\unit_fetch/unit_programCounter/ffi_4/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_5/n4 ), .ZN(n2825) );
  NOR2_X1 U3425 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(n2825), 
        .ZN(n2788) );
  NOR4_X1 U3426 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n2798)
         );
  NAND2_X1 U3427 ( .A1(n1559), .A2(n2798), .ZN(
        \unit_fetch/unit_instructionRegister/n68 ) );
  AOI21_X1 U3428 ( .B1(n2792), .B2(\unit_fetch/unit_instructionRegister/n68 ), 
        .A(n2924), .ZN(\unit_control/uut_second_stage/ffi_10/n5 ) );
  NOR2_X1 U3429 ( .A1(n2924), .A2(\unit_fetch/unit_instructionRegister/n68 ), 
        .ZN(\unit_control/uut_second_stage/ffi_12/n5 ) );
  NOR2_X1 U3430 ( .A1(n2793), .A2(n2927), .ZN(
        \unit_fetch/unit_instructionRegister/n72 ) );
  NAND2_X1 U3431 ( .A1(n2924), .A2(\unit_fetch/unit_instructionRegister/n72 ), 
        .ZN(n2797) );
  NAND2_X1 U3432 ( .A1(n2924), .A2(n1559), .ZN(
        \unit_fetch/unit_instructionRegister/n70 ) );
  NOR3_X1 U3433 ( .A1(n2794), .A2(n2929), .A3(
        \unit_fetch/unit_instructionRegister/n70 ), .ZN(n6) );
  NAND2_X1 U3434 ( .A1(n2797), .A2(n1614), .ZN(
        \unit_control/uut_second_stage/ffi_13/n5 ) );
  NAND2_X1 U3435 ( .A1(\unit_fetch/unit_instructionRegister/n72 ), .A2(n2794), 
        .ZN(n2796) );
  INV_X1 U3436 ( .A(n2796), .ZN(\unit_control/uut_second_stage/ffi_14/n5 ) );
  NOR2_X1 U3437 ( .A1(n1605), .A2(n1932), .ZN(
        \unit_control/uut_second_stage/ffi_24/n3 ) );
  OR2_X1 U3438 ( .A1(n6), .A2(\unit_control/uut_second_stage/ffi_24/n3 ), .ZN(
        \unit_control/uut_second_stage/ffi_17/n5 ) );
  OAI21_X1 U3439 ( .B1(n2798), .B2(n2797), .A(n2796), .ZN(
        \unit_control/uut_second_stage/ffi_21/n5 ) );
  NOR2_X1 U3440 ( .A1(n2798), .A2(n1614), .ZN(
        \unit_control/uut_second_stage/ffi_3/n5 ) );
  AND2_X1 U3441 ( .A1(\unit_control/cw1delay[10] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_10/n5 ) );
  AND2_X1 U3442 ( .A1(\unit_control/cw1delay[12] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_12/n5 ) );
  AND2_X1 U3443 ( .A1(\unit_control/cw1delay[13] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_13/n5 ) );
  AND2_X1 U3444 ( .A1(\unit_control/cw1delay[14] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_14/n5 ) );
  AND2_X1 U3445 ( .A1(\unit_control/cw1delay[17] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_17/n6 ) );
  AND2_X1 U3446 ( .A1(\unit_control/cw1delay[3] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_3/n5 ) );
  AND2_X1 U3447 ( .A1(\unit_control/cw1delay[4] ), .A2(n1943), .ZN(
        \unit_control/uut_third_stage/ffi_4/n5 ) );
  AND2_X1 U3448 ( .A1(\unit_control/cw1delay[9] ), .A2(n1942), .ZN(
        \unit_control/uut_third_stage/ffi_9/n6 ) );
  NAND2_X1 U3449 ( .A1(n2808), .A2(n1668), .ZN(n2799) );
  OAI211_X1 U3450 ( .C1(\unit_fetch/unit_instructionRegister/n54 ), .C2(n2810), 
        .A(n2799), .B(n2811), .ZN(\unit_decode/IMMreg/ffi_16/n5 ) );
  NAND2_X1 U3451 ( .A1(n2808), .A2(n1666), .ZN(n2800) );
  OAI211_X1 U3452 ( .C1(\unit_fetch/unit_instructionRegister/n55 ), .C2(n2810), 
        .A(n2800), .B(n2811), .ZN(\unit_decode/IMMreg/ffi_17/n5 ) );
  NAND2_X1 U3453 ( .A1(n2808), .A2(n1679), .ZN(n2801) );
  OAI211_X1 U3454 ( .C1(\unit_fetch/unit_instructionRegister/n56 ), .C2(n2810), 
        .A(n2801), .B(n2811), .ZN(\unit_decode/IMMreg/ffi_18/n5 ) );
  NAND2_X1 U3455 ( .A1(n2808), .A2(n1675), .ZN(n2802) );
  OAI211_X1 U3456 ( .C1(\unit_fetch/unit_instructionRegister/n57 ), .C2(n2810), 
        .A(n2802), .B(n2811), .ZN(\unit_decode/IMMreg/ffi_19/n5 ) );
  OAI21_X1 U3457 ( .B1(n2810), .B2(\unit_fetch/unit_instructionRegister/n60 ), 
        .A(n2811), .ZN(n2803) );
  INV_X1 U3458 ( .A(n2803), .ZN(n2805) );
  OAI21_X1 U3459 ( .B1(\unit_decode/IMMreg/ffi_20/n4 ), .B2(n2932), .A(n2805), 
        .ZN(\unit_decode/IMMreg/ffi_20/n5 ) );
  OAI22_X1 U3460 ( .A1(n2810), .A2(\unit_fetch/unit_instructionRegister/n59 ), 
        .B1(n2932), .B2(\unit_decode/IMMreg/ffi_21/n4 ), .ZN(n2804) );
  INV_X1 U3461 ( .A(n2811), .ZN(n2807) );
  OR2_X1 U3462 ( .A1(n2804), .A2(n2807), .ZN(\unit_decode/IMMreg/ffi_21/n5 )
         );
  OAI21_X1 U3463 ( .B1(\unit_decode/IMMreg/ffi_22/n4 ), .B2(n2932), .A(n2805), 
        .ZN(\unit_decode/IMMreg/ffi_22/n5 ) );
  AOI21_X1 U3464 ( .B1(n2808), .B2(n1674), .A(n2807), .ZN(n2806) );
  OAI21_X1 U3465 ( .B1(\unit_fetch/unit_instructionRegister/n61 ), .B2(n2810), 
        .A(n2806), .ZN(\unit_decode/IMMreg/ffi_23/n5 ) );
  AOI21_X1 U3466 ( .B1(n2808), .B2(n1670), .A(n2807), .ZN(n2809) );
  OAI21_X1 U3467 ( .B1(\unit_fetch/unit_instructionRegister/n62 ), .B2(n2810), 
        .A(n2809), .ZN(\unit_decode/IMMreg/ffi_24/n5 ) );
  OAI211_X1 U3468 ( .C1(\unit_decode/IMMreg/ffi_25/n4 ), .C2(n2932), .A(n2812), 
        .B(n2811), .ZN(\unit_decode/IMMreg/ffi_25/n5 ) );
  NAND2_X1 U3469 ( .A1(\unit_control/uut_third_stage/ffi_17/n5 ), .A2(n1942), 
        .ZN(n471) );
  NOR2_X1 U3470 ( .A1(n2818), .A2(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n67 ) );
  NOR2_X1 U3471 ( .A1(n2813), .A2(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n71 ) );
  NOR2_X1 U3472 ( .A1(n2814), .A2(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n74 ) );
  AND2_X1 U3473 ( .A1(n2815), .A2(n1559), .ZN(
        \unit_fetch/unit_instructionRegister/n75 ) );
  NOR2_X1 U3474 ( .A1(n2816), .A2(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n78 ) );
  INV_X1 U3475 ( .A(n2817), .ZN(n2826) );
  NOR2_X1 U3476 ( .A1(\unit_fetch/unit_programCounter/ffi_3/n4 ), .A2(n2825), 
        .ZN(n2883) );
  NAND2_X1 U3477 ( .A1(n2826), .A2(n2883), .ZN(n2873) );
  AOI21_X1 U3478 ( .B1(n2818), .B2(n2873), .A(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n77 ) );
  NAND2_X1 U3479 ( .A1(n2878), .A2(n2883), .ZN(n2823) );
  NAND2_X1 U3480 ( .A1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .ZN(n2856) );
  INV_X1 U3481 ( .A(n2878), .ZN(n2819) );
  NOR3_X1 U3482 ( .A1(n1607), .A2(n2824), .A3(n2867), .ZN(n2868) );
  INV_X1 U3483 ( .A(n2868), .ZN(n2820) );
  OAI221_X1 U3484 ( .B1(n2823), .B2(n1603), .C1(n2823), .C2(n2856), .A(n2820), 
        .ZN(n2842) );
  NOR3_X1 U3485 ( .A1(\unit_fetch/pc_regout[1] ), .A2(
        \unit_fetch/pc_regout[0] ), .A3(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .ZN(n2893) );
  NAND2_X1 U3486 ( .A1(n2889), .A2(n2893), .ZN(n2879) );
  OAI211_X1 U3487 ( .C1(n1587), .C2(n1603), .A(n2873), .B(n2879), .ZN(n2834)
         );
  NOR2_X1 U3488 ( .A1(n2842), .A2(n2834), .ZN(n2821) );
  NOR3_X1 U3489 ( .A1(\unit_fetch/pc_regout[1] ), .A2(
        \unit_fetch/unit_programCounter/ffi_2/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_0/n4 ), .ZN(n2827) );
  NAND2_X1 U3490 ( .A1(n2878), .A2(n2827), .ZN(n2838) );
  INV_X1 U3491 ( .A(n2838), .ZN(n2849) );
  NAND2_X1 U3492 ( .A1(n2883), .A2(n2849), .ZN(n2844) );
  AOI21_X1 U3493 ( .B1(n2821), .B2(n2844), .A(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n79 ) );
  OAI21_X1 U3494 ( .B1(n2822), .B2(n2893), .A(n2901), .ZN(n2846) );
  OR2_X1 U3495 ( .A1(n2824), .A2(n2823), .ZN(n2836) );
  NOR2_X1 U3496 ( .A1(n1607), .A2(n2825), .ZN(n2848) );
  NAND2_X1 U3497 ( .A1(n2826), .A2(n2848), .ZN(n2832) );
  INV_X1 U3498 ( .A(n2832), .ZN(n2843) );
  AOI211_X1 U3499 ( .C1(n2901), .C2(n2827), .A(n2834), .B(n2843), .ZN(n2831)
         );
  NOR2_X1 U3500 ( .A1(\unit_fetch/unit_programCounter/ffi_0/n4 ), .A2(n2829), 
        .ZN(n2855) );
  INV_X1 U3501 ( .A(n2855), .ZN(n2874) );
  AOI21_X1 U3502 ( .B1(n2847), .B2(n2874), .A(n2867), .ZN(n2896) );
  INV_X1 U3503 ( .A(n2896), .ZN(n2830) );
  AOI21_X1 U3504 ( .B1(n2831), .B2(n2830), .A(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n81 ) );
  OAI21_X1 U3505 ( .B1(n2867), .B2(n2833), .A(n2832), .ZN(n2906) );
  AOI211_X1 U3506 ( .C1(n2893), .C2(n2901), .A(n2834), .B(n2906), .ZN(n2835)
         );
  NOR2_X1 U3507 ( .A1(n2835), .A2(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n82 ) );
  OAI21_X1 U3508 ( .B1(n2847), .B2(n1587), .A(n2836), .ZN(n2871) );
  AOI21_X1 U3509 ( .B1(n2876), .B2(n2856), .A(n1587), .ZN(n2837) );
  OAI21_X1 U3510 ( .B1(n2871), .B2(n2837), .A(n1559), .ZN(n2841) );
  INV_X1 U3511 ( .A(n2841), .ZN(\unit_fetch/unit_instructionRegister/n83 ) );
  OAI22_X1 U3512 ( .A1(n2839), .A2(n2838), .B1(n1365), .B2(n2874), .ZN(n2840)
         );
  INV_X1 U3513 ( .A(n2840), .ZN(n2852) );
  OAI21_X1 U3514 ( .B1(n2852), .B2(n1932), .A(n2841), .ZN(
        \unit_fetch/unit_instructionRegister/n86 ) );
  OAI21_X1 U3515 ( .B1(n1932), .B2(n2844), .A(n2841), .ZN(
        \unit_fetch/unit_instructionRegister/n85 ) );
  NOR2_X1 U3516 ( .A1(n2843), .A2(n2842), .ZN(n2892) );
  INV_X1 U3517 ( .A(n2844), .ZN(n2898) );
  AOI21_X1 U3518 ( .B1(n2892), .B2(n2850), .A(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n87 ) );
  OAI211_X1 U3519 ( .C1(n2847), .C2(n2867), .A(n2846), .B(n2873), .ZN(n2851)
         );
  NAND2_X1 U3520 ( .A1(n2849), .A2(n2848), .ZN(n2890) );
  NAND2_X1 U3521 ( .A1(n2850), .A2(n2890), .ZN(n2854) );
  NOR2_X1 U3522 ( .A1(n2851), .A2(n2854), .ZN(n2853) );
  AOI21_X1 U3523 ( .B1(n2853), .B2(n2852), .A(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n88 ) );
  AOI21_X1 U3524 ( .B1(n2855), .B2(n2901), .A(n2854), .ZN(n2870) );
  AOI221_X1 U3525 ( .B1(n2856), .B2(n2870), .C1(n2867), .C2(n2870), .A(n1933), 
        .ZN(\unit_fetch/unit_instructionRegister/n89 ) );
  NOR4_X1 U3526 ( .A1(\unit_fetch/unit_programCounter/ffi_18/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_20/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_28/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_10/n4 ), .ZN(n2860) );
  NOR4_X1 U3527 ( .A1(\unit_fetch/unit_programCounter/ffi_7/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_22/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_30/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_26/n4 ), .ZN(n2859) );
  NOR4_X1 U3528 ( .A1(\unit_fetch/unit_programCounter/ffi_27/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_16/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_23/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_24/n4 ), .ZN(n2858) );
  NOR4_X1 U3529 ( .A1(\unit_fetch/unit_programCounter/ffi_12/n4 ), .A2(
        \unit_fetch/unit_adder/add_19/n47 ), .A3(
        \unit_fetch/unit_programCounter/ffi_6/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_14/n4 ), .ZN(n2857) );
  NAND4_X1 U3530 ( .A1(n2860), .A2(n2859), .A3(n2858), .A4(n2857), .ZN(n2866)
         );
  NOR4_X1 U3531 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_4/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_25/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_17/n4 ), .ZN(n2864) );
  NOR4_X1 U3532 ( .A1(\unit_fetch/unit_programCounter/ffi_8/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_9/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_21/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_29/n4 ), .ZN(n2863) );
  NOR4_X1 U3533 ( .A1(\unit_fetch/unit_programCounter/ffi_3/n4 ), .A2(
        \unit_fetch/unit_programCounter/ffi_5/n4 ), .A3(
        \unit_fetch/unit_programCounter/ffi_15/n4 ), .A4(
        \unit_fetch/unit_programCounter/ffi_19/n4 ), .ZN(n2862) );
  NAND4_X1 U3534 ( .A1(n2864), .A2(n2863), .A3(n2862), .A4(n2861), .ZN(n2865)
         );
  NOR2_X1 U3535 ( .A1(n2866), .A2(n2865), .ZN(n2907) );
  NOR2_X1 U3536 ( .A1(n2876), .A2(n2867), .ZN(n2897) );
  AOI211_X1 U3537 ( .C1(n2869), .C2(n2907), .A(n2897), .B(n2868), .ZN(n2904)
         );
  AOI21_X1 U3538 ( .B1(n2870), .B2(n2904), .A(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n90 ) );
  INV_X1 U3539 ( .A(n2871), .ZN(n2872) );
  OAI211_X1 U3540 ( .C1(n1587), .C2(n2874), .A(n2873), .B(n2872), .ZN(n2888)
         );
  NOR2_X1 U3541 ( .A1(n2876), .A2(n1587), .ZN(n2877) );
  OAI21_X1 U3542 ( .B1(n2888), .B2(n2877), .A(n1559), .ZN(n2885) );
  INV_X1 U3543 ( .A(n2885), .ZN(\unit_fetch/unit_instructionRegister/n91 ) );
  AND2_X1 U3544 ( .A1(n2878), .A2(n2893), .ZN(n2884) );
  OAI21_X1 U3545 ( .B1(n2887), .B2(n1365), .A(n2879), .ZN(n2881) );
  AOI21_X1 U3546 ( .B1(n2882), .B2(n2884), .A(n2881), .ZN(n2900) );
  OAI21_X1 U3547 ( .B1(n2900), .B2(n1932), .A(n2885), .ZN(
        \unit_fetch/unit_instructionRegister/n94 ) );
  NAND3_X1 U3548 ( .A1(n1559), .A2(n2884), .A3(n2883), .ZN(n2886) );
  NAND2_X1 U3549 ( .A1(n2886), .A2(n2885), .ZN(
        \unit_fetch/unit_instructionRegister/n93 ) );
  INV_X1 U3550 ( .A(n2887), .ZN(n2902) );
  AOI21_X1 U3551 ( .B1(n2889), .B2(n2902), .A(n2888), .ZN(n2895) );
  AND2_X1 U3552 ( .A1(n2890), .A2(n2895), .ZN(n2891) );
  AOI21_X1 U3553 ( .B1(n2892), .B2(n2891), .A(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n95 ) );
  NAND2_X1 U3554 ( .A1(n2893), .A2(n2901), .ZN(n2894) );
  NAND2_X1 U3555 ( .A1(n2895), .A2(n2894), .ZN(n2905) );
  NOR4_X1 U3556 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2905), .ZN(n2899)
         );
  AOI21_X1 U3557 ( .B1(n2900), .B2(n2899), .A(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n96 ) );
  AOI21_X1 U3558 ( .B1(n2902), .B2(n2901), .A(n2905), .ZN(n2903) );
  AOI21_X1 U3559 ( .B1(n2904), .B2(n2903), .A(n1932), .ZN(
        \unit_fetch/unit_instructionRegister/n97 ) );
  AOI211_X1 U3560 ( .C1(n2908), .C2(n2907), .A(n2906), .B(n2905), .ZN(n2909)
         );
  NOR2_X1 U3561 ( .A1(n2909), .A2(n1933), .ZN(
        \unit_fetch/unit_instructionRegister/n98 ) );
  NAND2_X1 U3562 ( .A1(n1931), .A2(n2910), .ZN(n2921) );
  NAND2_X1 U3563 ( .A1(n1926), .A2(\unit_fetch/pc_regout[1] ), .ZN(n2911) );
  OAI211_X1 U3564 ( .C1(\unit_fetch/unit_npcregister/ffi_1/n4 ), .C2(n1923), 
        .A(n2921), .B(n2911), .ZN(\unit_fetch/unit_npcregister/ffi_1/n5 ) );
  AOI22_X1 U3565 ( .A1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .A2(n1926), 
        .B1(n1929), .B2(n2915), .ZN(n2923) );
  OAI21_X1 U3566 ( .B1(\unit_fetch/unit_npcregister/ffi_2/n4 ), .B2(n1924), 
        .A(n2923), .ZN(\unit_fetch/unit_npcregister/ffi_2/n5 ) );
  OAI21_X1 U3567 ( .B1(\unit_fetch/unit_programCounter/ffi_1/n4 ), .B2(n2922), 
        .A(n2921), .ZN(\unit_fetch/unit_programCounter/ffi_1/n5 ) );
  OAI21_X1 U3568 ( .B1(\unit_fetch/unit_programCounter/ffi_2/n4 ), .B2(n1924), 
        .A(n2923), .ZN(\unit_fetch/unit_programCounter/ffi_2/n5 ) );
  AOI22_X1 U3569 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_0/n5 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_0/n4 ), .B2(n1685), .ZN(wr_data[0])
         );
  AOI22_X1 U3570 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_10/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_10/n4 ), .B2(n1685), .ZN(wr_data[10]) );
  AOI22_X1 U3571 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_11/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_11/n4 ), .B2(n1685), .ZN(wr_data[11]) );
  AOI22_X1 U3572 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_12/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_12/n4 ), .B2(n1685), .ZN(wr_data[12]) );
  AOI22_X1 U3573 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_13/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_13/n4 ), .B2(n1685), .ZN(wr_data[13]) );
  AOI22_X1 U3574 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_14/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_14/n4 ), .B2(n1685), .ZN(wr_data[14]) );
  AOI22_X1 U3575 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_15/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_15/n4 ), .B2(n1685), .ZN(wr_data[15]) );
  AOI22_X1 U3576 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_16/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_16/n4 ), .B2(n1685), .ZN(wr_data[16]) );
  AOI22_X1 U3577 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_17/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_17/n4 ), .B2(n1685), .ZN(wr_data[17]) );
  AOI22_X1 U3578 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_18/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_18/n4 ), .B2(n1685), .ZN(wr_data[18]) );
  AOI22_X1 U3579 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_19/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_19/n4 ), .B2(n1685), .ZN(wr_data[19]) );
  AOI22_X1 U3580 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_1/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_1/n4 ), .B2(n1685), .ZN(wr_data[1])
         );
  AOI22_X1 U3581 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_20/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_20/n4 ), .B2(n1685), .ZN(wr_data[20]) );
  AOI22_X1 U3582 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_21/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_21/n4 ), .B2(n1685), .ZN(wr_data[21]) );
  AOI22_X1 U3583 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_22/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_22/n4 ), .B2(n1685), .ZN(wr_data[22]) );
  AOI22_X1 U3584 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_23/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_23/n4 ), .B2(n1685), .ZN(wr_data[23]) );
  AOI22_X1 U3585 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_24/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_24/n4 ), .B2(n1685), .ZN(wr_data[24]) );
  AOI22_X1 U3586 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_25/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_25/n4 ), .B2(n1685), .ZN(wr_data[25]) );
  AOI22_X1 U3587 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_26/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_26/n4 ), .B2(n1685), .ZN(wr_data[26]) );
  AOI22_X1 U3588 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_27/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_27/n4 ), .B2(n1685), .ZN(wr_data[27]) );
  AOI22_X1 U3589 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_28/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_28/n4 ), .B2(n1685), .ZN(wr_data[28]) );
  AOI22_X1 U3590 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_29/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_29/n4 ), .B2(n1685), .ZN(wr_data[29]) );
  AOI22_X1 U3591 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_2/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_2/n4 ), .B2(n1685), .ZN(wr_data[2])
         );
  AOI22_X1 U3592 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_30/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_30/n4 ), .B2(n1685), .ZN(wr_data[30]) );
  AOI22_X1 U3593 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_31/n4 ), .B1(\unit_execution/COMP_NPC2/ffi_31/n4 ), .B2(n1685), .ZN(wr_data[31]) );
  AOI22_X1 U3594 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_3/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_3/n4 ), .B2(n1685), .ZN(wr_data[3])
         );
  AOI22_X1 U3595 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_4/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_4/n4 ), .B2(n1685), .ZN(wr_data[4])
         );
  AOI22_X1 U3596 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_5/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_5/n4 ), .B2(n1685), .ZN(wr_data[5])
         );
  AOI22_X1 U3597 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_6/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_6/n4 ), .B2(n1685), .ZN(wr_data[6])
         );
  AOI22_X1 U3598 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_7/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_7/n4 ), .B2(n1685), .ZN(wr_data[7])
         );
  AOI22_X1 U3599 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_8/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_8/n4 ), .B2(n1685), .ZN(wr_data[8])
         );
  AOI22_X1 U3600 ( .A1(n1650), .A2(\unit_execution/COMP_REGN_ALUOUT/ffi_9/n4 ), 
        .B1(\unit_execution/COMP_NPC2/ffi_9/n4 ), .B2(n1685), .ZN(wr_data[9])
         );
  INV_X1 U3601 ( .A(n2924), .ZN(n2928) );
  AOI21_X1 U3602 ( .B1(n2925), .B2(n2928), .A(n2929), .ZN(n2926) );
  AOI211_X1 U3603 ( .C1(n2929), .C2(n2928), .A(n1932), .B(n2926), .ZN(n2930)
         );
  OR3_X1 U3604 ( .A1(\unit_control/uut_second_stage/ffi_3/n5 ), .A2(n2930), 
        .A3(\unit_control/uut_second_stage/ffi_21/n5 ), .ZN(n4) );
endmodule

